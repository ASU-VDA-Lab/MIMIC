module fake_aes_9343_n_653 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_653);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_653;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_529;
wire n_455;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_24), .Y(n_80) );
BUFx2_ASAP7_75t_L g81 ( .A(n_69), .Y(n_81) );
BUFx2_ASAP7_75t_L g82 ( .A(n_34), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_60), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_30), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_47), .Y(n_85) );
CKINVDCx14_ASAP7_75t_R g86 ( .A(n_50), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_12), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_13), .Y(n_88) );
CKINVDCx16_ASAP7_75t_R g89 ( .A(n_65), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_70), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_16), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_39), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_5), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_36), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_8), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_54), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_1), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_3), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_78), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_68), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_6), .Y(n_101) );
CKINVDCx14_ASAP7_75t_R g102 ( .A(n_19), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_9), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_38), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_48), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_55), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_63), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_62), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_40), .Y(n_109) );
CKINVDCx14_ASAP7_75t_R g110 ( .A(n_6), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_42), .Y(n_111) );
INVxp67_ASAP7_75t_L g112 ( .A(n_31), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_51), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_9), .Y(n_114) );
CKINVDCx14_ASAP7_75t_R g115 ( .A(n_75), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_64), .Y(n_116) );
CKINVDCx16_ASAP7_75t_R g117 ( .A(n_8), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_22), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_85), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_80), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_80), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_102), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_83), .Y(n_123) );
NAND2xp33_ASAP7_75t_L g124 ( .A(n_84), .B(n_32), .Y(n_124) );
NOR2xp33_ASAP7_75t_SL g125 ( .A(n_89), .B(n_79), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_85), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_83), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_81), .B(n_0), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_90), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_94), .Y(n_130) );
OAI22xp5_ASAP7_75t_L g131 ( .A1(n_110), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_81), .B(n_2), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_94), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_107), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_90), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_107), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_92), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_92), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_96), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_89), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_82), .B(n_3), .Y(n_141) );
AO22x1_ASAP7_75t_L g142 ( .A1(n_87), .A2(n_4), .B1(n_5), .B2(n_7), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_96), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_100), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_100), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_104), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_82), .B(n_4), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_104), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_112), .B(n_7), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_106), .Y(n_150) );
BUFx10_ASAP7_75t_L g151 ( .A(n_140), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g152 ( .A(n_122), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_120), .B(n_106), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_120), .B(n_111), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_126), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_132), .B(n_117), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_126), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_121), .B(n_113), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_126), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_138), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_121), .B(n_109), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_126), .Y(n_162) );
AND2x2_ASAP7_75t_SL g163 ( .A(n_125), .B(n_111), .Y(n_163) );
INVx4_ASAP7_75t_SL g164 ( .A(n_126), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_126), .Y(n_165) );
INVxp33_ASAP7_75t_SL g166 ( .A(n_132), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_126), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_130), .Y(n_168) );
AND2x2_ASAP7_75t_L g169 ( .A(n_132), .B(n_86), .Y(n_169) );
NAND3xp33_ASAP7_75t_L g170 ( .A(n_123), .B(n_113), .C(n_101), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_123), .B(n_115), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_130), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_127), .B(n_99), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_130), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_130), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_127), .B(n_118), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_130), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_130), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_129), .B(n_105), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_130), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_119), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_144), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_129), .B(n_118), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_144), .Y(n_184) );
BUFx3_ASAP7_75t_L g185 ( .A(n_119), .Y(n_185) );
BUFx3_ASAP7_75t_L g186 ( .A(n_119), .Y(n_186) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_133), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_144), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_133), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_160), .Y(n_190) );
INVx2_ASAP7_75t_SL g191 ( .A(n_160), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_160), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_166), .B(n_128), .Y(n_193) );
HB1xp67_ASAP7_75t_L g194 ( .A(n_169), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_160), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_169), .B(n_156), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_171), .B(n_138), .Y(n_197) );
NOR2x1_ASAP7_75t_R g198 ( .A(n_171), .B(n_128), .Y(n_198) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_185), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_182), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_176), .B(n_141), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_182), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_176), .B(n_141), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_163), .A2(n_125), .B1(n_131), .B2(n_148), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_183), .B(n_147), .Y(n_205) );
BUFx3_ASAP7_75t_L g206 ( .A(n_185), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_163), .B(n_147), .Y(n_207) );
BUFx3_ASAP7_75t_L g208 ( .A(n_185), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_184), .Y(n_209) );
INVx4_ASAP7_75t_L g210 ( .A(n_163), .Y(n_210) );
INVx3_ASAP7_75t_L g211 ( .A(n_186), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_179), .B(n_138), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_173), .B(n_138), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_152), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_187), .Y(n_215) );
BUFx4f_ASAP7_75t_SL g216 ( .A(n_151), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_151), .B(n_149), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_183), .B(n_135), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_161), .B(n_149), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_187), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_187), .Y(n_221) );
OAI22xp5_ASAP7_75t_SL g222 ( .A1(n_153), .A2(n_131), .B1(n_116), .B2(n_98), .Y(n_222) );
INVx8_ASAP7_75t_L g223 ( .A(n_187), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_187), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_153), .B(n_135), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_158), .A2(n_148), .B1(n_143), .B2(n_137), .Y(n_226) );
INVx2_ASAP7_75t_SL g227 ( .A(n_186), .Y(n_227) );
AOI21xp33_ASAP7_75t_L g228 ( .A1(n_184), .A2(n_124), .B(n_143), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_170), .A2(n_139), .B1(n_137), .B2(n_142), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_187), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_188), .Y(n_231) );
NAND2xp33_ASAP7_75t_L g232 ( .A(n_158), .B(n_139), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_188), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_186), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_181), .Y(n_235) );
AND2x4_ASAP7_75t_L g236 ( .A(n_170), .B(n_150), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_154), .B(n_146), .Y(n_237) );
BUFx12f_ASAP7_75t_L g238 ( .A(n_151), .Y(n_238) );
BUFx2_ASAP7_75t_L g239 ( .A(n_238), .Y(n_239) );
NOR2x1_ASAP7_75t_L g240 ( .A(n_210), .B(n_146), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_235), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_235), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_192), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_200), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_197), .A2(n_181), .B(n_172), .Y(n_245) );
INVx3_ASAP7_75t_L g246 ( .A(n_206), .Y(n_246) );
AOI222xp33_ASAP7_75t_L g247 ( .A1(n_222), .A2(n_142), .B1(n_88), .B2(n_91), .C1(n_93), .C2(n_87), .Y(n_247) );
INVx5_ASAP7_75t_L g248 ( .A(n_223), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_203), .B(n_151), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_203), .B(n_146), .Y(n_250) );
BUFx3_ASAP7_75t_L g251 ( .A(n_238), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_197), .A2(n_181), .B(n_155), .Y(n_252) );
AOI222xp33_ASAP7_75t_L g253 ( .A1(n_222), .A2(n_88), .B1(n_91), .B2(n_93), .C1(n_114), .C2(n_97), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_192), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_193), .B(n_95), .Y(n_255) );
NAND2xp33_ASAP7_75t_L g256 ( .A(n_201), .B(n_189), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_204), .A2(n_150), .B1(n_146), .B2(n_145), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_200), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_203), .B(n_150), .Y(n_259) );
BUFx2_ASAP7_75t_L g260 ( .A(n_238), .Y(n_260) );
OR2x6_ASAP7_75t_L g261 ( .A(n_210), .B(n_97), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_192), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_202), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_202), .Y(n_264) );
AND2x4_ASAP7_75t_L g265 ( .A(n_203), .B(n_150), .Y(n_265) );
NOR2xp67_ASAP7_75t_SL g266 ( .A(n_206), .B(n_189), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_232), .A2(n_172), .B(n_180), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_201), .B(n_145), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_198), .B(n_101), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_205), .B(n_145), .Y(n_270) );
OR2x2_ASAP7_75t_L g271 ( .A(n_205), .B(n_114), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_218), .B(n_103), .Y(n_272) );
INVx3_ASAP7_75t_L g273 ( .A(n_206), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_209), .Y(n_274) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_194), .Y(n_275) );
NOR2xp33_ASAP7_75t_SL g276 ( .A(n_216), .B(n_108), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_227), .B(n_189), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_212), .A2(n_165), .B(n_180), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_209), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_231), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_212), .A2(n_165), .B(n_178), .Y(n_281) );
AOI221xp5_ASAP7_75t_L g282 ( .A1(n_196), .A2(n_103), .B1(n_133), .B2(n_134), .C(n_136), .Y(n_282) );
AND2x4_ASAP7_75t_L g283 ( .A(n_218), .B(n_136), .Y(n_283) );
BUFx6f_ASAP7_75t_L g284 ( .A(n_208), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_225), .B(n_196), .Y(n_285) );
A2O1A1Ixp33_ASAP7_75t_L g286 ( .A1(n_244), .A2(n_204), .B(n_219), .C(n_229), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_251), .Y(n_287) );
AND2x4_ASAP7_75t_L g288 ( .A(n_285), .B(n_225), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_270), .B(n_194), .Y(n_289) );
NOR2x1_ASAP7_75t_SL g290 ( .A(n_261), .B(n_210), .Y(n_290) );
OAI21x1_ASAP7_75t_L g291 ( .A1(n_278), .A2(n_220), .B(n_215), .Y(n_291) );
AOI21x1_ASAP7_75t_L g292 ( .A1(n_266), .A2(n_155), .B(n_175), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_270), .Y(n_293) );
OAI21x1_ASAP7_75t_L g294 ( .A1(n_281), .A2(n_224), .B(n_215), .Y(n_294) );
OAI21x1_ASAP7_75t_L g295 ( .A1(n_257), .A2(n_224), .B(n_215), .Y(n_295) );
AND2x4_ASAP7_75t_L g296 ( .A(n_248), .B(n_210), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_259), .Y(n_297) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_248), .Y(n_298) );
OAI21x1_ASAP7_75t_L g299 ( .A1(n_240), .A2(n_220), .B(n_224), .Y(n_299) );
OA21x2_ASAP7_75t_L g300 ( .A1(n_244), .A2(n_207), .B(n_178), .Y(n_300) );
AO32x2_ASAP7_75t_L g301 ( .A1(n_256), .A2(n_226), .A3(n_227), .B1(n_191), .B2(n_198), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_263), .Y(n_302) );
NAND2xp33_ASAP7_75t_L g303 ( .A(n_248), .B(n_227), .Y(n_303) );
O2A1O1Ixp33_ASAP7_75t_L g304 ( .A1(n_269), .A2(n_226), .B(n_213), .C(n_237), .Y(n_304) );
AOI21x1_ASAP7_75t_L g305 ( .A1(n_266), .A2(n_175), .B(n_177), .Y(n_305) );
OA21x2_ASAP7_75t_L g306 ( .A1(n_258), .A2(n_177), .B(n_168), .Y(n_306) );
OAI21x1_ASAP7_75t_L g307 ( .A1(n_240), .A2(n_220), .B(n_230), .Y(n_307) );
OR2x6_ASAP7_75t_L g308 ( .A(n_261), .B(n_249), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_271), .B(n_214), .Y(n_309) );
OAI21x1_ASAP7_75t_L g310 ( .A1(n_267), .A2(n_230), .B(n_231), .Y(n_310) );
A2O1A1Ixp33_ASAP7_75t_L g311 ( .A1(n_258), .A2(n_229), .B(n_237), .C(n_213), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_259), .B(n_233), .Y(n_312) );
OAI21x1_ASAP7_75t_L g313 ( .A1(n_280), .A2(n_230), .B(n_233), .Y(n_313) );
OAI21x1_ASAP7_75t_L g314 ( .A1(n_280), .A2(n_167), .B(n_157), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_248), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_259), .B(n_199), .Y(n_316) );
O2A1O1Ixp33_ASAP7_75t_L g317 ( .A1(n_272), .A2(n_217), .B(n_228), .C(n_199), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_259), .B(n_236), .Y(n_318) );
A2O1A1Ixp33_ASAP7_75t_L g319 ( .A1(n_263), .A2(n_236), .B(n_228), .C(n_195), .Y(n_319) );
OAI21x1_ASAP7_75t_L g320 ( .A1(n_264), .A2(n_157), .B(n_167), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g321 ( .A1(n_311), .A2(n_256), .B(n_277), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_288), .B(n_265), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g323 ( .A1(n_288), .A2(n_255), .B1(n_261), .B2(n_276), .Y(n_323) );
AND2x4_ASAP7_75t_L g324 ( .A(n_288), .B(n_265), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_309), .A2(n_261), .B1(n_247), .B2(n_253), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_308), .A2(n_271), .B1(n_264), .B2(n_279), .Y(n_326) );
AND2x4_ASAP7_75t_L g327 ( .A(n_296), .B(n_315), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_309), .A2(n_283), .B1(n_275), .B2(n_265), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_289), .B(n_265), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_308), .A2(n_283), .B1(n_282), .B2(n_239), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_293), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_312), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_308), .A2(n_279), .B1(n_274), .B2(n_283), .Y(n_333) );
OAI221xp5_ASAP7_75t_L g334 ( .A1(n_286), .A2(n_239), .B1(n_260), .B2(n_268), .C(n_251), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_302), .Y(n_335) );
O2A1O1Ixp33_ASAP7_75t_L g336 ( .A1(n_304), .A2(n_250), .B(n_283), .C(n_274), .Y(n_336) );
OAI21x1_ASAP7_75t_L g337 ( .A1(n_295), .A2(n_245), .B(n_252), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_308), .A2(n_260), .B1(n_242), .B2(n_241), .Y(n_338) );
AO21x1_ASAP7_75t_L g339 ( .A1(n_295), .A2(n_242), .B(n_241), .Y(n_339) );
AOI22xp33_ASAP7_75t_SL g340 ( .A1(n_290), .A2(n_248), .B1(n_284), .B2(n_246), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_312), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g342 ( .A1(n_297), .A2(n_236), .B1(n_134), .B2(n_136), .C(n_189), .Y(n_342) );
OAI222xp33_ASAP7_75t_L g343 ( .A1(n_287), .A2(n_248), .B1(n_254), .B2(n_243), .C1(n_262), .C2(n_134), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_316), .A2(n_284), .B1(n_243), .B2(n_262), .Y(n_344) );
AOI221xp5_ASAP7_75t_L g345 ( .A1(n_317), .A2(n_236), .B1(n_189), .B2(n_190), .C(n_195), .Y(n_345) );
AOI221xp5_ASAP7_75t_L g346 ( .A1(n_318), .A2(n_189), .B1(n_190), .B2(n_234), .C(n_191), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_318), .A2(n_273), .B1(n_246), .B2(n_191), .Y(n_347) );
A2O1A1Ixp33_ASAP7_75t_L g348 ( .A1(n_302), .A2(n_254), .B(n_234), .C(n_246), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_335), .B(n_301), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_335), .B(n_301), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_331), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_325), .B(n_287), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_326), .B(n_300), .Y(n_353) );
BUFx3_ASAP7_75t_L g354 ( .A(n_327), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_339), .Y(n_355) );
AOI22xp33_ASAP7_75t_SL g356 ( .A1(n_333), .A2(n_298), .B1(n_296), .B2(n_315), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_339), .Y(n_357) );
INVxp67_ASAP7_75t_SL g358 ( .A(n_336), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_332), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_337), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_344), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_341), .B(n_319), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_337), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_334), .A2(n_296), .B1(n_298), .B2(n_315), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_348), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_329), .B(n_300), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_348), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_327), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_327), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_322), .B(n_301), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_322), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_324), .B(n_301), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_324), .B(n_301), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_324), .B(n_313), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_321), .Y(n_375) );
INVx2_ASAP7_75t_SL g376 ( .A(n_340), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_345), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_338), .B(n_313), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_360), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_349), .Y(n_380) );
OAI21xp5_ASAP7_75t_L g381 ( .A1(n_377), .A2(n_323), .B(n_330), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_360), .A2(n_303), .B(n_310), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_370), .B(n_300), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_370), .B(n_300), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_349), .Y(n_385) );
BUFx2_ASAP7_75t_L g386 ( .A(n_374), .Y(n_386) );
INVxp67_ASAP7_75t_SL g387 ( .A(n_360), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_349), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_350), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_370), .B(n_306), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_352), .A2(n_328), .B1(n_346), .B2(n_347), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_372), .B(n_298), .Y(n_392) );
INVx5_ASAP7_75t_L g393 ( .A(n_376), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_352), .B(n_10), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_372), .B(n_298), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_372), .B(n_298), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_360), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_373), .B(n_306), .Y(n_398) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_351), .A2(n_342), .B1(n_343), .B2(n_303), .C(n_211), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_350), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_350), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_355), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_373), .B(n_306), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_355), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_357), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_351), .B(n_10), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_357), .Y(n_407) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_374), .Y(n_408) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_374), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_373), .B(n_306), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_363), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_371), .B(n_310), .Y(n_412) );
NOR3xp33_ASAP7_75t_L g413 ( .A(n_358), .B(n_307), .C(n_299), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_359), .B(n_294), .Y(n_414) );
AOI221xp5_ASAP7_75t_L g415 ( .A1(n_359), .A2(n_211), .B1(n_168), .B2(n_162), .C(n_167), .Y(n_415) );
OAI33xp33_ASAP7_75t_L g416 ( .A1(n_362), .A2(n_11), .A3(n_12), .B1(n_13), .B2(n_14), .B3(n_15), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_366), .B(n_11), .Y(n_417) );
OAI21x1_ASAP7_75t_L g418 ( .A1(n_363), .A2(n_291), .B(n_294), .Y(n_418) );
OAI321xp33_ASAP7_75t_L g419 ( .A1(n_376), .A2(n_292), .A3(n_305), .B1(n_284), .B2(n_159), .C(n_174), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_371), .B(n_299), .Y(n_420) );
INVx1_ASAP7_75t_SL g421 ( .A(n_354), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_380), .B(n_368), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_394), .A2(n_376), .B1(n_377), .B2(n_356), .Y(n_423) );
OAI211xp5_ASAP7_75t_L g424 ( .A1(n_381), .A2(n_356), .B(n_364), .C(n_358), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_408), .B(n_353), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_408), .B(n_409), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_406), .B(n_354), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_409), .B(n_378), .Y(n_428) );
AND2x4_ASAP7_75t_L g429 ( .A(n_393), .B(n_363), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_386), .B(n_353), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_417), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_386), .B(n_378), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_380), .B(n_353), .Y(n_433) );
BUFx2_ASAP7_75t_L g434 ( .A(n_393), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_417), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_385), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_379), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_385), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_416), .A2(n_362), .B1(n_375), .B2(n_364), .C(n_367), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_388), .B(n_378), .Y(n_440) );
BUFx3_ASAP7_75t_L g441 ( .A(n_421), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_388), .B(n_363), .Y(n_442) );
INVx1_ASAP7_75t_SL g443 ( .A(n_421), .Y(n_443) );
NAND5xp2_ASAP7_75t_SL g444 ( .A(n_381), .B(n_14), .C(n_15), .D(n_16), .E(n_17), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_389), .B(n_375), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_389), .B(n_369), .Y(n_446) );
NAND4xp25_ASAP7_75t_L g447 ( .A(n_391), .B(n_369), .C(n_368), .D(n_354), .Y(n_447) );
INVx1_ASAP7_75t_SL g448 ( .A(n_392), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_379), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_400), .B(n_365), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_400), .B(n_365), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_402), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_401), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_401), .Y(n_454) );
AOI31xp33_ASAP7_75t_L g455 ( .A1(n_416), .A2(n_369), .A3(n_368), .B(n_366), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_384), .B(n_367), .Y(n_456) );
INVx2_ASAP7_75t_SL g457 ( .A(n_393), .Y(n_457) );
INVx2_ASAP7_75t_SL g458 ( .A(n_393), .Y(n_458) );
NOR2xp67_ASAP7_75t_L g459 ( .A(n_393), .B(n_17), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_383), .B(n_420), .Y(n_460) );
OR2x6_ASAP7_75t_L g461 ( .A(n_382), .B(n_361), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_402), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_384), .B(n_361), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_393), .B(n_354), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_404), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_414), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_383), .B(n_18), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_383), .B(n_291), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_414), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_393), .B(n_307), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_420), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_392), .B(n_18), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_395), .B(n_19), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_379), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_395), .B(n_20), .Y(n_475) );
AND2x4_ASAP7_75t_L g476 ( .A(n_396), .B(n_61), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_397), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_396), .B(n_20), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_431), .B(n_412), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_448), .B(n_398), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_423), .B(n_404), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_460), .B(n_426), .Y(n_482) );
INVxp67_ASAP7_75t_L g483 ( .A(n_469), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_436), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_441), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_438), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_435), .B(n_412), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_453), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_454), .B(n_407), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_426), .B(n_403), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_450), .B(n_407), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_440), .B(n_403), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_452), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_450), .B(n_405), .Y(n_494) );
NAND3xp33_ASAP7_75t_L g495 ( .A(n_439), .B(n_413), .C(n_405), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_451), .B(n_390), .Y(n_496) );
NAND2x1p5_ASAP7_75t_L g497 ( .A(n_459), .B(n_418), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_451), .B(n_390), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_467), .B(n_390), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_437), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_440), .B(n_398), .Y(n_501) );
INVx1_ASAP7_75t_SL g502 ( .A(n_443), .Y(n_502) );
INVx2_ASAP7_75t_SL g503 ( .A(n_441), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_467), .B(n_410), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_452), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_471), .B(n_410), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_462), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_462), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_465), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_425), .B(n_387), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_465), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_425), .B(n_463), .Y(n_512) );
AND2x4_ASAP7_75t_L g513 ( .A(n_434), .B(n_413), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_445), .Y(n_514) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_424), .A2(n_399), .B(n_382), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_432), .B(n_397), .Y(n_516) );
INVxp67_ASAP7_75t_L g517 ( .A(n_445), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_422), .Y(n_518) );
INVx3_ASAP7_75t_L g519 ( .A(n_434), .Y(n_519) );
AND2x2_ASAP7_75t_SL g520 ( .A(n_464), .B(n_399), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_428), .B(n_397), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_446), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_428), .B(n_411), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_466), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_444), .A2(n_415), .B1(n_411), .B2(n_387), .Y(n_525) );
INVxp67_ASAP7_75t_SL g526 ( .A(n_437), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_449), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_442), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_447), .B(n_21), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_442), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_432), .B(n_411), .Y(n_531) );
NOR3xp33_ASAP7_75t_SL g532 ( .A(n_427), .B(n_419), .C(n_415), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_463), .B(n_418), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_433), .B(n_418), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_433), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_472), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_449), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_535), .B(n_456), .Y(n_538) );
NAND2x1_ASAP7_75t_L g539 ( .A(n_519), .B(n_457), .Y(n_539) );
OAI322xp33_ASAP7_75t_L g540 ( .A1(n_517), .A2(n_430), .A3(n_456), .B1(n_475), .B2(n_473), .C1(n_472), .C2(n_478), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_514), .B(n_468), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_512), .Y(n_542) );
AOI32xp33_ASAP7_75t_L g543 ( .A1(n_529), .A2(n_478), .A3(n_475), .B1(n_473), .B2(n_457), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_537), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_524), .Y(n_545) );
OAI21xp5_ASAP7_75t_L g546 ( .A1(n_529), .A2(n_476), .B(n_455), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_518), .B(n_468), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_482), .B(n_430), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_520), .A2(n_476), .B1(n_464), .B2(n_458), .Y(n_549) );
OAI21xp5_ASAP7_75t_L g550 ( .A1(n_525), .A2(n_476), .B(n_458), .Y(n_550) );
AOI21xp33_ASAP7_75t_L g551 ( .A1(n_481), .A2(n_461), .B(n_444), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_517), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_537), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_522), .B(n_477), .Y(n_554) );
O2A1O1Ixp33_ASAP7_75t_SL g555 ( .A1(n_485), .A2(n_477), .B(n_474), .C(n_464), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_490), .B(n_470), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_520), .A2(n_461), .B1(n_470), .B2(n_429), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_484), .Y(n_558) );
NAND2x1_ASAP7_75t_L g559 ( .A(n_519), .B(n_461), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_481), .A2(n_461), .B1(n_470), .B2(n_429), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_483), .B(n_474), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_483), .B(n_429), .Y(n_562) );
XOR2x2_ASAP7_75t_L g563 ( .A(n_504), .B(n_21), .Y(n_563) );
INVxp67_ASAP7_75t_L g564 ( .A(n_485), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_510), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_528), .B(n_22), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_536), .A2(n_174), .B1(n_159), .B2(n_273), .Y(n_567) );
AOI322xp5_ASAP7_75t_L g568 ( .A1(n_492), .A2(n_23), .A3(n_419), .B1(n_157), .B2(n_162), .C1(n_168), .C2(n_174), .Y(n_568) );
INVxp67_ASAP7_75t_SL g569 ( .A(n_526), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_501), .B(n_23), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_502), .B(n_480), .Y(n_571) );
OAI221xp5_ASAP7_75t_L g572 ( .A1(n_515), .A2(n_162), .B1(n_159), .B2(n_174), .C(n_273), .Y(n_572) );
OAI21xp5_ASAP7_75t_SL g573 ( .A1(n_513), .A2(n_305), .B(n_292), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_486), .Y(n_574) );
AO22x1_ASAP7_75t_L g575 ( .A1(n_519), .A2(n_284), .B1(n_26), .B2(n_27), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_488), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_479), .A2(n_159), .B1(n_174), .B2(n_284), .Y(n_577) );
INVx1_ASAP7_75t_SL g578 ( .A(n_503), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_503), .B(n_25), .Y(n_579) );
OAI21xp5_ASAP7_75t_L g580 ( .A1(n_525), .A2(n_320), .B(n_314), .Y(n_580) );
OAI21xp5_ASAP7_75t_SL g581 ( .A1(n_513), .A2(n_174), .B(n_159), .Y(n_581) );
O2A1O1Ixp33_ASAP7_75t_SL g582 ( .A1(n_499), .A2(n_28), .B(n_29), .C(n_33), .Y(n_582) );
OAI21xp5_ASAP7_75t_L g583 ( .A1(n_563), .A2(n_495), .B(n_532), .Y(n_583) );
OAI21xp33_ASAP7_75t_SL g584 ( .A1(n_569), .A2(n_526), .B(n_498), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_552), .B(n_530), .Y(n_585) );
NAND2x1_ASAP7_75t_L g586 ( .A(n_557), .B(n_513), .Y(n_586) );
OAI21xp5_ASAP7_75t_L g587 ( .A1(n_546), .A2(n_532), .B(n_497), .Y(n_587) );
INVx1_ASAP7_75t_SL g588 ( .A(n_578), .Y(n_588) );
INVxp67_ASAP7_75t_L g589 ( .A(n_570), .Y(n_589) );
AOI222xp33_ASAP7_75t_L g590 ( .A1(n_550), .A2(n_487), .B1(n_494), .B2(n_491), .C1(n_496), .C2(n_521), .Y(n_590) );
NOR2x1_ASAP7_75t_L g591 ( .A(n_581), .B(n_533), .Y(n_591) );
AOI222xp33_ASAP7_75t_L g592 ( .A1(n_566), .A2(n_523), .B1(n_516), .B2(n_531), .C1(n_493), .C2(n_508), .Y(n_592) );
NOR3xp33_ASAP7_75t_L g593 ( .A(n_551), .B(n_489), .C(n_505), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_571), .B(n_506), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_551), .A2(n_534), .B1(n_497), .B2(n_511), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_561), .Y(n_596) );
XNOR2xp5_ASAP7_75t_L g597 ( .A(n_549), .B(n_509), .Y(n_597) );
OAI222xp33_ASAP7_75t_L g598 ( .A1(n_543), .A2(n_507), .B1(n_500), .B2(n_527), .C1(n_43), .C2(n_44), .Y(n_598) );
OAI22xp33_ASAP7_75t_L g599 ( .A1(n_560), .A2(n_527), .B1(n_500), .B2(n_159), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_558), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_574), .Y(n_601) );
XOR2x2_ASAP7_75t_L g602 ( .A(n_542), .B(n_35), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g603 ( .A1(n_540), .A2(n_221), .B1(n_223), .B2(n_211), .C(n_208), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_547), .B(n_320), .Y(n_604) );
OAI21xp5_ASAP7_75t_SL g605 ( .A1(n_580), .A2(n_211), .B(n_41), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_576), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_545), .Y(n_607) );
INVxp67_ASAP7_75t_L g608 ( .A(n_562), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_547), .B(n_37), .Y(n_609) );
OAI22xp5_ASAP7_75t_SL g610 ( .A1(n_539), .A2(n_45), .B1(n_46), .B2(n_49), .Y(n_610) );
OAI222xp33_ASAP7_75t_L g611 ( .A1(n_586), .A2(n_559), .B1(n_548), .B2(n_562), .C1(n_564), .C2(n_538), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_583), .A2(n_538), .B1(n_565), .B2(n_541), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_600), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_589), .B(n_566), .Y(n_614) );
AOI21x1_ASAP7_75t_L g615 ( .A1(n_602), .A2(n_575), .B(n_579), .Y(n_615) );
OAI221xp5_ASAP7_75t_L g616 ( .A1(n_584), .A2(n_555), .B1(n_568), .B2(n_572), .C(n_573), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_596), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_601), .Y(n_618) );
OAI21xp5_ASAP7_75t_SL g619 ( .A1(n_598), .A2(n_556), .B(n_567), .Y(n_619) );
OAI21x1_ASAP7_75t_SL g620 ( .A1(n_587), .A2(n_553), .B(n_544), .Y(n_620) );
AOI322xp5_ASAP7_75t_L g621 ( .A1(n_593), .A2(n_541), .A3(n_554), .B1(n_577), .B2(n_582), .C1(n_58), .C2(n_59), .Y(n_621) );
OAI221xp5_ASAP7_75t_L g622 ( .A1(n_593), .A2(n_554), .B1(n_208), .B2(n_221), .C(n_57), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g623 ( .A1(n_598), .A2(n_314), .B(n_223), .Y(n_623) );
OAI22x1_ASAP7_75t_L g624 ( .A1(n_588), .A2(n_52), .B1(n_53), .B2(n_56), .Y(n_624) );
INVxp67_ASAP7_75t_L g625 ( .A(n_606), .Y(n_625) );
OAI21xp33_ASAP7_75t_L g626 ( .A1(n_590), .A2(n_221), .B(n_67), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_592), .A2(n_221), .B1(n_164), .B2(n_223), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_612), .A2(n_589), .B1(n_595), .B2(n_591), .Y(n_628) );
OAI22xp5_ASAP7_75t_SL g629 ( .A1(n_622), .A2(n_610), .B1(n_597), .B2(n_608), .Y(n_629) );
NAND4xp25_ASAP7_75t_L g630 ( .A(n_626), .B(n_603), .C(n_605), .D(n_609), .Y(n_630) );
NOR3xp33_ASAP7_75t_L g631 ( .A(n_615), .B(n_599), .C(n_608), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_617), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_619), .A2(n_607), .B1(n_585), .B2(n_594), .Y(n_633) );
INVx1_ASAP7_75t_SL g634 ( .A(n_624), .Y(n_634) );
AOI211xp5_ASAP7_75t_L g635 ( .A1(n_611), .A2(n_604), .B(n_221), .C(n_72), .Y(n_635) );
INVx2_ASAP7_75t_SL g636 ( .A(n_613), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_618), .Y(n_637) );
NOR2x1_ASAP7_75t_L g638 ( .A(n_634), .B(n_622), .Y(n_638) );
O2A1O1Ixp33_ASAP7_75t_L g639 ( .A1(n_631), .A2(n_620), .B(n_616), .C(n_614), .Y(n_639) );
INVx2_ASAP7_75t_SL g640 ( .A(n_636), .Y(n_640) );
OAI22xp5_ASAP7_75t_SL g641 ( .A1(n_629), .A2(n_616), .B1(n_627), .B2(n_625), .Y(n_641) );
AND3x4_ASAP7_75t_L g642 ( .A(n_633), .B(n_621), .C(n_623), .Y(n_642) );
NAND3xp33_ASAP7_75t_SL g643 ( .A(n_639), .B(n_635), .C(n_628), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_640), .Y(n_644) );
NAND4xp25_ASAP7_75t_L g645 ( .A(n_638), .B(n_630), .C(n_632), .D(n_637), .Y(n_645) );
OAI211xp5_ASAP7_75t_SL g646 ( .A1(n_644), .A2(n_641), .B(n_642), .C(n_73), .Y(n_646) );
AND3x1_ASAP7_75t_L g647 ( .A(n_643), .B(n_66), .C(n_71), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_646), .A2(n_645), .B1(n_223), .B2(n_164), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_647), .Y(n_649) );
O2A1O1Ixp33_ASAP7_75t_L g650 ( .A1(n_649), .A2(n_74), .B(n_76), .C(n_77), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_650), .A2(n_648), .B1(n_223), .B2(n_221), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_651), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_652), .A2(n_164), .B1(n_641), .B2(n_643), .Y(n_653) );
endmodule