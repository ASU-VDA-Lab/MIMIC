module fake_netlist_6_797_n_1587 (n_52, n_1, n_91, n_326, n_256, n_209, n_63, n_223, n_278, n_341, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_342, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_350, n_78, n_84, n_142, n_143, n_180, n_62, n_349, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_280, n_287, n_353, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_338, n_56, n_119, n_235, n_147, n_191, n_340, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_352, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_348, n_69, n_293, n_31, n_334, n_53, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1587);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_341;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_342;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_350;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_280;
input n_287;
input n_353;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_338;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_352;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_293;
input n_31;
input n_334;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1587;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_1575;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1558;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_513;
wire n_645;
wire n_1381;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_702;
wire n_1175;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_1033;
wire n_462;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1483;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1339;
wire n_537;
wire n_1427;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_1429;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_828;
wire n_607;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1586;
wire n_380;
wire n_1535;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1443;
wire n_1272;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_934;
wire n_482;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_1522;
wire n_548;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_799;
wire n_1548;
wire n_1155;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1373;
wire n_1292;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_712;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_1582;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1576;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1240;

INVx1_ASAP7_75t_SL g358 ( 
.A(n_121),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_142),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_192),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_55),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_270),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_10),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_25),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_297),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_274),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_331),
.Y(n_367)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_44),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_156),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_320),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_212),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_300),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_183),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_190),
.Y(n_374)
);

CKINVDCx14_ASAP7_75t_R g375 ( 
.A(n_165),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_132),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_23),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_68),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_110),
.Y(n_379)
);

BUFx8_ASAP7_75t_SL g380 ( 
.A(n_4),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_15),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_265),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_103),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_353),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_63),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_293),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_219),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_326),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_79),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_286),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_136),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_3),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_196),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_94),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_339),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_144),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_287),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_207),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_202),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_269),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_100),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_176),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_119),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_349),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_154),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_208),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_120),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_245),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_162),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_210),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_344),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_72),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_77),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_76),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_109),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_39),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_182),
.Y(n_417)
);

CKINVDCx11_ASAP7_75t_R g418 ( 
.A(n_347),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_312),
.Y(n_419)
);

CKINVDCx14_ASAP7_75t_R g420 ( 
.A(n_184),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_24),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_259),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_197),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_135),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_198),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_341),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_62),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_279),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_17),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_337),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_248),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_26),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_308),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_249),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_34),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_332),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_7),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_56),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_80),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_16),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_14),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_153),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_4),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_50),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_329),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_168),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_113),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_125),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_240),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_348),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_31),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_350),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_108),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_48),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_138),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_216),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_73),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_114),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_67),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_284),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_2),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_34),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_241),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_123),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_317),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_14),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_75),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_36),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_8),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_281),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_346),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_86),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_351),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_129),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_28),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_84),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_7),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_230),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_278),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_36),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_340),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_316),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_252),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_134),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_272),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_276),
.Y(n_486)
);

INVx2_ASAP7_75t_SL g487 ( 
.A(n_345),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_28),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_33),
.Y(n_489)
);

BUFx8_ASAP7_75t_SL g490 ( 
.A(n_49),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_239),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_146),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_53),
.Y(n_493)
);

BUFx10_ASAP7_75t_L g494 ( 
.A(n_2),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_26),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_23),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_47),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_228),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_65),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_158),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_127),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_315),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_199),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_30),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_310),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_37),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_32),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_319),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_311),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_163),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_131),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_222),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_140),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_203),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_253),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_17),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_223),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_47),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_18),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_98),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_10),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_231),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_35),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_321),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_71),
.Y(n_525)
);

BUFx2_ASAP7_75t_SL g526 ( 
.A(n_33),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_188),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_236),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_21),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_101),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_266),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_357),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_37),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_354),
.Y(n_534)
);

CKINVDCx14_ASAP7_75t_R g535 ( 
.A(n_8),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_145),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_149),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_25),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_260),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_81),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_232),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_186),
.Y(n_542)
);

BUFx10_ASAP7_75t_L g543 ( 
.A(n_24),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_247),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_296),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_338),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_227),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_234),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_6),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_96),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_469),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_469),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_469),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_469),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_380),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_506),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_396),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_428),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_506),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_506),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_490),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_506),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_429),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_440),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_437),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_459),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_418),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_464),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_359),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_365),
.Y(n_570)
);

CKINVDCx16_ASAP7_75t_R g571 ( 
.A(n_370),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_451),
.Y(n_572)
);

CKINVDCx16_ASAP7_75t_R g573 ( 
.A(n_368),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_371),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_462),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_482),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_494),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_468),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_521),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_523),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_499),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_533),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_367),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_368),
.B(n_0),
.Y(n_584)
);

NOR2xp67_ASAP7_75t_L g585 ( 
.A(n_453),
.B(n_0),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_549),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_367),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_535),
.B(n_1),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_466),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_361),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_372),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_395),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_395),
.Y(n_593)
);

INVxp67_ASAP7_75t_SL g594 ( 
.A(n_402),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_412),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_412),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_360),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_362),
.Y(n_598)
);

INVxp67_ASAP7_75t_L g599 ( 
.A(n_494),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_366),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_535),
.B(n_1),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_453),
.B(n_3),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_376),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_378),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_379),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_385),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_388),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_391),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_397),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_398),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_373),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_406),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_408),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_537),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_374),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_382),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_363),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_383),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_410),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_413),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_503),
.B(n_5),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_384),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_386),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_414),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_387),
.Y(n_625)
);

NOR2xp67_ASAP7_75t_L g626 ( 
.A(n_363),
.B(n_5),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_390),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_475),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_475),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_415),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_422),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_393),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_364),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_394),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_358),
.B(n_399),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_433),
.Y(n_636)
);

INVxp67_ASAP7_75t_SL g637 ( 
.A(n_438),
.Y(n_637)
);

CKINVDCx20_ASAP7_75t_R g638 ( 
.A(n_539),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_400),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_494),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_375),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_401),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_375),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_420),
.Y(n_644)
);

HB1xp67_ASAP7_75t_L g645 ( 
.A(n_377),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_477),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_488),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_455),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_488),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_456),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_403),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_457),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_381),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_463),
.Y(n_654)
);

CKINVDCx20_ASAP7_75t_R g655 ( 
.A(n_480),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_472),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_474),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_404),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_478),
.Y(n_659)
);

INVxp67_ASAP7_75t_SL g660 ( 
.A(n_481),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_511),
.B(n_6),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_405),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_409),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_411),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_483),
.Y(n_665)
);

INVxp67_ASAP7_75t_L g666 ( 
.A(n_543),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_486),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_417),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_551),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_552),
.Y(n_670)
);

HB1xp67_ASAP7_75t_L g671 ( 
.A(n_590),
.Y(n_671)
);

XOR2xp5_ASAP7_75t_L g672 ( 
.A(n_557),
.B(n_419),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_635),
.B(n_389),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_602),
.B(n_487),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_633),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_553),
.Y(n_676)
);

BUFx2_ASAP7_75t_L g677 ( 
.A(n_569),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_583),
.B(n_369),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_554),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_573),
.B(n_543),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_556),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_559),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_560),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_562),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_617),
.Y(n_685)
);

NAND2xp33_ASAP7_75t_L g686 ( 
.A(n_601),
.B(n_392),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_617),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_597),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_598),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_583),
.Y(n_690)
);

NOR2x1_ASAP7_75t_L g691 ( 
.A(n_585),
.B(n_491),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_635),
.B(n_543),
.Y(n_692)
);

INVx3_ASAP7_75t_L g693 ( 
.A(n_628),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_600),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_603),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_628),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_570),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_629),
.Y(n_698)
);

INVxp67_ASAP7_75t_L g699 ( 
.A(n_645),
.Y(n_699)
);

CKINVDCx8_ASAP7_75t_R g700 ( 
.A(n_555),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_602),
.B(n_369),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_629),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_647),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_647),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_SL g705 ( 
.A(n_641),
.B(n_416),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_604),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_605),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_649),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_606),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_637),
.B(n_550),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_649),
.Y(n_711)
);

INVx5_ASAP7_75t_L g712 ( 
.A(n_571),
.Y(n_712)
);

INVx1_ASAP7_75t_SL g713 ( 
.A(n_589),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_607),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_608),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_609),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_610),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_660),
.B(n_407),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_563),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_612),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_565),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_584),
.B(n_421),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_572),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_653),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_575),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_613),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_578),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_579),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_580),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_619),
.B(n_423),
.Y(n_730)
);

OAI21x1_ASAP7_75t_L g731 ( 
.A1(n_620),
.A2(n_425),
.B(n_407),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_624),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_584),
.B(n_432),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_630),
.B(n_424),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_582),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_588),
.B(n_594),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_586),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_631),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_636),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_648),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_650),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_652),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_654),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_656),
.B(n_426),
.Y(n_744)
);

NAND2x1p5_ASAP7_75t_L g745 ( 
.A(n_588),
.B(n_498),
.Y(n_745)
);

OA21x2_ASAP7_75t_L g746 ( 
.A1(n_657),
.A2(n_436),
.B(n_425),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_659),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_665),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_667),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_587),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_592),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_593),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_595),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_596),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_621),
.B(n_427),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_621),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_626),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_661),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_574),
.Y(n_759)
);

INVx1_ASAP7_75t_SL g760 ( 
.A(n_589),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_736),
.A2(n_663),
.B1(n_664),
.B2(n_643),
.Y(n_761)
);

AND2x6_ASAP7_75t_L g762 ( 
.A(n_701),
.B(n_436),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_690),
.B(n_508),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_673),
.B(n_591),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_756),
.B(n_611),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_703),
.Y(n_766)
);

INVx4_ASAP7_75t_SL g767 ( 
.A(n_680),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_703),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_703),
.Y(n_769)
);

INVx1_ASAP7_75t_SL g770 ( 
.A(n_713),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_740),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_673),
.B(n_615),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_690),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_678),
.B(n_513),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_688),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_756),
.B(n_616),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_692),
.B(n_577),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_678),
.B(n_514),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_689),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_756),
.B(n_618),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_SL g781 ( 
.A(n_697),
.B(n_561),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_669),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_756),
.B(n_755),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_759),
.B(n_622),
.Y(n_784)
);

BUFx3_ASAP7_75t_L g785 ( 
.A(n_751),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_703),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_755),
.B(n_623),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_694),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_679),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_695),
.Y(n_790)
);

AND2x6_ASAP7_75t_L g791 ( 
.A(n_701),
.B(n_450),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_710),
.B(n_625),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_706),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_707),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_709),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_710),
.B(n_627),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_679),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_679),
.Y(n_798)
);

AND2x2_ASAP7_75t_SL g799 ( 
.A(n_677),
.B(n_661),
.Y(n_799)
);

INVx4_ASAP7_75t_L g800 ( 
.A(n_740),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_740),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_714),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_679),
.Y(n_803)
);

BUFx8_ASAP7_75t_SL g804 ( 
.A(n_700),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_674),
.B(n_736),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_699),
.B(n_632),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_683),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_745),
.B(n_634),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_712),
.B(n_639),
.Y(n_809)
);

BUFx10_ASAP7_75t_L g810 ( 
.A(n_718),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_745),
.B(n_642),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_715),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_758),
.B(n_651),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_740),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_683),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_699),
.B(n_658),
.Y(n_816)
);

AND2x6_ASAP7_75t_L g817 ( 
.A(n_691),
.B(n_450),
.Y(n_817)
);

INVx4_ASAP7_75t_L g818 ( 
.A(n_741),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_712),
.B(n_662),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_683),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_692),
.B(n_668),
.Y(n_821)
);

INVxp67_ASAP7_75t_L g822 ( 
.A(n_671),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_683),
.Y(n_823)
);

AND2x6_ASAP7_75t_L g824 ( 
.A(n_718),
.B(n_473),
.Y(n_824)
);

INVx4_ASAP7_75t_L g825 ( 
.A(n_741),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_730),
.B(n_430),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_684),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_671),
.B(n_599),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_670),
.Y(n_829)
);

INVx4_ASAP7_75t_L g830 ( 
.A(n_741),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_721),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_730),
.B(n_431),
.Y(n_832)
);

BUFx10_ASAP7_75t_L g833 ( 
.A(n_757),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_712),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_734),
.B(n_434),
.Y(n_835)
);

NAND2xp33_ASAP7_75t_L g836 ( 
.A(n_734),
.B(n_439),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_676),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_681),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_744),
.B(n_442),
.Y(n_839)
);

AND2x6_ASAP7_75t_L g840 ( 
.A(n_752),
.B(n_473),
.Y(n_840)
);

BUFx4f_ASAP7_75t_L g841 ( 
.A(n_721),
.Y(n_841)
);

INVx1_ASAP7_75t_SL g842 ( 
.A(n_760),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_722),
.B(n_644),
.Y(n_843)
);

BUFx3_ASAP7_75t_L g844 ( 
.A(n_712),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_682),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_716),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_717),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_741),
.Y(n_848)
);

INVx8_ASAP7_75t_L g849 ( 
.A(n_721),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_827),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_783),
.B(n_744),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_782),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_805),
.A2(n_733),
.B(n_686),
.C(n_731),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_762),
.B(n_733),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_813),
.B(n_675),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_787),
.A2(n_566),
.B1(n_568),
.B2(n_558),
.Y(n_856)
);

NAND2x1p5_ASAP7_75t_L g857 ( 
.A(n_834),
.B(n_725),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_782),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_775),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_762),
.B(n_686),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_829),
.Y(n_861)
);

AO22x2_ASAP7_75t_L g862 ( 
.A1(n_777),
.A2(n_772),
.B1(n_764),
.B2(n_828),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_779),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_806),
.B(n_675),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_762),
.B(n_750),
.Y(n_865)
);

AO22x2_ASAP7_75t_L g866 ( 
.A1(n_822),
.A2(n_672),
.B1(n_526),
.B2(n_666),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_837),
.Y(n_867)
);

AO22x2_ASAP7_75t_L g868 ( 
.A1(n_770),
.A2(n_640),
.B1(n_525),
.B2(n_546),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_804),
.Y(n_869)
);

OAI221xp5_ASAP7_75t_L g870 ( 
.A1(n_821),
.A2(n_732),
.B1(n_742),
.B2(n_738),
.C(n_726),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_842),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_788),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_762),
.B(n_750),
.Y(n_873)
);

AO22x2_ASAP7_75t_L g874 ( 
.A1(n_767),
.A2(n_525),
.B1(n_546),
.B2(n_527),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_776),
.A2(n_705),
.B1(n_581),
.B2(n_614),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_765),
.Y(n_876)
);

AO22x2_ASAP7_75t_L g877 ( 
.A1(n_767),
.A2(n_536),
.B1(n_548),
.B2(n_515),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_790),
.Y(n_878)
);

OAI221xp5_ASAP7_75t_L g879 ( 
.A1(n_780),
.A2(n_748),
.B1(n_743),
.B2(n_564),
.C(n_753),
.Y(n_879)
);

AO22x2_ASAP7_75t_L g880 ( 
.A1(n_774),
.A2(n_778),
.B1(n_811),
.B2(n_808),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_773),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_810),
.B(n_724),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_810),
.B(n_724),
.Y(n_883)
);

BUFx8_ASAP7_75t_L g884 ( 
.A(n_844),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_793),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_791),
.B(n_754),
.Y(n_886)
);

AO22x2_ASAP7_75t_L g887 ( 
.A1(n_774),
.A2(n_655),
.B1(n_646),
.B2(n_12),
.Y(n_887)
);

NOR2xp67_ASAP7_75t_L g888 ( 
.A(n_761),
.B(n_567),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_794),
.Y(n_889)
);

AO22x2_ASAP7_75t_L g890 ( 
.A1(n_778),
.A2(n_655),
.B1(n_646),
.B2(n_12),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_795),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_838),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_816),
.Y(n_893)
);

INVxp67_ASAP7_75t_SL g894 ( 
.A(n_771),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_845),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_792),
.B(n_705),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_802),
.Y(n_897)
);

BUFx8_ASAP7_75t_L g898 ( 
.A(n_812),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_846),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_785),
.B(n_847),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_843),
.A2(n_638),
.B1(n_576),
.B2(n_446),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_791),
.A2(n_447),
.B1(n_448),
.B2(n_445),
.Y(n_902)
);

OR2x6_ASAP7_75t_L g903 ( 
.A(n_809),
.B(n_819),
.Y(n_903)
);

INVxp67_ASAP7_75t_L g904 ( 
.A(n_833),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_763),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_833),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_766),
.Y(n_907)
);

HB1xp67_ASAP7_75t_L g908 ( 
.A(n_763),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_768),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_769),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_786),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_796),
.Y(n_912)
);

AO22x2_ASAP7_75t_L g913 ( 
.A1(n_799),
.A2(n_13),
.B1(n_9),
.B2(n_11),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_791),
.B(n_754),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_831),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_831),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_791),
.B(n_747),
.Y(n_917)
);

NAND2x1p5_ASAP7_75t_L g918 ( 
.A(n_841),
.B(n_725),
.Y(n_918)
);

NAND2x1_ASAP7_75t_L g919 ( 
.A(n_824),
.B(n_746),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_826),
.B(n_747),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_803),
.Y(n_921)
);

AO22x2_ASAP7_75t_L g922 ( 
.A1(n_832),
.A2(n_13),
.B1(n_9),
.B2(n_11),
.Y(n_922)
);

NAND2x1p5_ASAP7_75t_L g923 ( 
.A(n_841),
.B(n_749),
.Y(n_923)
);

OAI221xp5_ASAP7_75t_L g924 ( 
.A1(n_835),
.A2(n_720),
.B1(n_739),
.B2(n_727),
.C(n_728),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_807),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_784),
.B(n_749),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_789),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_815),
.B(n_719),
.Y(n_928)
);

AO22x2_ASAP7_75t_L g929 ( 
.A1(n_839),
.A2(n_18),
.B1(n_15),
.B2(n_16),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_824),
.B(n_747),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_820),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_800),
.B(n_729),
.Y(n_932)
);

AO22x2_ASAP7_75t_L g933 ( 
.A1(n_781),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_933)
);

INVxp67_ASAP7_75t_L g934 ( 
.A(n_817),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_817),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_789),
.Y(n_936)
);

NAND2x1p5_ASAP7_75t_L g937 ( 
.A(n_800),
.B(n_735),
.Y(n_937)
);

HAxp5_ASAP7_75t_SL g938 ( 
.A(n_817),
.B(n_435),
.CON(n_938),
.SN(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_824),
.B(n_747),
.Y(n_939)
);

OAI221xp5_ASAP7_75t_L g940 ( 
.A1(n_836),
.A2(n_720),
.B1(n_737),
.B2(n_444),
.C(n_454),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_797),
.Y(n_941)
);

OAI221xp5_ASAP7_75t_L g942 ( 
.A1(n_818),
.A2(n_461),
.B1(n_489),
.B2(n_443),
.C(n_441),
.Y(n_942)
);

NAND2x1p5_ASAP7_75t_L g943 ( 
.A(n_818),
.B(n_693),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_824),
.Y(n_944)
);

NAND2x1p5_ASAP7_75t_L g945 ( 
.A(n_825),
.B(n_693),
.Y(n_945)
);

AO22x2_ASAP7_75t_L g946 ( 
.A1(n_825),
.A2(n_22),
.B1(n_19),
.B2(n_20),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_771),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_797),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_851),
.B(n_830),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_893),
.B(n_926),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_876),
.B(n_771),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_864),
.B(n_855),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_871),
.B(n_896),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_852),
.B(n_801),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_882),
.B(n_801),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_858),
.B(n_801),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_883),
.B(n_854),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_920),
.B(n_814),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_900),
.B(n_906),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_859),
.B(n_814),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_905),
.B(n_814),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_875),
.B(n_848),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_912),
.B(n_848),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_932),
.B(n_848),
.Y(n_964)
);

NAND2xp33_ASAP7_75t_SL g965 ( 
.A(n_935),
.B(n_449),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_863),
.B(n_849),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_872),
.B(n_849),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_878),
.B(n_721),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_885),
.B(n_723),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_889),
.B(n_723),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_891),
.B(n_798),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_897),
.B(n_723),
.Y(n_972)
);

NAND2xp33_ASAP7_75t_SL g973 ( 
.A(n_908),
.B(n_452),
.Y(n_973)
);

NAND2xp33_ASAP7_75t_SL g974 ( 
.A(n_860),
.B(n_458),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_899),
.B(n_798),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_904),
.B(n_723),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_947),
.B(n_460),
.Y(n_977)
);

NAND2xp33_ASAP7_75t_SL g978 ( 
.A(n_881),
.B(n_465),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_853),
.B(n_823),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_947),
.B(n_467),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_861),
.B(n_823),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_928),
.B(n_470),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_850),
.B(n_817),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_867),
.B(n_471),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_892),
.B(n_476),
.Y(n_985)
);

NAND2xp33_ASAP7_75t_SL g986 ( 
.A(n_938),
.B(n_479),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_895),
.B(n_484),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_901),
.B(n_685),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_902),
.B(n_856),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_934),
.B(n_865),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_873),
.B(n_485),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_886),
.B(n_914),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_862),
.B(n_840),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_862),
.B(n_840),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_918),
.B(n_492),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_880),
.B(n_840),
.Y(n_996)
);

NAND2xp33_ASAP7_75t_SL g997 ( 
.A(n_944),
.B(n_500),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_923),
.B(n_501),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_917),
.B(n_888),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_930),
.B(n_502),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_939),
.B(n_505),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_857),
.B(n_509),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_937),
.B(n_510),
.Y(n_1003)
);

NAND2xp33_ASAP7_75t_SL g1004 ( 
.A(n_869),
.B(n_512),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_903),
.B(n_687),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_927),
.B(n_517),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_880),
.B(n_840),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_894),
.B(n_702),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_936),
.B(n_520),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_941),
.B(n_948),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_915),
.B(n_522),
.Y(n_1011)
);

NAND2xp33_ASAP7_75t_SL g1012 ( 
.A(n_919),
.B(n_524),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_916),
.B(n_528),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_921),
.B(n_530),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_925),
.B(n_531),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_931),
.B(n_532),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_868),
.B(n_887),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_903),
.B(n_708),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_943),
.B(n_534),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_945),
.B(n_540),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_909),
.B(n_711),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_910),
.B(n_541),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_911),
.B(n_542),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_907),
.B(n_544),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_884),
.B(n_545),
.Y(n_1025)
);

NAND2xp33_ASAP7_75t_SL g1026 ( 
.A(n_919),
.B(n_547),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_898),
.B(n_698),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_870),
.B(n_698),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_940),
.B(n_704),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_942),
.B(n_704),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_979),
.A2(n_992),
.B(n_990),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_949),
.A2(n_746),
.B(n_924),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_950),
.B(n_868),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_952),
.B(n_887),
.Y(n_1034)
);

NAND2x1_ASAP7_75t_L g1035 ( 
.A(n_981),
.B(n_874),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_954),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_953),
.B(n_696),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_989),
.A2(n_879),
.B(n_495),
.C(n_496),
.Y(n_1038)
);

INVx4_ASAP7_75t_L g1039 ( 
.A(n_961),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_957),
.B(n_877),
.Y(n_1040)
);

NOR4xp25_ASAP7_75t_L g1041 ( 
.A(n_1017),
.B(n_913),
.C(n_933),
.D(n_890),
.Y(n_1041)
);

NOR3xp33_ASAP7_75t_SL g1042 ( 
.A(n_986),
.B(n_963),
.C(n_978),
.Y(n_1042)
);

AO22x2_ASAP7_75t_L g1043 ( 
.A1(n_993),
.A2(n_913),
.B1(n_946),
.B2(n_933),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_994),
.A2(n_497),
.B(n_504),
.C(n_493),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_958),
.A2(n_877),
.B(n_696),
.Y(n_1045)
);

BUFx2_ASAP7_75t_L g1046 ( 
.A(n_1005),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_983),
.A2(n_516),
.B(n_507),
.Y(n_1047)
);

AOI221x1_ASAP7_75t_L g1048 ( 
.A1(n_996),
.A2(n_929),
.B1(n_922),
.B2(n_946),
.C(n_866),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_999),
.A2(n_929),
.B(n_922),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_991),
.A2(n_866),
.B(n_890),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_L g1051 ( 
.A1(n_956),
.A2(n_58),
.B(n_57),
.Y(n_1051)
);

NAND2xp33_ASAP7_75t_L g1052 ( 
.A(n_1007),
.B(n_518),
.Y(n_1052)
);

NOR3xp33_ASAP7_75t_L g1053 ( 
.A(n_959),
.B(n_529),
.C(n_519),
.Y(n_1053)
);

HB1xp67_ASAP7_75t_L g1054 ( 
.A(n_951),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_964),
.A2(n_60),
.B(n_59),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_1005),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_1029),
.A2(n_538),
.B(n_64),
.Y(n_1057)
);

AO21x1_ASAP7_75t_L g1058 ( 
.A1(n_974),
.A2(n_22),
.B(n_27),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_1018),
.Y(n_1059)
);

OA21x2_ASAP7_75t_L g1060 ( 
.A1(n_971),
.A2(n_66),
.B(n_61),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_988),
.B(n_27),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_1000),
.A2(n_70),
.B(n_69),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_975),
.A2(n_78),
.B(n_74),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_L g1064 ( 
.A1(n_1010),
.A2(n_83),
.B(n_82),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_962),
.B(n_29),
.Y(n_1065)
);

INVx2_ASAP7_75t_SL g1066 ( 
.A(n_1018),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_955),
.B(n_29),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_961),
.B(n_30),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_960),
.B(n_31),
.Y(n_1069)
);

AOI21x1_ASAP7_75t_L g1070 ( 
.A1(n_1001),
.A2(n_1030),
.B(n_1013),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_965),
.A2(n_32),
.B(n_35),
.C(n_38),
.Y(n_1071)
);

OA21x2_ASAP7_75t_L g1072 ( 
.A1(n_1028),
.A2(n_87),
.B(n_85),
.Y(n_1072)
);

AO21x2_ASAP7_75t_L g1073 ( 
.A1(n_995),
.A2(n_89),
.B(n_88),
.Y(n_1073)
);

AO21x2_ASAP7_75t_L g1074 ( 
.A1(n_998),
.A2(n_91),
.B(n_90),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_1008),
.A2(n_93),
.B(n_92),
.Y(n_1075)
);

INVx2_ASAP7_75t_SL g1076 ( 
.A(n_1021),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1012),
.A2(n_97),
.B(n_95),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_968),
.A2(n_102),
.B(n_99),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_1026),
.A2(n_105),
.B(n_104),
.Y(n_1079)
);

NAND3xp33_ASAP7_75t_L g1080 ( 
.A(n_973),
.B(n_38),
.C(n_39),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1021),
.B(n_40),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_1004),
.Y(n_1082)
);

BUFx12f_ASAP7_75t_L g1083 ( 
.A(n_981),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_966),
.B(n_40),
.Y(n_1084)
);

AO31x2_ASAP7_75t_L g1085 ( 
.A1(n_997),
.A2(n_41),
.A3(n_42),
.B(n_43),
.Y(n_1085)
);

INVxp67_ASAP7_75t_L g1086 ( 
.A(n_982),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_969),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_967),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_1027),
.Y(n_1089)
);

NAND2xp33_ASAP7_75t_L g1090 ( 
.A(n_1003),
.B(n_106),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_1014),
.A2(n_41),
.B(n_42),
.C(n_43),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_976),
.A2(n_44),
.B(n_45),
.C(n_46),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_1015),
.A2(n_45),
.B(n_46),
.C(n_48),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1016),
.B(n_49),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_970),
.A2(n_972),
.B(n_1019),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_1011),
.A2(n_235),
.B1(n_356),
.B2(n_355),
.Y(n_1096)
);

OAI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_1022),
.A2(n_111),
.B(n_107),
.Y(n_1097)
);

AOI21x1_ASAP7_75t_L g1098 ( 
.A1(n_1006),
.A2(n_115),
.B(n_112),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1020),
.A2(n_117),
.B(n_116),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_1009),
.A2(n_122),
.B(n_118),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_1002),
.B(n_124),
.Y(n_1101)
);

CKINVDCx20_ASAP7_75t_R g1102 ( 
.A(n_1046),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1036),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1054),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1087),
.Y(n_1105)
);

CKINVDCx11_ASAP7_75t_R g1106 ( 
.A(n_1083),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_1059),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_1031),
.A2(n_1024),
.B(n_1023),
.Y(n_1108)
);

AOI22x1_ASAP7_75t_L g1109 ( 
.A1(n_1057),
.A2(n_980),
.B1(n_977),
.B2(n_985),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_1065),
.A2(n_987),
.B1(n_984),
.B2(n_1025),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_1064),
.A2(n_128),
.B(n_126),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1061),
.B(n_50),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_1070),
.A2(n_133),
.B(n_130),
.Y(n_1113)
);

INVxp67_ASAP7_75t_SL g1114 ( 
.A(n_1068),
.Y(n_1114)
);

AO21x1_ASAP7_75t_L g1115 ( 
.A1(n_1049),
.A2(n_51),
.B(n_52),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1081),
.Y(n_1116)
);

AO21x2_ASAP7_75t_L g1117 ( 
.A1(n_1032),
.A2(n_139),
.B(n_137),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1090),
.A2(n_143),
.B(n_141),
.Y(n_1118)
);

AO21x2_ASAP7_75t_L g1119 ( 
.A1(n_1045),
.A2(n_148),
.B(n_147),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1033),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_1095),
.A2(n_151),
.B(n_150),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_1078),
.A2(n_255),
.B(n_352),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1069),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_1089),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1076),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_SL g1126 ( 
.A(n_1039),
.B(n_51),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1040),
.Y(n_1127)
);

NOR2xp67_ASAP7_75t_L g1128 ( 
.A(n_1086),
.B(n_152),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1084),
.Y(n_1129)
);

INVxp67_ASAP7_75t_SL g1130 ( 
.A(n_1039),
.Y(n_1130)
);

OR2x6_ASAP7_75t_L g1131 ( 
.A(n_1035),
.B(n_1088),
.Y(n_1131)
);

AO32x2_ASAP7_75t_L g1132 ( 
.A1(n_1048),
.A2(n_52),
.A3(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1066),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_1088),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1094),
.Y(n_1135)
);

AOI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1037),
.A2(n_258),
.B(n_155),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_SL g1137 ( 
.A1(n_1097),
.A2(n_261),
.B(n_157),
.Y(n_1137)
);

OR2x6_ASAP7_75t_L g1138 ( 
.A(n_1088),
.B(n_159),
.Y(n_1138)
);

HB1xp67_ASAP7_75t_L g1139 ( 
.A(n_1056),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_1063),
.A2(n_262),
.B(n_160),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1051),
.A2(n_263),
.B(n_161),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1067),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1072),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1075),
.A2(n_264),
.B(n_164),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_1056),
.Y(n_1145)
);

INVx1_ASAP7_75t_SL g1146 ( 
.A(n_1034),
.Y(n_1146)
);

INVx1_ASAP7_75t_SL g1147 ( 
.A(n_1056),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1072),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_1082),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_1100),
.A2(n_267),
.B(n_166),
.Y(n_1150)
);

OA21x2_ASAP7_75t_L g1151 ( 
.A1(n_1077),
.A2(n_268),
.B(n_167),
.Y(n_1151)
);

AO21x2_ASAP7_75t_L g1152 ( 
.A1(n_1079),
.A2(n_271),
.B(n_169),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1043),
.B(n_54),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1098),
.A2(n_170),
.B(n_171),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1043),
.Y(n_1155)
);

INVx4_ASAP7_75t_L g1156 ( 
.A(n_1073),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_1085),
.Y(n_1157)
);

OA21x2_ASAP7_75t_L g1158 ( 
.A1(n_1044),
.A2(n_172),
.B(n_173),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1050),
.A2(n_174),
.B1(n_175),
.B2(n_177),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1073),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1041),
.B(n_178),
.Y(n_1161)
);

NAND2x1p5_ASAP7_75t_L g1162 ( 
.A(n_1101),
.B(n_179),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1062),
.A2(n_180),
.B(n_181),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1085),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_1080),
.A2(n_185),
.B1(n_187),
.B2(n_189),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1074),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_1042),
.Y(n_1167)
);

OAI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1038),
.A2(n_191),
.B(n_193),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1085),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1092),
.Y(n_1170)
);

NAND2x1p5_ASAP7_75t_L g1171 ( 
.A(n_1060),
.B(n_194),
.Y(n_1171)
);

OAI22xp33_ASAP7_75t_SL g1172 ( 
.A1(n_1047),
.A2(n_195),
.B1(n_200),
.B2(n_201),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1074),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_1096),
.Y(n_1174)
);

INVx6_ASAP7_75t_L g1175 ( 
.A(n_1053),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1103),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1105),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1123),
.B(n_1091),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1146),
.B(n_1114),
.Y(n_1179)
);

INVx4_ASAP7_75t_L g1180 ( 
.A(n_1131),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1143),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_1131),
.B(n_1139),
.Y(n_1182)
);

AO21x2_ASAP7_75t_L g1183 ( 
.A1(n_1164),
.A2(n_1052),
.B(n_1058),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1148),
.Y(n_1184)
);

HB1xp67_ASAP7_75t_L g1185 ( 
.A(n_1104),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1146),
.B(n_1114),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1155),
.B(n_1093),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1127),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1113),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1120),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1169),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1142),
.B(n_1071),
.Y(n_1192)
);

OR2x6_ASAP7_75t_L g1193 ( 
.A(n_1138),
.B(n_1099),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1129),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1135),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1157),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_1131),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1157),
.Y(n_1198)
);

NAND2x1p5_ASAP7_75t_L g1199 ( 
.A(n_1158),
.B(n_1121),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1116),
.B(n_1060),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_1161),
.B(n_1112),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1112),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1153),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_1102),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1171),
.Y(n_1205)
);

INVxp67_ASAP7_75t_L g1206 ( 
.A(n_1149),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1153),
.Y(n_1207)
);

OR2x2_ASAP7_75t_L g1208 ( 
.A(n_1161),
.B(n_1055),
.Y(n_1208)
);

INVxp67_ASAP7_75t_SL g1209 ( 
.A(n_1130),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1171),
.Y(n_1210)
);

BUFx2_ASAP7_75t_L g1211 ( 
.A(n_1130),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1139),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1144),
.A2(n_204),
.B(n_205),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1115),
.Y(n_1214)
);

INVx4_ASAP7_75t_L g1215 ( 
.A(n_1107),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1133),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1117),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1117),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1132),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_1163),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1154),
.Y(n_1221)
);

INVx1_ASAP7_75t_SL g1222 ( 
.A(n_1124),
.Y(n_1222)
);

HB1xp67_ASAP7_75t_L g1223 ( 
.A(n_1134),
.Y(n_1223)
);

AO21x2_ASAP7_75t_L g1224 ( 
.A1(n_1160),
.A2(n_206),
.B(n_209),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1151),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1140),
.A2(n_211),
.B(n_213),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1141),
.A2(n_214),
.B(n_215),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1151),
.Y(n_1228)
);

AOI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1166),
.A2(n_217),
.B(n_218),
.Y(n_1229)
);

INVx2_ASAP7_75t_SL g1230 ( 
.A(n_1145),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1132),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1132),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1174),
.A2(n_220),
.B1(n_221),
.B2(n_224),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1173),
.Y(n_1234)
);

INVx2_ASAP7_75t_SL g1235 ( 
.A(n_1134),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1125),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1111),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1170),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1136),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1122),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1108),
.Y(n_1241)
);

A2O1A1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1168),
.A2(n_225),
.B(n_226),
.C(n_229),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1147),
.Y(n_1243)
);

OAI221xp5_ASAP7_75t_L g1244 ( 
.A1(n_1110),
.A2(n_233),
.B1(n_237),
.B2(n_238),
.C(n_242),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1138),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1150),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1138),
.B(n_243),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1147),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1158),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1126),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1202),
.B(n_1167),
.Y(n_1251)
);

OR2x6_ASAP7_75t_L g1252 ( 
.A(n_1247),
.B(n_1197),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_1204),
.B(n_1128),
.Y(n_1253)
);

OR2x6_ASAP7_75t_L g1254 ( 
.A(n_1247),
.B(n_1175),
.Y(n_1254)
);

NAND2xp33_ASAP7_75t_R g1255 ( 
.A(n_1247),
.B(n_1168),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1204),
.B(n_1118),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_1215),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1179),
.B(n_1126),
.Y(n_1258)
);

NAND2xp33_ASAP7_75t_R g1259 ( 
.A(n_1245),
.B(n_1118),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_1201),
.B(n_1172),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1215),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1182),
.B(n_1152),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_R g1263 ( 
.A(n_1230),
.B(n_1106),
.Y(n_1263)
);

NAND2xp33_ASAP7_75t_R g1264 ( 
.A(n_1201),
.B(n_1175),
.Y(n_1264)
);

NAND2xp33_ASAP7_75t_R g1265 ( 
.A(n_1192),
.B(n_244),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1179),
.B(n_1162),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1211),
.Y(n_1267)
);

INVxp67_ASAP7_75t_L g1268 ( 
.A(n_1185),
.Y(n_1268)
);

NAND2xp33_ASAP7_75t_SL g1269 ( 
.A(n_1215),
.B(n_1159),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1176),
.Y(n_1270)
);

NAND2xp33_ASAP7_75t_R g1271 ( 
.A(n_1192),
.B(n_246),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_1182),
.B(n_1152),
.Y(n_1272)
);

AND2x2_ASAP7_75t_SL g1273 ( 
.A(n_1197),
.B(n_1165),
.Y(n_1273)
);

CKINVDCx9p33_ASAP7_75t_R g1274 ( 
.A(n_1211),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_1230),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1182),
.B(n_1119),
.Y(n_1276)
);

INVx2_ASAP7_75t_SL g1277 ( 
.A(n_1243),
.Y(n_1277)
);

INVxp67_ASAP7_75t_L g1278 ( 
.A(n_1236),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1222),
.Y(n_1279)
);

INVxp67_ASAP7_75t_L g1280 ( 
.A(n_1216),
.Y(n_1280)
);

NAND2xp33_ASAP7_75t_R g1281 ( 
.A(n_1186),
.B(n_250),
.Y(n_1281)
);

OR2x6_ASAP7_75t_L g1282 ( 
.A(n_1197),
.B(n_1162),
.Y(n_1282)
);

XOR2x2_ASAP7_75t_SL g1283 ( 
.A(n_1194),
.B(n_1172),
.Y(n_1283)
);

OR2x2_ASAP7_75t_L g1284 ( 
.A(n_1203),
.B(n_1119),
.Y(n_1284)
);

NAND2xp33_ASAP7_75t_R g1285 ( 
.A(n_1186),
.B(n_251),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1195),
.B(n_1109),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1207),
.B(n_254),
.Y(n_1287)
);

CKINVDCx16_ASAP7_75t_R g1288 ( 
.A(n_1223),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1176),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1250),
.B(n_256),
.Y(n_1290)
);

INVxp67_ASAP7_75t_L g1291 ( 
.A(n_1206),
.Y(n_1291)
);

NAND2xp33_ASAP7_75t_R g1292 ( 
.A(n_1193),
.B(n_257),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1178),
.B(n_1137),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1177),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1180),
.B(n_1156),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_R g1296 ( 
.A(n_1197),
.B(n_1235),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1188),
.Y(n_1297)
);

INVxp67_ASAP7_75t_L g1298 ( 
.A(n_1248),
.Y(n_1298)
);

BUFx10_ASAP7_75t_L g1299 ( 
.A(n_1212),
.Y(n_1299)
);

OR2x6_ASAP7_75t_L g1300 ( 
.A(n_1197),
.B(n_1156),
.Y(n_1300)
);

INVxp67_ASAP7_75t_L g1301 ( 
.A(n_1235),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1180),
.B(n_1209),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1190),
.Y(n_1303)
);

NAND2xp33_ASAP7_75t_R g1304 ( 
.A(n_1193),
.B(n_273),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1187),
.B(n_275),
.Y(n_1305)
);

INVx2_ASAP7_75t_SL g1306 ( 
.A(n_1180),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1191),
.Y(n_1307)
);

XNOR2xp5_ASAP7_75t_L g1308 ( 
.A(n_1187),
.B(n_277),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_1193),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1238),
.Y(n_1310)
);

INVxp67_ASAP7_75t_L g1311 ( 
.A(n_1200),
.Y(n_1311)
);

INVxp67_ASAP7_75t_L g1312 ( 
.A(n_1200),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1214),
.B(n_280),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_R g1314 ( 
.A(n_1208),
.B(n_1229),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_SL g1315 ( 
.A(n_1242),
.B(n_282),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1193),
.B(n_283),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1208),
.B(n_285),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1191),
.Y(n_1318)
);

BUFx10_ASAP7_75t_L g1319 ( 
.A(n_1196),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_SL g1320 ( 
.A(n_1242),
.B(n_288),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_R g1321 ( 
.A(n_1229),
.B(n_289),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1198),
.Y(n_1322)
);

INVxp67_ASAP7_75t_L g1323 ( 
.A(n_1183),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_1233),
.Y(n_1324)
);

XNOR2xp5_ASAP7_75t_L g1325 ( 
.A(n_1244),
.B(n_290),
.Y(n_1325)
);

AND2x4_ASAP7_75t_L g1326 ( 
.A(n_1205),
.B(n_291),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1307),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1311),
.B(n_1234),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1322),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1312),
.B(n_1318),
.Y(n_1330)
);

AOI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1255),
.A2(n_1183),
.B1(n_1205),
.B2(n_1210),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1267),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1309),
.B(n_1210),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1309),
.B(n_1234),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1294),
.B(n_1219),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1268),
.B(n_1181),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1270),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1297),
.B(n_1303),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1267),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1289),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1310),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1284),
.Y(n_1342)
);

OR2x2_ASAP7_75t_L g1343 ( 
.A(n_1323),
.B(n_1249),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1258),
.B(n_1231),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1319),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1288),
.B(n_1249),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1298),
.B(n_1181),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1286),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1272),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1280),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1272),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1277),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1278),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1262),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1299),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1276),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1266),
.B(n_1184),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_1274),
.Y(n_1358)
);

OR2x2_ASAP7_75t_L g1359 ( 
.A(n_1260),
.B(n_1217),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1300),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_1302),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1300),
.B(n_1232),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1302),
.Y(n_1363)
);

BUFx4f_ASAP7_75t_SL g1364 ( 
.A(n_1279),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1315),
.A2(n_1183),
.B1(n_1220),
.B2(n_1224),
.Y(n_1365)
);

OR2x2_ASAP7_75t_L g1366 ( 
.A(n_1293),
.B(n_1218),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1295),
.Y(n_1367)
);

INVxp67_ASAP7_75t_L g1368 ( 
.A(n_1251),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1301),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1256),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1305),
.B(n_1184),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1264),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1316),
.B(n_1217),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1259),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1320),
.A2(n_1220),
.B1(n_1224),
.B2(n_1239),
.Y(n_1375)
);

INVx2_ASAP7_75t_SL g1376 ( 
.A(n_1257),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1317),
.B(n_1218),
.Y(n_1377)
);

AND2x4_ASAP7_75t_L g1378 ( 
.A(n_1306),
.B(n_1241),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1261),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1252),
.B(n_1241),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1252),
.B(n_1225),
.Y(n_1381)
);

INVx8_ASAP7_75t_L g1382 ( 
.A(n_1254),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1282),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1254),
.B(n_1225),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1275),
.Y(n_1385)
);

OAI33xp33_ASAP7_75t_L g1386 ( 
.A1(n_1348),
.A2(n_1291),
.A3(n_1324),
.B1(n_1283),
.B2(n_1228),
.B3(n_1265),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1338),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1344),
.B(n_1314),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1349),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1332),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1372),
.A2(n_1308),
.B1(n_1325),
.B2(n_1273),
.Y(n_1391)
);

BUFx6f_ASAP7_75t_L g1392 ( 
.A(n_1382),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1342),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1344),
.B(n_1228),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1368),
.B(n_1253),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1329),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1338),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1337),
.Y(n_1398)
);

NAND3xp33_ASAP7_75t_L g1399 ( 
.A(n_1374),
.B(n_1285),
.C(n_1281),
.Y(n_1399)
);

AO21x2_ASAP7_75t_L g1400 ( 
.A1(n_1331),
.A2(n_1321),
.B(n_1348),
.Y(n_1400)
);

AOI221xp5_ASAP7_75t_L g1401 ( 
.A1(n_1350),
.A2(n_1308),
.B1(n_1269),
.B2(n_1287),
.C(n_1325),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1349),
.B(n_1224),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1337),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1353),
.B(n_1341),
.Y(n_1404)
);

AND2x4_ASAP7_75t_SL g1405 ( 
.A(n_1352),
.B(n_1345),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1379),
.Y(n_1406)
);

BUFx2_ASAP7_75t_L g1407 ( 
.A(n_1361),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1327),
.Y(n_1408)
);

INVx1_ASAP7_75t_SL g1409 ( 
.A(n_1364),
.Y(n_1409)
);

INVx1_ASAP7_75t_SL g1410 ( 
.A(n_1379),
.Y(n_1410)
);

INVx1_ASAP7_75t_SL g1411 ( 
.A(n_1361),
.Y(n_1411)
);

INVx1_ASAP7_75t_SL g1412 ( 
.A(n_1358),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1351),
.B(n_1199),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1357),
.B(n_1313),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1351),
.B(n_1282),
.Y(n_1415)
);

INVxp67_ASAP7_75t_L g1416 ( 
.A(n_1369),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1390),
.B(n_1342),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1407),
.B(n_1354),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1396),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1396),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1393),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1411),
.B(n_1346),
.Y(n_1422)
);

NOR2x1_ASAP7_75t_L g1423 ( 
.A(n_1399),
.B(n_1358),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1403),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1398),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1407),
.B(n_1346),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1398),
.Y(n_1427)
);

INVxp33_ASAP7_75t_L g1428 ( 
.A(n_1392),
.Y(n_1428)
);

AND2x4_ASAP7_75t_SL g1429 ( 
.A(n_1392),
.B(n_1345),
.Y(n_1429)
);

INVx1_ASAP7_75t_SL g1430 ( 
.A(n_1410),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1408),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1408),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1416),
.B(n_1377),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1388),
.B(n_1354),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1387),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1388),
.B(n_1356),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1397),
.B(n_1356),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1404),
.B(n_1366),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1389),
.B(n_1362),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1394),
.Y(n_1440)
);

OAI221xp5_ASAP7_75t_L g1441 ( 
.A1(n_1423),
.A2(n_1391),
.B1(n_1401),
.B2(n_1412),
.C(n_1271),
.Y(n_1441)
);

OAI221xp5_ASAP7_75t_L g1442 ( 
.A1(n_1433),
.A2(n_1395),
.B1(n_1304),
.B2(n_1292),
.C(n_1355),
.Y(n_1442)
);

OAI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1428),
.A2(n_1392),
.B1(n_1382),
.B2(n_1370),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_SL g1444 ( 
.A(n_1438),
.B(n_1392),
.Y(n_1444)
);

AOI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1430),
.A2(n_1386),
.B1(n_1400),
.B2(n_1383),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1421),
.B(n_1405),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1422),
.B(n_1405),
.Y(n_1447)
);

AO221x2_ASAP7_75t_L g1448 ( 
.A1(n_1419),
.A2(n_1385),
.B1(n_1383),
.B2(n_1400),
.C(n_1360),
.Y(n_1448)
);

BUFx2_ASAP7_75t_L g1449 ( 
.A(n_1426),
.Y(n_1449)
);

AOI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1428),
.A2(n_1400),
.B1(n_1392),
.B2(n_1382),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1429),
.Y(n_1451)
);

NOR4xp25_ASAP7_75t_SL g1452 ( 
.A(n_1420),
.B(n_1360),
.C(n_1339),
.D(n_1340),
.Y(n_1452)
);

INVx3_ASAP7_75t_L g1453 ( 
.A(n_1429),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1437),
.B(n_1414),
.Y(n_1454)
);

INVx3_ASAP7_75t_SL g1455 ( 
.A(n_1417),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1434),
.B(n_1406),
.Y(n_1456)
);

NOR4xp25_ASAP7_75t_SL g1457 ( 
.A(n_1424),
.B(n_1363),
.C(n_1406),
.D(n_1296),
.Y(n_1457)
);

AO221x2_ASAP7_75t_L g1458 ( 
.A1(n_1435),
.A2(n_1425),
.B1(n_1432),
.B2(n_1431),
.C(n_1367),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1449),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1445),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1458),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1454),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1455),
.B(n_1437),
.Y(n_1463)
);

INVxp67_ASAP7_75t_L g1464 ( 
.A(n_1441),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1448),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1446),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1444),
.B(n_1447),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1448),
.Y(n_1468)
);

BUFx3_ASAP7_75t_L g1469 ( 
.A(n_1451),
.Y(n_1469)
);

NOR3x1_ASAP7_75t_L g1470 ( 
.A(n_1442),
.B(n_1376),
.C(n_1336),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1453),
.B(n_1439),
.Y(n_1471)
);

INVx1_ASAP7_75t_SL g1472 ( 
.A(n_1456),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1450),
.B(n_1436),
.Y(n_1473)
);

AOI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1443),
.A2(n_1415),
.B1(n_1382),
.B2(n_1376),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1452),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1457),
.B(n_1439),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1455),
.B(n_1418),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1441),
.A2(n_1365),
.B1(n_1290),
.B2(n_1359),
.Y(n_1478)
);

INVxp67_ASAP7_75t_L g1479 ( 
.A(n_1459),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1462),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1463),
.Y(n_1481)
);

AOI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1460),
.A2(n_1415),
.B1(n_1362),
.B2(n_1367),
.Y(n_1482)
);

INVx1_ASAP7_75t_SL g1483 ( 
.A(n_1469),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1477),
.B(n_1418),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1472),
.B(n_1440),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1466),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1460),
.B(n_1440),
.Y(n_1487)
);

NAND2x1_ASAP7_75t_L g1488 ( 
.A(n_1476),
.B(n_1389),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1469),
.B(n_1409),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1461),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_SL g1491 ( 
.A(n_1483),
.B(n_1464),
.Y(n_1491)
);

INVx1_ASAP7_75t_SL g1492 ( 
.A(n_1483),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1485),
.B(n_1461),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1489),
.B(n_1464),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1486),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1490),
.B(n_1468),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1488),
.Y(n_1497)
);

AND2x2_ASAP7_75t_SL g1498 ( 
.A(n_1481),
.B(n_1470),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1480),
.Y(n_1499)
);

OAI21xp33_ASAP7_75t_L g1500 ( 
.A1(n_1479),
.A2(n_1478),
.B(n_1465),
.Y(n_1500)
);

BUFx4f_ASAP7_75t_SL g1501 ( 
.A(n_1492),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_1491),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1495),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1499),
.Y(n_1504)
);

CKINVDCx20_ASAP7_75t_R g1505 ( 
.A(n_1494),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1496),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1493),
.Y(n_1507)
);

NOR3xp33_ASAP7_75t_L g1508 ( 
.A(n_1502),
.B(n_1500),
.C(n_1497),
.Y(n_1508)
);

AOI211x1_ASAP7_75t_SL g1509 ( 
.A1(n_1501),
.A2(n_1487),
.B(n_1465),
.C(n_1475),
.Y(n_1509)
);

AOI221xp5_ASAP7_75t_L g1510 ( 
.A1(n_1506),
.A2(n_1500),
.B1(n_1478),
.B2(n_1497),
.C(n_1498),
.Y(n_1510)
);

NOR2x1_ASAP7_75t_L g1511 ( 
.A(n_1505),
.B(n_1467),
.Y(n_1511)
);

O2A1O1Ixp33_ASAP7_75t_L g1512 ( 
.A1(n_1503),
.A2(n_1473),
.B(n_1484),
.C(n_1471),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_SL g1513 ( 
.A(n_1507),
.B(n_1482),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1504),
.B(n_1474),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1501),
.Y(n_1515)
);

A2O1A1Ixp33_ASAP7_75t_L g1516 ( 
.A1(n_1502),
.A2(n_1359),
.B(n_1375),
.C(n_1415),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1502),
.B(n_1427),
.Y(n_1517)
);

OAI211xp5_ASAP7_75t_L g1518 ( 
.A1(n_1510),
.A2(n_1263),
.B(n_1347),
.C(n_1366),
.Y(n_1518)
);

OAI211xp5_ASAP7_75t_L g1519 ( 
.A1(n_1508),
.A2(n_1384),
.B(n_1427),
.C(n_1377),
.Y(n_1519)
);

AOI221xp5_ASAP7_75t_L g1520 ( 
.A1(n_1513),
.A2(n_1389),
.B1(n_1334),
.B2(n_1330),
.C(n_1378),
.Y(n_1520)
);

AOI221xp5_ASAP7_75t_L g1521 ( 
.A1(n_1515),
.A2(n_1334),
.B1(n_1330),
.B2(n_1378),
.C(n_1333),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1517),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1511),
.B(n_1333),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1514),
.A2(n_1384),
.B1(n_1343),
.B2(n_1333),
.Y(n_1524)
);

AOI221xp5_ASAP7_75t_L g1525 ( 
.A1(n_1512),
.A2(n_1334),
.B1(n_1378),
.B2(n_1381),
.C(n_1327),
.Y(n_1525)
);

AOI211xp5_ASAP7_75t_L g1526 ( 
.A1(n_1516),
.A2(n_1326),
.B(n_1381),
.C(n_1226),
.Y(n_1526)
);

AOI211xp5_ASAP7_75t_L g1527 ( 
.A1(n_1509),
.A2(n_1227),
.B(n_1226),
.C(n_1213),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1523),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1522),
.B(n_1394),
.Y(n_1529)
);

NOR2x1_ASAP7_75t_L g1530 ( 
.A(n_1518),
.B(n_1343),
.Y(n_1530)
);

XNOR2xp5_ASAP7_75t_L g1531 ( 
.A(n_1519),
.B(n_1371),
.Y(n_1531)
);

CKINVDCx16_ASAP7_75t_R g1532 ( 
.A(n_1524),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1521),
.Y(n_1533)
);

OAI221xp5_ASAP7_75t_L g1534 ( 
.A1(n_1526),
.A2(n_1525),
.B1(n_1520),
.B2(n_1527),
.C(n_1199),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_SL g1535 ( 
.A1(n_1523),
.A2(n_1402),
.B1(n_1373),
.B2(n_1413),
.Y(n_1535)
);

AND3x4_ASAP7_75t_L g1536 ( 
.A(n_1523),
.B(n_1189),
.C(n_1239),
.Y(n_1536)
);

NOR2xp33_ASAP7_75t_R g1537 ( 
.A(n_1532),
.B(n_292),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_R g1538 ( 
.A(n_1528),
.B(n_294),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_R g1539 ( 
.A(n_1533),
.B(n_295),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_R g1540 ( 
.A(n_1531),
.B(n_298),
.Y(n_1540)
);

NAND2xp33_ASAP7_75t_SL g1541 ( 
.A(n_1536),
.B(n_1373),
.Y(n_1541)
);

NAND2xp33_ASAP7_75t_SL g1542 ( 
.A(n_1529),
.B(n_1371),
.Y(n_1542)
);

NOR3xp33_ASAP7_75t_SL g1543 ( 
.A(n_1534),
.B(n_299),
.C(n_301),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_R g1544 ( 
.A(n_1530),
.B(n_302),
.Y(n_1544)
);

NAND2xp33_ASAP7_75t_SL g1545 ( 
.A(n_1535),
.B(n_1402),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_R g1546 ( 
.A(n_1532),
.B(n_303),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1532),
.B(n_1413),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1537),
.B(n_1335),
.Y(n_1548)
);

NAND3xp33_ASAP7_75t_SL g1549 ( 
.A(n_1546),
.B(n_1199),
.C(n_1380),
.Y(n_1549)
);

NAND4xp25_ASAP7_75t_L g1550 ( 
.A(n_1547),
.B(n_1380),
.C(n_1328),
.D(n_1220),
.Y(n_1550)
);

XOR2x1_ASAP7_75t_L g1551 ( 
.A(n_1538),
.B(n_304),
.Y(n_1551)
);

NAND3xp33_ASAP7_75t_SL g1552 ( 
.A(n_1544),
.B(n_1328),
.C(n_1221),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1543),
.A2(n_1540),
.B1(n_1539),
.B2(n_1545),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1542),
.B(n_1335),
.Y(n_1554)
);

AND3x2_ASAP7_75t_L g1555 ( 
.A(n_1541),
.B(n_305),
.C(n_306),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1547),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1547),
.Y(n_1557)
);

BUFx2_ASAP7_75t_L g1558 ( 
.A(n_1537),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1547),
.B(n_1227),
.Y(n_1559)
);

BUFx3_ASAP7_75t_L g1560 ( 
.A(n_1547),
.Y(n_1560)
);

HB1xp67_ASAP7_75t_L g1561 ( 
.A(n_1551),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1558),
.B(n_307),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1560),
.B(n_309),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1556),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1555),
.Y(n_1565)
);

INVx2_ASAP7_75t_SL g1566 ( 
.A(n_1557),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1548),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1553),
.Y(n_1568)
);

XNOR2xp5_ASAP7_75t_L g1569 ( 
.A(n_1552),
.B(n_1549),
.Y(n_1569)
);

OR4x1_ASAP7_75t_L g1570 ( 
.A(n_1550),
.B(n_313),
.C(n_314),
.D(n_318),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1561),
.Y(n_1571)
);

XNOR2xp5_ASAP7_75t_L g1572 ( 
.A(n_1569),
.B(n_1554),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1565),
.B(n_1566),
.Y(n_1573)
);

INVxp67_ASAP7_75t_SL g1574 ( 
.A(n_1563),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1564),
.A2(n_1559),
.B1(n_1189),
.B2(n_1221),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_SL g1576 ( 
.A1(n_1568),
.A2(n_1246),
.B1(n_1240),
.B2(n_1237),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1571),
.A2(n_1567),
.B1(n_1573),
.B2(n_1574),
.Y(n_1577)
);

AOI31xp33_ASAP7_75t_L g1578 ( 
.A1(n_1572),
.A2(n_1562),
.A3(n_1567),
.B(n_1570),
.Y(n_1578)
);

AOI31xp33_ASAP7_75t_L g1579 ( 
.A1(n_1575),
.A2(n_322),
.A3(n_323),
.B(n_324),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1577),
.B(n_1576),
.Y(n_1580)
);

OAI322xp33_ASAP7_75t_L g1581 ( 
.A1(n_1578),
.A2(n_1246),
.A3(n_1240),
.B1(n_1237),
.B2(n_330),
.C1(n_333),
.C2(n_334),
.Y(n_1581)
);

OR2x6_ASAP7_75t_L g1582 ( 
.A(n_1580),
.B(n_1579),
.Y(n_1582)
);

XNOR2xp5_ASAP7_75t_L g1583 ( 
.A(n_1581),
.B(n_325),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1582),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1583),
.Y(n_1585)
);

OAI221xp5_ASAP7_75t_R g1586 ( 
.A1(n_1584),
.A2(n_327),
.B1(n_328),
.B2(n_335),
.C(n_336),
.Y(n_1586)
);

AOI211xp5_ASAP7_75t_L g1587 ( 
.A1(n_1586),
.A2(n_1585),
.B(n_342),
.C(n_343),
.Y(n_1587)
);


endmodule