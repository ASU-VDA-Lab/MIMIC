module fake_jpeg_14016_n_235 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_235);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_235;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp33_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_54),
.Y(n_66)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_26),
.B(n_0),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_49),
.B(n_18),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_28),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_50),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_91)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_52),
.Y(n_80)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g97 ( 
.A(n_53),
.Y(n_97)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_57),
.Y(n_70)
);

BUFx4f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_56),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_59),
.Y(n_72)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_17),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_27),
.B(n_1),
.C(n_2),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_5),
.C(n_6),
.Y(n_92)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_62),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_21),
.B(n_15),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_32),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_33),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_81),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_30),
.B1(n_25),
.B2(n_23),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_67),
.A2(n_69),
.B1(n_86),
.B2(n_95),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_48),
.A2(n_30),
.B1(n_25),
.B2(n_23),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_L g110 ( 
.A1(n_73),
.A2(n_81),
.B(n_66),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_52),
.A2(n_37),
.B1(n_33),
.B2(n_31),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_74),
.A2(n_91),
.B1(n_58),
.B2(n_43),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_40),
.B(n_37),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_59),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_31),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_87),
.C(n_94),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_54),
.A2(n_35),
.B1(n_26),
.B2(n_29),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_84),
.A2(n_90),
.B1(n_68),
.B2(n_74),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_53),
.A2(n_32),
.B1(n_29),
.B2(n_21),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_1),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_38),
.A2(n_35),
.B1(n_3),
.B2(n_4),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_61),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_6),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_55),
.A2(n_8),
.B1(n_10),
.B2(n_14),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_44),
.A2(n_10),
.B1(n_47),
.B2(n_56),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_96),
.A2(n_56),
.B1(n_43),
.B2(n_42),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_72),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_100),
.B(n_102),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_101),
.A2(n_106),
.B1(n_71),
.B2(n_75),
.Y(n_134)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_121),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_104),
.B(n_117),
.Y(n_147)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_42),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_107),
.B(n_108),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_64),
.A2(n_46),
.B(n_83),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_119),
.B(n_128),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_110),
.B(n_120),
.Y(n_142)
);

BUFx4f_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_85),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_113),
.A2(n_75),
.B(n_71),
.Y(n_133)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

OR2x2_ASAP7_75t_SL g115 ( 
.A(n_94),
.B(n_92),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_118),
.Y(n_137)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_77),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_123),
.B(n_124),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_67),
.A2(n_75),
.B(n_80),
.C(n_78),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_125),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_78),
.B(n_79),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g129 ( 
.A(n_127),
.Y(n_129)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_SL g130 ( 
.A(n_115),
.B(n_75),
.C(n_79),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_146),
.C(n_139),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_149),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_101),
.A2(n_65),
.B1(n_89),
.B2(n_109),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_SL g163 ( 
.A1(n_141),
.A2(n_146),
.B(n_139),
.C(n_134),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_104),
.A2(n_89),
.B(n_99),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_L g172 ( 
.A1(n_143),
.A2(n_149),
.B(n_152),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_122),
.B1(n_124),
.B2(n_113),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_144),
.A2(n_148),
.B1(n_150),
.B2(n_137),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_108),
.A2(n_114),
.B(n_113),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_108),
.A2(n_99),
.B1(n_126),
.B2(n_105),
.Y(n_148)
);

AOI32xp33_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_123),
.A3(n_118),
.B1(n_111),
.B2(n_128),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_125),
.A2(n_112),
.B1(n_111),
.B2(n_116),
.Y(n_150)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_161),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_145),
.B(n_147),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_156),
.B(n_160),
.Y(n_183)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_158),
.A2(n_163),
.B(n_172),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_148),
.C(n_130),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_133),
.C(n_135),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_147),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_140),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_166),
.Y(n_185)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_164),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_137),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_167),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_142),
.B(n_145),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_169),
.A2(n_170),
.B1(n_136),
.B2(n_138),
.Y(n_188)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_141),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_135),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_173),
.B(n_132),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_142),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_174),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_191),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_190),
.C(n_173),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_154),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_186),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_168),
.A2(n_136),
.B1(n_138),
.B2(n_163),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_188),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_158),
.C(n_165),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_171),
.A2(n_163),
.B(n_168),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_194),
.C(n_197),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_190),
.B(n_163),
.C(n_167),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_157),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_198),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_163),
.C(n_164),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_161),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_179),
.C(n_184),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_177),
.C(n_176),
.Y(n_212)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_201),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_185),
.B(n_184),
.Y(n_202)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_202),
.Y(n_211)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_175),
.Y(n_203)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_203),
.Y(n_213)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_181),
.Y(n_204)
);

OA21x2_ASAP7_75t_SL g210 ( 
.A1(n_204),
.A2(n_186),
.B(n_181),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_179),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_209),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_191),
.Y(n_209)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_210),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_199),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_209),
.A2(n_177),
.B1(n_194),
.B2(n_197),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_217),
.Y(n_223)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_213),
.Y(n_216)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_216),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_212),
.A2(n_195),
.B(n_192),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_213),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_219),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_214),
.A2(n_205),
.B(n_177),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_222),
.A2(n_217),
.B(n_206),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_205),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_220),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_211),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_226),
.A2(n_227),
.B1(n_229),
.B2(n_223),
.Y(n_231)
);

BUFx24_ASAP7_75t_SL g230 ( 
.A(n_228),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_222),
.B(n_208),
.Y(n_229)
);

NAND3xp33_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_226),
.C(n_225),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_232),
.B(n_233),
.Y(n_234)
);

NOR4xp25_ASAP7_75t_L g233 ( 
.A(n_230),
.B(n_220),
.C(n_176),
.D(n_221),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_234),
.B(n_207),
.Y(n_235)
);


endmodule