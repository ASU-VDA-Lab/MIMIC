module fake_jpeg_26316_n_119 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_119);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_119;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_2),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_20),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_17),
.B1(n_37),
.B2(n_33),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_39),
.B1(n_14),
.B2(n_16),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_1),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_64),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_1),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_54),
.A2(n_51),
.B1(n_40),
.B2(n_49),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_70),
.B1(n_2),
.B2(n_3),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_50),
.Y(n_71)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_71),
.A2(n_46),
.B1(n_43),
.B2(n_44),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_75),
.A2(n_76),
.B1(n_4),
.B2(n_5),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_69),
.A2(n_46),
.B1(n_44),
.B2(n_42),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_67),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_83),
.Y(n_96)
);

AO21x1_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_50),
.B(n_3),
.Y(n_78)
);

AO21x1_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_82),
.B(n_6),
.Y(n_95)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_22),
.B1(n_32),
.B2(n_31),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_88),
.A2(n_87),
.B1(n_74),
.B2(n_81),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_95),
.B1(n_94),
.B2(n_96),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_93),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_21),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_79),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_78),
.B(n_88),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_100),
.A2(n_104),
.B(n_98),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_103),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_96),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_6),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_7),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_108),
.C(n_100),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_109),
.Y(n_110)
);

AOI322xp5_ASAP7_75t_L g112 ( 
.A1(n_110),
.A2(n_111),
.A3(n_99),
.B1(n_107),
.B2(n_9),
.C1(n_11),
.C2(n_12),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_27),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_24),
.C(n_30),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_19),
.C(n_23),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

MAJx2_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_28),
.C(n_29),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_117),
.B(n_38),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_7),
.Y(n_119)
);


endmodule