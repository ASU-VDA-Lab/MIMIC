module fake_jpeg_18703_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_20),
.B1(n_32),
.B2(n_27),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_48),
.A2(n_44),
.B1(n_20),
.B2(n_27),
.Y(n_96)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_28),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_50),
.B(n_21),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_30),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_54),
.A2(n_60),
.B(n_65),
.Y(n_90)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_17),
.Y(n_60)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_30),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_36),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_21),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_75),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_28),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_73),
.B(n_82),
.Y(n_114)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_76),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_45),
.Y(n_77)
);

AOI21xp33_ASAP7_75t_L g119 ( 
.A1(n_77),
.A2(n_33),
.B(n_23),
.Y(n_119)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_78),
.B(n_79),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_52),
.Y(n_79)
);

OAI32xp33_ASAP7_75t_L g80 ( 
.A1(n_57),
.A2(n_46),
.A3(n_22),
.B1(n_31),
.B2(n_34),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_98),
.Y(n_112)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_26),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_84),
.B(n_86),
.Y(n_136)
);

AOI32xp33_ASAP7_75t_L g85 ( 
.A1(n_60),
.A2(n_20),
.A3(n_46),
.B1(n_27),
.B2(n_32),
.Y(n_85)
);

AOI32xp33_ASAP7_75t_L g121 ( 
.A1(n_85),
.A2(n_67),
.A3(n_45),
.B1(n_43),
.B2(n_42),
.Y(n_121)
);

INVx5_ASAP7_75t_SL g86 ( 
.A(n_64),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_87),
.B(n_88),
.Y(n_137)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_89),
.B(n_93),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_L g91 ( 
.A1(n_58),
.A2(n_44),
.B1(n_46),
.B2(n_20),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_91),
.A2(n_100),
.B1(n_67),
.B2(n_33),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_32),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_56),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_96),
.A2(n_31),
.B1(n_35),
.B2(n_29),
.Y(n_138)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_26),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_47),
.A2(n_43),
.B1(n_42),
.B2(n_37),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_65),
.A2(n_27),
.B1(n_34),
.B2(n_22),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_109),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_54),
.B(n_34),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_107),
.A2(n_65),
.B(n_33),
.C(n_23),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_123),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_119),
.B(n_121),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_90),
.A2(n_0),
.B(n_1),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_69),
.B(n_63),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_80),
.A2(n_43),
.B1(n_42),
.B2(n_37),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_131),
.B1(n_100),
.B2(n_91),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_31),
.B1(n_86),
.B2(n_35),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_134),
.A2(n_90),
.B(n_77),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_141),
.A2(n_126),
.B(n_130),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_142),
.A2(n_150),
.B1(n_151),
.B2(n_155),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_112),
.A2(n_101),
.B1(n_87),
.B2(n_78),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_158),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_112),
.A2(n_88),
.B1(n_104),
.B2(n_106),
.Y(n_146)
);

MAJx2_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_77),
.C(n_83),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_147),
.A2(n_152),
.B(n_135),
.Y(n_191)
);

OAI32xp33_ASAP7_75t_L g148 ( 
.A1(n_113),
.A2(n_104),
.A3(n_29),
.B1(n_25),
.B2(n_16),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_149),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_113),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_108),
.B1(n_103),
.B2(n_95),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_131),
.A2(n_70),
.B1(n_95),
.B2(n_81),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_139),
.A2(n_70),
.B1(n_74),
.B2(n_16),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_118),
.B(n_71),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_153),
.B(n_161),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_125),
.A2(n_76),
.B1(n_25),
.B2(n_13),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_157),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_119),
.A2(n_25),
.B1(n_18),
.B2(n_24),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_122),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_117),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_124),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_168),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_118),
.B(n_25),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_162),
.A2(n_127),
.B1(n_132),
.B2(n_136),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_53),
.C(n_24),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_167),
.C(n_127),
.Y(n_180)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_114),
.B(n_30),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_136),
.Y(n_177)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_111),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_166),
.B(n_171),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_114),
.B(n_24),
.C(n_99),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_110),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_133),
.A2(n_16),
.B1(n_17),
.B2(n_13),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_169),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_196)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_111),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_176),
.A2(n_179),
.B1(n_194),
.B2(n_195),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_177),
.B(n_178),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_110),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_150),
.A2(n_128),
.B1(n_115),
.B2(n_133),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_163),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_117),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_181),
.B(n_183),
.Y(n_213)
);

AO22x1_ASAP7_75t_L g182 ( 
.A1(n_140),
.A2(n_128),
.B1(n_115),
.B2(n_129),
.Y(n_182)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_117),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_185),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_116),
.Y(n_186)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_126),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_187),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_164),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_188),
.B(n_193),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_189),
.A2(n_192),
.B(n_143),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_191),
.A2(n_196),
.B(n_6),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_154),
.A2(n_170),
.B(n_156),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_162),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_142),
.A2(n_135),
.B1(n_130),
.B2(n_129),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_151),
.A2(n_129),
.B1(n_24),
.B2(n_17),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_144),
.B(n_0),
.Y(n_199)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_146),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_202),
.B(n_2),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_155),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_203),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_157),
.B(n_2),
.Y(n_204)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_189),
.A2(n_154),
.B(n_170),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_205),
.A2(n_212),
.B(n_219),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_173),
.A2(n_170),
.B1(n_148),
.B2(n_152),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_206),
.A2(n_211),
.B1(n_194),
.B2(n_201),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_182),
.C(n_200),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_173),
.A2(n_171),
.B1(n_166),
.B2(n_147),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_217),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_216),
.A2(n_229),
.B1(n_199),
.B2(n_204),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_198),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_191),
.A2(n_4),
.B(n_5),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_186),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_223),
.Y(n_254)
);

INVxp67_ASAP7_75t_SL g223 ( 
.A(n_188),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_198),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_200),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_172),
.A2(n_9),
.B1(n_12),
.B2(n_11),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_225),
.A2(n_230),
.B1(n_199),
.B2(n_196),
.Y(n_240)
);

INVx3_ASAP7_75t_SL g226 ( 
.A(n_174),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_174),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_192),
.A2(n_4),
.B(n_6),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_227),
.A2(n_176),
.B(n_178),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_181),
.B(n_183),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_180),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_172),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_230)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_236),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_190),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_190),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_243),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_238),
.B(n_240),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_241),
.A2(n_252),
.B1(n_253),
.B2(n_209),
.Y(n_262)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_242),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_177),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_251),
.Y(n_266)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_182),
.C(n_184),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_246),
.B(n_247),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_214),
.B(n_175),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_221),
.Y(n_248)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_211),
.B(n_184),
.C(n_197),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_250),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_205),
.B(n_197),
.C(n_179),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_212),
.B(n_175),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_206),
.A2(n_195),
.B1(n_201),
.B2(n_203),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_210),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_255),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_254),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_257),
.B(n_258),
.Y(n_286)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_234),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_261),
.B(n_269),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_262),
.A2(n_268),
.B1(n_240),
.B2(n_222),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_253),
.A2(n_230),
.B1(n_225),
.B2(n_241),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_251),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_239),
.A2(n_220),
.B(n_207),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_271),
.A2(n_239),
.B(n_207),
.Y(n_280)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_249),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_237),
.Y(n_275)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_275),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_235),
.C(n_243),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_277),
.C(n_282),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_256),
.C(n_264),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_273),
.Y(n_278)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_278),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_236),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_283),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_280),
.A2(n_229),
.B(n_219),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_281),
.A2(n_257),
.B1(n_258),
.B2(n_222),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_246),
.C(n_244),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_250),
.Y(n_283)
);

INVxp33_ASAP7_75t_L g285 ( 
.A(n_273),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_289),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_267),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_218),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_261),
.A2(n_252),
.B1(n_209),
.B2(n_274),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_288),
.A2(n_265),
.B1(n_231),
.B2(n_218),
.Y(n_301)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_259),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_232),
.C(n_224),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_283),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_291),
.A2(n_292),
.B1(n_286),
.B2(n_285),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_290),
.A2(n_272),
.B1(n_270),
.B2(n_263),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_294),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_302),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_284),
.A2(n_265),
.B(n_231),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_300),
.B(n_297),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_287),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_279),
.B(n_227),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_302),
.C(n_282),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_308),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_277),
.C(n_276),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_307),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_293),
.A2(n_296),
.B1(n_303),
.B2(n_298),
.Y(n_306)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_306),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_311),
.A2(n_295),
.B1(n_13),
.B2(n_8),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_226),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_312),
.A2(n_226),
.B1(n_299),
.B2(n_216),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_315),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_295),
.C(n_7),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_309),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_312),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_319),
.B(n_320),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_309),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_322),
.A2(n_313),
.B(n_314),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_324),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_325),
.A2(n_323),
.B(n_321),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_326),
.B(n_315),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_310),
.C(n_6),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_8),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_8),
.B(n_327),
.Y(n_330)
);


endmodule