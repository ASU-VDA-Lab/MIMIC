module real_jpeg_3842_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_1),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_1),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_1),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_1),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_1),
.B(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_1),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_1),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_1),
.B(n_242),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_2),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_2),
.B(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_2),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_2),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_2),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_2),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_2),
.B(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_4),
.B(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_4),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_4),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_4),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_4),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_4),
.B(n_280),
.Y(n_279)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_6),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_6),
.Y(n_264)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_7),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_7),
.Y(n_96)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_9),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_9),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_9),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_9),
.B(n_101),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_9),
.B(n_179),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_10),
.Y(n_86)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_10),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_11),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_11),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_11),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_12),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g167 ( 
.A(n_12),
.B(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_13),
.Y(n_114)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_13),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_14),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_14),
.B(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_14),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_14),
.B(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_15),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_15),
.B(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_SL g166 ( 
.A(n_15),
.B(n_101),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_196),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_194),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_154),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_19),
.B(n_154),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_97),
.C(n_138),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_20),
.B(n_200),
.Y(n_199)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_20),
.Y(n_336)
);

FAx1_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_62),
.CI(n_79),
.CON(n_20),
.SN(n_20)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_21),
.B(n_62),
.C(n_79),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_38),
.C(n_52),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_22),
.B(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_33),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_24),
.B(n_29),
.C(n_33),
.Y(n_153)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_27),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_28),
.Y(n_273)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_36),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_37),
.Y(n_126)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_37),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_38),
.A2(n_52),
.B1(n_53),
.B2(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_38),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_43),
.C(n_49),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_39),
.A2(n_49),
.B1(n_173),
.B2(n_209),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_39),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

OR2x2_ASAP7_75t_SL g64 ( 
.A(n_40),
.B(n_65),
.Y(n_64)
);

OR2x2_ASAP7_75t_SL g162 ( 
.A(n_40),
.B(n_163),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_40),
.B(n_175),
.Y(n_174)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_43),
.B(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVx11_ASAP7_75t_L g239 ( 
.A(n_48),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_49),
.A2(n_173),
.B1(n_174),
.B2(n_176),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_49),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_50),
.Y(n_234)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_51),
.Y(n_220)
);

BUFx8_ASAP7_75t_L g298 ( 
.A(n_51),
.Y(n_298)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_58),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_54),
.A2(n_55),
.B1(n_58),
.B2(n_59),
.Y(n_221)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_57),
.Y(n_290)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_61),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_69),
.B2(n_70),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_64),
.B(n_71),
.C(n_76),
.Y(n_185)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_65),
.Y(n_217)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_67),
.Y(n_252)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_75),
.B1(n_76),
.B2(n_78),
.Y(n_70)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_71),
.A2(n_78),
.B1(n_122),
.B2(n_123),
.Y(n_258)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_78),
.B(n_122),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_88),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_80),
.A2(n_81),
.B(n_83),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_80),
.B(n_89),
.C(n_92),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_83),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_87),
.B(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_93),
.B(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_93),
.B(n_255),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_93),
.B(n_288),
.Y(n_287)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_97),
.B(n_138),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_117),
.C(n_119),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_98),
.A2(n_117),
.B1(n_118),
.B2(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_98),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_104),
.B2(n_116),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_105),
.C(n_110),
.Y(n_140)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_109),
.B1(n_110),
.B2(n_115),
.Y(n_104)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_114),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_114),
.Y(n_281)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_119),
.B(n_204),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_127),
.C(n_133),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_120),
.A2(n_121),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_127),
.A2(n_128),
.B1(n_133),
.B2(n_134),
.Y(n_326)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_132),
.Y(n_179)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_153),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_141),
.C(n_153),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_148),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_144),
.C(n_148),
.Y(n_159)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_147),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_180),
.B1(n_192),
.B2(n_193),
.Y(n_156)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_157),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_170),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_165),
.B2(n_169),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_177),
.B2(n_178),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_174),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_174),
.A2(n_176),
.B1(n_249),
.B2(n_250),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_176),
.B(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_180),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_225),
.B(n_334),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_199),
.B(n_201),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_206),
.C(n_222),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_202),
.A2(n_203),
.B1(n_331),
.B2(n_332),
.Y(n_330)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_206),
.B(n_222),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.C(n_221),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_207),
.B(n_318),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_210),
.B(n_221),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_215),
.C(n_218),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_211),
.A2(n_212),
.B1(n_215),
.B2(n_216),
.Y(n_245)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_218),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_218),
.Y(n_246)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_328),
.B(n_333),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_313),
.B(n_327),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_268),
.B(n_312),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_259),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_229),
.B(n_259),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_247),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_243),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_231),
.B(n_243),
.C(n_247),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_235),
.C(n_240),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_232),
.A2(n_233),
.B1(n_235),
.B2(n_236),
.Y(n_261)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_240),
.B(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_253),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_248),
.B(n_322),
.C(n_323),
.Y(n_321)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_258),
.Y(n_253)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_254),
.Y(n_322)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_258),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.C(n_267),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_260),
.B(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_262),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_262),
.A2(n_267),
.B1(n_304),
.B2(n_310),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_263),
.Y(n_302)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_264),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_265),
.Y(n_303)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_267),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_306),
.B(n_311),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_292),
.B(n_305),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_277),
.B(n_291),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_287),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_287),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_282),
.B(n_286),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_282),
.Y(n_286)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_286),
.A2(n_294),
.B1(n_299),
.B2(n_300),
.Y(n_293)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_286),
.Y(n_299)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx8_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_301),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_301),
.Y(n_305)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_294),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_295),
.A2(n_296),
.B(n_299),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_303),
.B(n_304),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_308),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_315),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_319),
.B2(n_320),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_321),
.C(n_324),
.Y(n_329)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_324),
.Y(n_320)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_330),
.Y(n_333)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_331),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);


endmodule