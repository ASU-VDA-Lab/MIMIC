module real_aes_1032_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_0), .B(n_140), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_1), .A2(n_149), .B(n_154), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_2), .B(n_820), .Y(n_819) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_3), .B(n_156), .Y(n_194) );
INVx1_ASAP7_75t_L g147 ( .A(n_4), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_5), .B(n_156), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_6), .B(n_166), .Y(n_570) );
INVx1_ASAP7_75t_L g550 ( .A(n_7), .Y(n_550) );
CKINVDCx16_ASAP7_75t_R g820 ( .A(n_8), .Y(n_820) );
CKINVDCx5p33_ASAP7_75t_R g516 ( .A(n_9), .Y(n_516) );
NAND2xp33_ASAP7_75t_L g183 ( .A(n_10), .B(n_158), .Y(n_183) );
INVx2_ASAP7_75t_L g137 ( .A(n_11), .Y(n_137) );
AOI221x1_ASAP7_75t_L g229 ( .A1(n_12), .A2(n_24), .B1(n_140), .B2(n_149), .C(n_230), .Y(n_229) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_13), .Y(n_111) );
NOR3xp33_ASAP7_75t_L g818 ( .A(n_13), .B(n_819), .C(n_821), .Y(n_818) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_14), .B(n_140), .Y(n_179) );
AO21x2_ASAP7_75t_L g176 ( .A1(n_15), .A2(n_177), .B(n_178), .Y(n_176) );
INVx1_ASAP7_75t_L g578 ( .A(n_16), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_17), .B(n_160), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_18), .B(n_156), .Y(n_170) );
AO21x1_ASAP7_75t_L g189 ( .A1(n_19), .A2(n_140), .B(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g115 ( .A(n_20), .Y(n_115) );
INVx1_ASAP7_75t_L g576 ( .A(n_21), .Y(n_576) );
INVx1_ASAP7_75t_SL g498 ( .A(n_22), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_23), .B(n_141), .Y(n_566) );
NAND2x1_ASAP7_75t_L g202 ( .A(n_25), .B(n_156), .Y(n_202) );
AOI33xp33_ASAP7_75t_L g536 ( .A1(n_26), .A2(n_54), .A3(n_481), .B1(n_486), .B2(n_537), .B3(n_538), .Y(n_536) );
NAND2x1_ASAP7_75t_L g221 ( .A(n_27), .B(n_158), .Y(n_221) );
INVx1_ASAP7_75t_L g509 ( .A(n_28), .Y(n_509) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_29), .A2(n_89), .B(n_137), .Y(n_136) );
OR2x2_ASAP7_75t_L g162 ( .A(n_29), .B(n_89), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_30), .B(n_489), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_31), .B(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_32), .B(n_156), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_33), .B(n_158), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_34), .A2(n_149), .B(n_210), .Y(n_209) );
AOI22xp5_ASAP7_75t_SL g797 ( .A1(n_35), .A2(n_798), .B1(n_804), .B2(n_805), .Y(n_797) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_35), .Y(n_804) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_36), .Y(n_823) );
AND2x2_ASAP7_75t_L g146 ( .A(n_37), .B(n_147), .Y(n_146) );
AND2x2_ASAP7_75t_L g150 ( .A(n_37), .B(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g480 ( .A(n_37), .Y(n_480) );
OR2x6_ASAP7_75t_L g113 ( .A(n_38), .B(n_114), .Y(n_113) );
INVxp67_ASAP7_75t_L g821 ( .A(n_38), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_39), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_40), .B(n_140), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_41), .B(n_489), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_42), .A2(n_135), .B1(n_166), .B2(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_43), .B(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_44), .B(n_141), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_45), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_46), .B(n_158), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_47), .B(n_177), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_48), .B(n_141), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_49), .A2(n_149), .B(n_220), .Y(n_219) );
CKINVDCx5p33_ASAP7_75t_R g563 ( .A(n_50), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g121 ( .A1(n_51), .A2(n_86), .B1(n_122), .B2(n_123), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_51), .Y(n_123) );
AOI22xp5_ASAP7_75t_L g800 ( .A1(n_52), .A2(n_81), .B1(n_801), .B2(n_802), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_52), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_53), .B(n_158), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_55), .B(n_141), .Y(n_527) );
INVx1_ASAP7_75t_L g143 ( .A(n_56), .Y(n_143) );
INVx1_ASAP7_75t_L g153 ( .A(n_56), .Y(n_153) );
AOI22xp5_ASAP7_75t_L g117 ( .A1(n_57), .A2(n_118), .B1(n_444), .B2(n_445), .Y(n_117) );
INVxp67_ASAP7_75t_L g445 ( .A(n_57), .Y(n_445) );
AND2x2_ASAP7_75t_L g528 ( .A(n_57), .B(n_160), .Y(n_528) );
AOI221xp5_ASAP7_75t_L g548 ( .A1(n_58), .A2(n_75), .B1(n_478), .B2(n_489), .C(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_59), .B(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_60), .B(n_156), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_61), .B(n_135), .Y(n_518) );
AOI21xp5_ASAP7_75t_SL g477 ( .A1(n_62), .A2(n_478), .B(n_483), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_63), .A2(n_149), .B(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g573 ( .A(n_64), .Y(n_573) );
AO21x1_ASAP7_75t_L g191 ( .A1(n_65), .A2(n_149), .B(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_66), .B(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_67), .B(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g526 ( .A(n_68), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_69), .B(n_140), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_70), .A2(n_478), .B(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g214 ( .A(n_71), .B(n_161), .Y(n_214) );
INVx1_ASAP7_75t_L g145 ( .A(n_72), .Y(n_145) );
INVx1_ASAP7_75t_L g151 ( .A(n_72), .Y(n_151) );
AND2x2_ASAP7_75t_L g225 ( .A(n_73), .B(n_134), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_74), .B(n_489), .Y(n_539) );
AND2x2_ASAP7_75t_L g500 ( .A(n_76), .B(n_134), .Y(n_500) );
INVx1_ASAP7_75t_L g574 ( .A(n_77), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_78), .A2(n_478), .B(n_497), .Y(n_496) );
OAI22xp5_ASAP7_75t_SL g119 ( .A1(n_79), .A2(n_120), .B1(n_121), .B2(n_124), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_79), .Y(n_124) );
A2O1A1Ixp33_ASAP7_75t_L g564 ( .A1(n_80), .A2(n_478), .B(n_531), .C(n_565), .Y(n_564) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_81), .Y(n_801) );
INVx1_ASAP7_75t_L g116 ( .A(n_82), .Y(n_116) );
AND2x2_ASAP7_75t_L g133 ( .A(n_83), .B(n_134), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_84), .B(n_140), .Y(n_172) );
AND2x2_ASAP7_75t_SL g475 ( .A(n_85), .B(n_134), .Y(n_475) );
INVx1_ASAP7_75t_L g122 ( .A(n_86), .Y(n_122) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_87), .A2(n_478), .B1(n_534), .B2(n_535), .Y(n_533) );
AND2x2_ASAP7_75t_L g190 ( .A(n_88), .B(n_166), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_90), .B(n_158), .Y(n_171) );
AND2x2_ASAP7_75t_L g206 ( .A(n_91), .B(n_134), .Y(n_206) );
INVx1_ASAP7_75t_L g484 ( .A(n_92), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_93), .B(n_156), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g798 ( .A1(n_94), .A2(n_799), .B1(n_800), .B2(n_803), .Y(n_798) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_94), .Y(n_799) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_95), .A2(n_149), .B(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_96), .B(n_158), .Y(n_231) );
AND2x2_ASAP7_75t_L g540 ( .A(n_97), .B(n_134), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_98), .B(n_156), .Y(n_155) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_99), .A2(n_507), .B(n_508), .C(n_511), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_100), .Y(n_812) );
BUFx2_ASAP7_75t_L g453 ( .A(n_101), .Y(n_453) );
BUFx2_ASAP7_75t_SL g457 ( .A(n_101), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_102), .A2(n_149), .B(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_103), .B(n_141), .Y(n_487) );
AOI21xp33_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_814), .B(n_822), .Y(n_104) );
OA22x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_449), .B1(n_454), .B2(n_458), .Y(n_105) );
OAI21x1_ASAP7_75t_SL g106 ( .A1(n_107), .A2(n_117), .B(n_446), .Y(n_106) );
BUFx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
BUFx3_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_L g448 ( .A(n_110), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
AND2x6_ASAP7_75t_SL g462 ( .A(n_111), .B(n_113), .Y(n_462) );
OR2x6_ASAP7_75t_SL g464 ( .A(n_111), .B(n_112), .Y(n_464) );
OR2x2_ASAP7_75t_L g813 ( .A(n_111), .B(n_113), .Y(n_813) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g817 ( .A(n_114), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
INVx1_ASAP7_75t_L g444 ( .A(n_118), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_125), .B1(n_442), .B2(n_443), .Y(n_118) );
INVx1_ASAP7_75t_L g442 ( .A(n_119), .Y(n_442) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g443 ( .A(n_125), .Y(n_443) );
INVx3_ASAP7_75t_L g809 ( .A(n_125), .Y(n_809) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_351), .Y(n_125) );
NOR4xp25_ASAP7_75t_L g126 ( .A(n_127), .B(n_269), .C(n_295), .D(n_335), .Y(n_126) );
OAI211xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_184), .B(n_215), .C(n_255), .Y(n_127) );
INVxp67_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_163), .Y(n_129) );
AND2x2_ASAP7_75t_L g422 ( .A(n_130), .B(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_131), .B(n_163), .Y(n_289) );
BUFx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g216 ( .A(n_132), .B(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_132), .B(n_242), .Y(n_241) );
INVx5_ASAP7_75t_L g275 ( .A(n_132), .Y(n_275) );
NOR2x1_ASAP7_75t_SL g317 ( .A(n_132), .B(n_164), .Y(n_317) );
AND2x2_ASAP7_75t_L g373 ( .A(n_132), .B(n_176), .Y(n_373) );
OR2x6_ASAP7_75t_L g132 ( .A(n_133), .B(n_138), .Y(n_132) );
INVx3_ASAP7_75t_L g205 ( .A(n_134), .Y(n_205) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_134), .A2(n_205), .B1(n_506), .B2(n_512), .Y(n_505) );
INVx4_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_135), .B(n_515), .Y(n_514) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx4f_ASAP7_75t_L g177 ( .A(n_136), .Y(n_177) );
AND2x2_ASAP7_75t_SL g161 ( .A(n_137), .B(n_162), .Y(n_161) );
AND2x4_ASAP7_75t_L g166 ( .A(n_137), .B(n_162), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_148), .B(n_160), .Y(n_138) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_146), .Y(n_140) );
INVx1_ASAP7_75t_L g510 ( .A(n_141), .Y(n_510) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
AND2x6_ASAP7_75t_L g158 ( .A(n_142), .B(n_151), .Y(n_158) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x4_ASAP7_75t_L g156 ( .A(n_144), .B(n_153), .Y(n_156) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx5_ASAP7_75t_L g159 ( .A(n_146), .Y(n_159) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_146), .Y(n_511) );
AND2x2_ASAP7_75t_L g152 ( .A(n_147), .B(n_153), .Y(n_152) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_147), .Y(n_491) );
AND2x6_ASAP7_75t_L g149 ( .A(n_150), .B(n_152), .Y(n_149) );
BUFx3_ASAP7_75t_L g492 ( .A(n_150), .Y(n_492) );
INVx2_ASAP7_75t_L g482 ( .A(n_151), .Y(n_482) );
AND2x4_ASAP7_75t_L g478 ( .A(n_152), .B(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g486 ( .A(n_153), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_157), .B(n_159), .Y(n_154) );
INVxp67_ASAP7_75t_L g579 ( .A(n_156), .Y(n_579) );
INVxp67_ASAP7_75t_L g577 ( .A(n_158), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_159), .A2(n_170), .B(n_171), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_159), .A2(n_182), .B(n_183), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_159), .A2(n_193), .B(n_194), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_159), .A2(n_202), .B(n_203), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_159), .A2(n_211), .B(n_212), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_159), .A2(n_221), .B(n_222), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_159), .A2(n_231), .B(n_232), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g483 ( .A1(n_159), .A2(n_484), .B(n_485), .C(n_487), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_SL g497 ( .A1(n_159), .A2(n_485), .B(n_498), .C(n_499), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_L g525 ( .A1(n_159), .A2(n_485), .B(n_526), .C(n_527), .Y(n_525) );
INVx1_ASAP7_75t_L g534 ( .A(n_159), .Y(n_534) );
O2A1O1Ixp33_ASAP7_75t_SL g549 ( .A1(n_159), .A2(n_485), .B(n_550), .C(n_551), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_159), .A2(n_566), .B(n_567), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_159), .B(n_166), .Y(n_580) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_160), .Y(n_224) );
OA21x2_ASAP7_75t_L g228 ( .A1(n_160), .A2(n_229), .B(n_233), .Y(n_228) );
OA21x2_ASAP7_75t_L g268 ( .A1(n_160), .A2(n_229), .B(n_233), .Y(n_268) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_175), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_164), .B(n_176), .Y(n_245) );
AND2x2_ASAP7_75t_L g306 ( .A(n_164), .B(n_275), .Y(n_306) );
AO21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_167), .B(n_173), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_165), .B(n_174), .Y(n_173) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_165), .A2(n_167), .B(n_173), .Y(n_259) );
INVx1_ASAP7_75t_SL g165 ( .A(n_166), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_166), .A2(n_179), .B(n_180), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_166), .B(n_196), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_166), .A2(n_477), .B(n_488), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_168), .B(n_172), .Y(n_167) );
AND2x2_ASAP7_75t_L g318 ( .A(n_175), .B(n_242), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_175), .B(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g362 ( .A(n_175), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g395 ( .A(n_175), .B(n_216), .Y(n_395) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g239 ( .A(n_176), .Y(n_239) );
AND2x2_ASAP7_75t_L g272 ( .A(n_176), .B(n_273), .Y(n_272) );
BUFx3_ASAP7_75t_L g307 ( .A(n_176), .Y(n_307) );
OR2x2_ASAP7_75t_L g383 ( .A(n_176), .B(n_242), .Y(n_383) );
INVx2_ASAP7_75t_SL g531 ( .A(n_177), .Y(n_531) );
OA21x2_ASAP7_75t_L g547 ( .A1(n_177), .A2(n_548), .B(n_552), .Y(n_547) );
INVx1_ASAP7_75t_SL g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_197), .Y(n_185) );
AOI211x1_ASAP7_75t_SL g312 ( .A1(n_186), .A2(n_304), .B(n_313), .C(n_315), .Y(n_312) );
AND2x2_ASAP7_75t_SL g357 ( .A(n_186), .B(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_186), .B(n_355), .Y(n_402) );
BUFx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g252 ( .A(n_187), .Y(n_252) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g227 ( .A(n_188), .Y(n_227) );
OAI21x1_ASAP7_75t_SL g188 ( .A1(n_189), .A2(n_191), .B(n_195), .Y(n_188) );
INVx1_ASAP7_75t_L g196 ( .A(n_190), .Y(n_196) );
AOI322xp5_ASAP7_75t_L g215 ( .A1(n_197), .A2(n_216), .A3(n_226), .B1(n_234), .B2(n_237), .C1(n_243), .C2(n_246), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_197), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_207), .Y(n_197) );
INVx2_ASAP7_75t_L g250 ( .A(n_198), .Y(n_250) );
INVxp67_ASAP7_75t_L g292 ( .A(n_198), .Y(n_292) );
BUFx3_ASAP7_75t_L g356 ( .A(n_198), .Y(n_356) );
AO21x2_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_205), .B(n_206), .Y(n_198) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_199), .A2(n_205), .B(n_206), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_200), .B(n_204), .Y(n_199) );
AO21x2_ASAP7_75t_L g207 ( .A1(n_205), .A2(n_208), .B(n_214), .Y(n_207) );
AO21x2_ASAP7_75t_L g254 ( .A1(n_205), .A2(n_208), .B(n_214), .Y(n_254) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_205), .A2(n_522), .B(n_528), .Y(n_521) );
AO21x2_ASAP7_75t_L g544 ( .A1(n_205), .A2(n_522), .B(n_528), .Y(n_544) );
INVx2_ASAP7_75t_L g265 ( .A(n_207), .Y(n_265) );
AND2x2_ASAP7_75t_L g314 ( .A(n_207), .B(n_228), .Y(n_314) );
AND2x2_ASAP7_75t_L g358 ( .A(n_207), .B(n_267), .Y(n_358) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_209), .B(n_213), .Y(n_208) );
AND2x2_ASAP7_75t_L g243 ( .A(n_216), .B(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_216), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_SL g437 ( .A(n_216), .B(n_272), .Y(n_437) );
INVx4_ASAP7_75t_L g242 ( .A(n_217), .Y(n_242) );
AND2x2_ASAP7_75t_L g274 ( .A(n_217), .B(n_275), .Y(n_274) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_217), .Y(n_327) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_224), .B(n_225), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_219), .B(n_223), .Y(n_218) );
AO21x2_ASAP7_75t_L g493 ( .A1(n_224), .A2(n_494), .B(n_500), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g336 ( .A(n_226), .B(n_311), .Y(n_336) );
INVx1_ASAP7_75t_SL g375 ( .A(n_226), .Y(n_375) );
AND2x4_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
AND2x4_ASAP7_75t_L g266 ( .A(n_227), .B(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_227), .B(n_265), .Y(n_334) );
AND2x2_ASAP7_75t_L g386 ( .A(n_227), .B(n_236), .Y(n_386) );
OR2x2_ASAP7_75t_L g410 ( .A(n_227), .B(n_228), .Y(n_410) );
AND2x2_ASAP7_75t_L g234 ( .A(n_228), .B(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g284 ( .A(n_228), .B(n_265), .Y(n_284) );
AND2x2_ASAP7_75t_SL g340 ( .A(n_228), .B(n_252), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_234), .B(n_347), .Y(n_364) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
BUFx2_ASAP7_75t_L g299 ( .A(n_236), .Y(n_299) );
AND2x4_ASAP7_75t_SL g339 ( .A(n_236), .B(n_253), .Y(n_339) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_240), .Y(n_237) );
OR2x2_ASAP7_75t_L g287 ( .A(n_238), .B(n_241), .Y(n_287) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g256 ( .A(n_239), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g404 ( .A(n_239), .B(n_317), .Y(n_404) );
AND2x2_ASAP7_75t_L g420 ( .A(n_239), .B(n_274), .Y(n_420) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AOI311xp33_ASAP7_75t_L g390 ( .A1(n_241), .A2(n_329), .A3(n_391), .B(n_393), .C(n_400), .Y(n_390) );
AND2x4_ASAP7_75t_L g257 ( .A(n_242), .B(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g261 ( .A(n_242), .Y(n_261) );
NAND2x1p5_ASAP7_75t_L g331 ( .A(n_242), .B(n_275), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_242), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g374 ( .A(n_242), .B(n_361), .Y(n_374) );
AND2x2_ASAP7_75t_L g260 ( .A(n_244), .B(n_261), .Y(n_260) );
INVxp67_ASAP7_75t_SL g244 ( .A(n_245), .Y(n_244) );
INVxp67_ASAP7_75t_SL g278 ( .A(n_245), .Y(n_278) );
OR2x2_ASAP7_75t_L g367 ( .A(n_245), .B(n_331), .Y(n_367) );
INVx1_ASAP7_75t_L g423 ( .A(n_245), .Y(n_423) );
INVx1_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_251), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g332 ( .A(n_249), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g346 ( .A(n_249), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g421 ( .A(n_249), .B(n_294), .Y(n_421) );
BUFx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g264 ( .A(n_250), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g283 ( .A(n_250), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g345 ( .A(n_251), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_251), .A2(n_401), .B1(n_402), .B2(n_403), .Y(n_400) );
OR2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
AND2x2_ASAP7_75t_L g294 ( .A(n_252), .B(n_265), .Y(n_294) );
AND2x4_ASAP7_75t_L g347 ( .A(n_252), .B(n_254), .Y(n_347) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OAI21xp33_ASAP7_75t_SL g255 ( .A1(n_256), .A2(n_260), .B(n_262), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g341 ( .A1(n_256), .A2(n_342), .B1(n_346), .B2(n_348), .Y(n_341) );
AND2x2_ASAP7_75t_SL g301 ( .A(n_257), .B(n_275), .Y(n_301) );
INVx2_ASAP7_75t_L g363 ( .A(n_257), .Y(n_363) );
AND2x2_ASAP7_75t_L g377 ( .A(n_257), .B(n_373), .Y(n_377) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g273 ( .A(n_259), .Y(n_273) );
INVx1_ASAP7_75t_L g326 ( .A(n_259), .Y(n_326) );
INVx1_ASAP7_75t_L g277 ( .A(n_261), .Y(n_277) );
AND3x2_ASAP7_75t_L g305 ( .A(n_261), .B(n_306), .C(n_307), .Y(n_305) );
INVx1_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
INVx1_ASAP7_75t_L g369 ( .A(n_264), .Y(n_369) );
AND2x2_ASAP7_75t_L g297 ( .A(n_266), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g368 ( .A(n_266), .B(n_369), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g379 ( .A1(n_266), .A2(n_380), .B1(n_384), .B2(n_387), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_266), .B(n_414), .Y(n_418) );
BUFx2_ASAP7_75t_L g309 ( .A(n_267), .Y(n_309) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g280 ( .A(n_268), .Y(n_280) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_268), .Y(n_399) );
OAI221xp5_ASAP7_75t_SL g269 ( .A1(n_270), .A2(n_279), .B1(n_281), .B2(n_282), .C(n_285), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_271), .B(n_276), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
INVx1_ASAP7_75t_L g361 ( .A(n_273), .Y(n_361) );
INVx2_ASAP7_75t_SL g350 ( .A(n_274), .Y(n_350) );
AND2x2_ASAP7_75t_L g432 ( .A(n_274), .B(n_299), .Y(n_432) );
INVx4_ASAP7_75t_L g323 ( .A(n_275), .Y(n_323) );
INVx1_ASAP7_75t_L g281 ( .A(n_276), .Y(n_281) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AND2x4_ASAP7_75t_L g392 ( .A(n_280), .B(n_347), .Y(n_392) );
INVx1_ASAP7_75t_SL g431 ( .A(n_280), .Y(n_431) );
AND2x2_ASAP7_75t_L g436 ( .A(n_280), .B(n_339), .Y(n_436) );
INVx1_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g378 ( .A(n_284), .Y(n_378) );
OAI21xp5_ASAP7_75t_SL g285 ( .A1(n_286), .A2(n_288), .B(n_290), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
INVx1_ASAP7_75t_L g311 ( .A(n_292), .Y(n_311) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g308 ( .A(n_294), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g398 ( .A(n_294), .B(n_399), .Y(n_398) );
OAI211xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_300), .B(n_302), .C(n_319), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g391 ( .A(n_298), .B(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_299), .B(n_314), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_299), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g424 ( .A(n_299), .B(n_347), .Y(n_424) );
OAI221xp5_ASAP7_75t_SL g335 ( .A1(n_300), .A2(n_324), .B1(n_336), .B2(n_337), .C(n_341), .Y(n_335) );
INVx3_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g406 ( .A(n_301), .B(n_307), .Y(n_406) );
OAI32xp33_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_308), .A3(n_310), .B1(n_312), .B2(n_316), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVxp67_ASAP7_75t_SL g396 ( .A(n_306), .Y(n_396) );
INVx2_ASAP7_75t_L g329 ( .A(n_307), .Y(n_329) );
O2A1O1Ixp33_ASAP7_75t_L g438 ( .A1(n_307), .A2(n_359), .B(n_439), .C(n_440), .Y(n_438) );
INVx1_ASAP7_75t_L g344 ( .A(n_309), .Y(n_344) );
OR2x2_ASAP7_75t_L g440 ( .A(n_309), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_313), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g401 ( .A(n_316), .Y(n_401) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx1_ASAP7_75t_L g382 ( .A(n_317), .Y(n_382) );
OAI21xp33_ASAP7_75t_SL g319 ( .A1(n_320), .A2(n_328), .B(n_332), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
OR2x2_ASAP7_75t_L g359 ( .A(n_322), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_323), .B(n_326), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_327), .Y(n_324) );
AOI221xp5_ASAP7_75t_L g425 ( .A1(n_325), .A2(n_357), .B1(n_426), .B2(n_429), .C(n_433), .Y(n_425) );
INVx2_ASAP7_75t_L g428 ( .A(n_325), .Y(n_428) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
OR2x2_ASAP7_75t_L g349 ( .A(n_329), .B(n_350), .Y(n_349) );
AND2x4_ASAP7_75t_L g416 ( .A(n_329), .B(n_374), .Y(n_416) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVxp67_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx1_ASAP7_75t_L g414 ( .A(n_339), .Y(n_414) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_347), .B(n_377), .Y(n_434) );
INVx2_ASAP7_75t_L g441 ( .A(n_347), .Y(n_441) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OAI221xp5_ASAP7_75t_L g411 ( .A1(n_349), .A2(n_412), .B1(n_415), .B2(n_417), .C(n_419), .Y(n_411) );
AND5x1_ASAP7_75t_L g351 ( .A(n_352), .B(n_390), .C(n_405), .D(n_425), .E(n_435), .Y(n_351) );
NOR2xp33_ASAP7_75t_SL g352 ( .A(n_353), .B(n_370), .Y(n_352) );
OAI221xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_359), .B1(n_362), .B2(n_364), .C(n_365), .Y(n_353) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_355), .B(n_357), .Y(n_354) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_368), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OAI221xp5_ASAP7_75t_SL g370 ( .A1(n_371), .A2(n_375), .B1(n_376), .B2(n_378), .C(n_379), .Y(n_370) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
AND2x4_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_375), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
OR2x2_ASAP7_75t_L g388 ( .A(n_383), .B(n_389), .Y(n_388) );
CKINVDCx16_ASAP7_75t_R g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
AOI21xp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_396), .B(n_397), .Y(n_393) );
INVx1_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_407), .B(n_411), .Y(n_405) );
INVx1_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVxp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B1(n_422), .B2(n_424), .Y(n_419) );
O2A1O1Ixp33_ASAP7_75t_L g435 ( .A1(n_421), .A2(n_436), .B(n_437), .C(n_438), .Y(n_435) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx1_ASAP7_75t_L g439 ( .A(n_432), .Y(n_439) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AOI22x1_ASAP7_75t_L g459 ( .A1(n_443), .A2(n_460), .B1(n_463), .B2(n_465), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_446), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
CKINVDCx11_ASAP7_75t_R g455 ( .A(n_456), .Y(n_455) );
CKINVDCx8_ASAP7_75t_R g456 ( .A(n_457), .Y(n_456) );
OAI21xp33_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_797), .B(n_806), .Y(n_458) );
INVx3_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
CKINVDCx5p33_ASAP7_75t_R g461 ( .A(n_462), .Y(n_461) );
CKINVDCx11_ASAP7_75t_R g810 ( .A(n_462), .Y(n_810) );
INVx1_ASAP7_75t_SL g808 ( .A(n_463), .Y(n_808) );
CKINVDCx11_ASAP7_75t_R g463 ( .A(n_464), .Y(n_463) );
OAI22x1_ASAP7_75t_L g807 ( .A1(n_465), .A2(n_808), .B1(n_809), .B2(n_810), .Y(n_807) );
INVx1_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
AND3x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_687), .C(n_750), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_651), .Y(n_468) );
NOR3xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_592), .C(n_621), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_471), .B(n_581), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_501), .B1(n_541), .B2(n_553), .Y(n_471) );
NAND2x1_ASAP7_75t_L g736 ( .A(n_472), .B(n_582), .Y(n_736) );
INVx2_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_493), .Y(n_473) );
INVx2_ASAP7_75t_L g555 ( .A(n_474), .Y(n_555) );
INVx4_ASAP7_75t_L g597 ( .A(n_474), .Y(n_597) );
BUFx6f_ASAP7_75t_L g617 ( .A(n_474), .Y(n_617) );
AND2x4_ASAP7_75t_L g628 ( .A(n_474), .B(n_596), .Y(n_628) );
AND2x2_ASAP7_75t_L g634 ( .A(n_474), .B(n_558), .Y(n_634) );
NOR2x1_ASAP7_75t_SL g764 ( .A(n_474), .B(n_569), .Y(n_764) );
OR2x6_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
INVxp67_ASAP7_75t_L g517 ( .A(n_478), .Y(n_517) );
NOR2x1p5_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
INVx1_ASAP7_75t_L g538 ( .A(n_481), .Y(n_538) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OR2x6_ASAP7_75t_L g485 ( .A(n_482), .B(n_486), .Y(n_485) );
INVxp67_ASAP7_75t_L g507 ( .A(n_485), .Y(n_507) );
INVx2_ASAP7_75t_L g568 ( .A(n_485), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_485), .A2(n_510), .B1(n_573), .B2(n_574), .Y(n_572) );
AND2x2_ASAP7_75t_L g490 ( .A(n_486), .B(n_491), .Y(n_490) );
INVxp33_ASAP7_75t_L g537 ( .A(n_486), .Y(n_537) );
INVx1_ASAP7_75t_L g519 ( .A(n_489), .Y(n_519) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_492), .Y(n_489) );
INVx1_ASAP7_75t_L g561 ( .A(n_490), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_492), .Y(n_562) );
INVx2_ASAP7_75t_L g600 ( .A(n_493), .Y(n_600) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_493), .Y(n_614) );
INVx1_ASAP7_75t_L g625 ( .A(n_493), .Y(n_625) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_493), .Y(n_637) );
AND2x2_ASAP7_75t_L g669 ( .A(n_493), .B(n_569), .Y(n_669) );
AND2x2_ASAP7_75t_L g701 ( .A(n_493), .B(n_585), .Y(n_701) );
INVx1_ASAP7_75t_L g708 ( .A(n_493), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_520), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g650 ( .A(n_503), .B(n_589), .Y(n_650) );
INVx2_ASAP7_75t_L g724 ( .A(n_503), .Y(n_724) );
AND2x2_ASAP7_75t_L g747 ( .A(n_503), .B(n_520), .Y(n_747) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_504), .B(n_544), .Y(n_588) );
INVx2_ASAP7_75t_L g609 ( .A(n_504), .Y(n_609) );
AND2x4_ASAP7_75t_L g631 ( .A(n_504), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g666 ( .A(n_504), .Y(n_666) );
AND2x2_ASAP7_75t_L g743 ( .A(n_504), .B(n_547), .Y(n_743) );
OR2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_513), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_509), .B(n_510), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_517), .B1(n_518), .B2(n_519), .Y(n_513) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g714 ( .A(n_520), .Y(n_714) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_529), .Y(n_520) );
NOR2xp67_ASAP7_75t_L g639 ( .A(n_521), .B(n_609), .Y(n_639) );
AND2x2_ASAP7_75t_L g644 ( .A(n_521), .B(n_609), .Y(n_644) );
INVx2_ASAP7_75t_L g657 ( .A(n_521), .Y(n_657) );
NOR2x1_ASAP7_75t_L g705 ( .A(n_521), .B(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
AND2x4_ASAP7_75t_L g630 ( .A(n_529), .B(n_543), .Y(n_630) );
AND2x2_ASAP7_75t_L g645 ( .A(n_529), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g698 ( .A(n_529), .Y(n_698) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_530), .B(n_547), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_530), .B(n_544), .Y(n_702) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_532), .B(n_540), .Y(n_530) );
AO21x2_ASAP7_75t_L g591 ( .A1(n_531), .A2(n_532), .B(n_540), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_533), .B(n_539), .Y(n_532) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVxp33_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2x1p5_ASAP7_75t_L g542 ( .A(n_543), .B(n_545), .Y(n_542) );
INVx3_ASAP7_75t_L g606 ( .A(n_543), .Y(n_606) );
INVx3_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_544), .Y(n_604) );
AND2x2_ASAP7_75t_L g773 ( .A(n_544), .B(n_774), .Y(n_773) );
INVx3_ASAP7_75t_L g661 ( .A(n_545), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_545), .B(n_698), .Y(n_793) );
BUFx3_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g608 ( .A(n_546), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x4_ASAP7_75t_L g589 ( .A(n_547), .B(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g632 ( .A(n_547), .Y(n_632) );
INVxp67_ASAP7_75t_L g646 ( .A(n_547), .Y(n_646) );
INVx1_ASAP7_75t_L g706 ( .A(n_547), .Y(n_706) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_547), .Y(n_774) );
INVx1_ASAP7_75t_L g758 ( .A(n_553), .Y(n_758) );
NOR2x1_ASAP7_75t_L g553 ( .A(n_554), .B(n_556), .Y(n_553) );
NOR2x1_ASAP7_75t_L g678 ( .A(n_554), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g712 ( .A(n_555), .B(n_584), .Y(n_712) );
OR2x2_ASAP7_75t_L g748 ( .A(n_556), .B(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g730 ( .A(n_557), .B(n_708), .Y(n_730) );
AND2x2_ASAP7_75t_L g782 ( .A(n_557), .B(n_617), .Y(n_782) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_569), .Y(n_557) );
AND2x4_ASAP7_75t_L g584 ( .A(n_558), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g596 ( .A(n_558), .Y(n_596) );
INVx2_ASAP7_75t_L g613 ( .A(n_558), .Y(n_613) );
HB1xp67_ASAP7_75t_L g791 ( .A(n_558), .Y(n_791) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_564), .Y(n_558) );
NOR3xp33_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .C(n_563), .Y(n_560) );
INVx3_ASAP7_75t_L g585 ( .A(n_569), .Y(n_585) );
INVx2_ASAP7_75t_L g679 ( .A(n_569), .Y(n_679) );
AND2x4_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
OAI21xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_575), .B(n_580), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_577), .B1(n_578), .B2(n_579), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_586), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_583), .B(n_659), .Y(n_676) );
NOR2x1_ASAP7_75t_L g718 ( .A(n_583), .B(n_597), .Y(n_718) );
INVx4_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_584), .B(n_659), .Y(n_796) );
AND2x2_ASAP7_75t_L g612 ( .A(n_585), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g626 ( .A(n_585), .Y(n_626) );
AOI22xp5_ASAP7_75t_SL g674 ( .A1(n_586), .A2(n_675), .B1(n_676), .B2(n_677), .Y(n_674) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
NAND2x1p5_ASAP7_75t_L g671 ( .A(n_587), .B(n_645), .Y(n_671) );
INVx2_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g732 ( .A(n_588), .B(n_620), .Y(n_732) );
AND2x2_ASAP7_75t_L g602 ( .A(n_589), .B(n_603), .Y(n_602) );
AND2x4_ASAP7_75t_L g638 ( .A(n_589), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g734 ( .A(n_589), .B(n_724), .Y(n_734) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x4_ASAP7_75t_L g656 ( .A(n_591), .B(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g682 ( .A(n_591), .Y(n_682) );
AND2x2_ASAP7_75t_L g772 ( .A(n_591), .B(n_609), .Y(n_772) );
OAI221xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_601), .B1(n_605), .B2(n_610), .C(n_615), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_598), .Y(n_594) );
INVx1_ASAP7_75t_L g673 ( .A(n_595), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_595), .B(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_595), .B(n_669), .Y(n_788) );
AND2x4_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
NOR2xp67_ASAP7_75t_SL g641 ( .A(n_597), .B(n_642), .Y(n_641) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_597), .Y(n_654) );
OR2x2_ASAP7_75t_L g738 ( .A(n_597), .B(n_739), .Y(n_738) );
AND2x4_ASAP7_75t_SL g790 ( .A(n_597), .B(n_791), .Y(n_790) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx3_ASAP7_75t_L g659 ( .A(n_599), .Y(n_659) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
HB1xp67_ASAP7_75t_L g749 ( .A(n_600), .Y(n_749) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AOI221x1_ASAP7_75t_L g689 ( .A1(n_602), .A2(n_690), .B1(n_692), .B2(n_695), .C(n_699), .Y(n_689) );
AND2x2_ASAP7_75t_L g675 ( .A(n_603), .B(n_631), .Y(n_675) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
AND2x2_ASAP7_75t_L g618 ( .A(n_606), .B(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_606), .B(n_608), .Y(n_745) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
AND2x2_ASAP7_75t_SL g616 ( .A(n_612), .B(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_612), .B(n_625), .Y(n_642) );
INVx2_ASAP7_75t_L g649 ( .A(n_612), .Y(n_649) );
INVx1_ASAP7_75t_L g694 ( .A(n_613), .Y(n_694) );
BUFx2_ASAP7_75t_L g783 ( .A(n_614), .Y(n_783) );
NAND2xp33_ASAP7_75t_SL g615 ( .A(n_616), .B(n_618), .Y(n_615) );
OR2x6_ASAP7_75t_L g648 ( .A(n_617), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g729 ( .A(n_617), .B(n_669), .Y(n_729) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_640), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_629), .B1(n_633), .B2(n_638), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_624), .B(n_627), .Y(n_623) );
AND2x2_ASAP7_75t_SL g686 ( .A(n_624), .B(n_628), .Y(n_686) );
AND2x4_ASAP7_75t_L g692 ( .A(n_624), .B(n_693), .Y(n_692) );
AND2x4_ASAP7_75t_SL g624 ( .A(n_625), .B(n_626), .Y(n_624) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_625), .Y(n_717) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_628), .B(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_628), .B(n_659), .Y(n_691) );
HB1xp67_ASAP7_75t_L g775 ( .A(n_628), .Y(n_775) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
AND2x2_ASAP7_75t_L g722 ( .A(n_630), .B(n_723), .Y(n_722) );
INVx3_ASAP7_75t_L g683 ( .A(n_631), .Y(n_683) );
NAND2x1_ASAP7_75t_SL g727 ( .A(n_631), .B(n_682), .Y(n_727) );
AND2x2_ASAP7_75t_L g761 ( .A(n_631), .B(n_656), .Y(n_761) );
AND2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_643), .B1(n_647), .B2(n_650), .Y(n_640) );
BUFx2_ASAP7_75t_L g756 ( .A(n_642), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_643), .A2(n_712), .B1(n_786), .B2(n_795), .Y(n_794) );
AND2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
NAND2x1p5_ASAP7_75t_L g697 ( .A(n_644), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g664 ( .A(n_645), .B(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND3xp33_ASAP7_75t_L g780 ( .A(n_649), .B(n_781), .C(n_783), .Y(n_780) );
INVx1_ASAP7_75t_L g684 ( .A(n_650), .Y(n_684) );
AOI211x1_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_660), .B(n_662), .C(n_680), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g711 ( .A(n_655), .B(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_658), .Y(n_655) );
AND2x2_ASAP7_75t_L g742 ( .A(n_656), .B(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_656), .B(n_723), .Y(n_754) );
AND2x2_ASAP7_75t_L g786 ( .A(n_656), .B(n_724), .Y(n_786) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g767 ( .A(n_659), .Y(n_767) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OR2x2_ASAP7_75t_L g696 ( .A(n_661), .B(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_674), .Y(n_662) );
AOI22xp5_ASAP7_75t_SL g663 ( .A1(n_664), .A2(n_667), .B1(n_670), .B2(n_672), .Y(n_663) );
BUFx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g704 ( .A(n_666), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_SL g719 ( .A(n_666), .Y(n_719) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_SL g789 ( .A(n_669), .B(n_790), .Y(n_789) );
INVx3_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVxp67_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g725 ( .A(n_678), .B(n_708), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_684), .B(n_685), .Y(n_680) );
OR2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_682), .B(n_704), .Y(n_779) );
OR2x2_ASAP7_75t_L g757 ( .A(n_683), .B(n_702), .Y(n_757) );
INVx1_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NAND3x1_ASAP7_75t_L g688 ( .A(n_689), .B(n_709), .C(n_733), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_692), .A2(n_722), .B1(n_725), .B2(n_726), .Y(n_721) );
NAND2xp5_ASAP7_75t_SL g707 ( .A(n_693), .B(n_708), .Y(n_707) );
INVx2_ASAP7_75t_SL g766 ( .A(n_693), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_693), .B(n_767), .Y(n_770) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
OAI222xp33_ASAP7_75t_L g753 ( .A1(n_697), .A2(n_754), .B1(n_755), .B2(n_756), .C1(n_757), .C2(n_758), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_702), .B1(n_703), .B2(n_707), .Y(n_699) );
INVx1_ASAP7_75t_SL g739 ( .A(n_701), .Y(n_739) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g776 ( .A(n_705), .B(n_772), .Y(n_776) );
NOR2x1_ASAP7_75t_L g709 ( .A(n_710), .B(n_720), .Y(n_709) );
AOI21xp5_ASAP7_75t_SL g710 ( .A1(n_711), .A2(n_713), .B(n_719), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_728), .Y(n_720) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_727), .B(n_741), .Y(n_740) );
OAI21xp5_ASAP7_75t_SL g728 ( .A1(n_729), .A2(n_730), .B(n_731), .Y(n_728) );
INVx1_ASAP7_75t_L g755 ( .A(n_730), .Y(n_755) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
AOI221xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_735), .B1(n_737), .B2(n_740), .C(n_744), .Y(n_733) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVxp67_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
AOI21xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B(n_748), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVxp67_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
NAND3x1_ASAP7_75t_L g751 ( .A(n_752), .B(n_777), .C(n_784), .Y(n_751) );
NOR2x1_ASAP7_75t_L g752 ( .A(n_753), .B(n_759), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_760), .B(n_768), .Y(n_759) );
NAND2xp5_ASAP7_75t_SL g760 ( .A(n_761), .B(n_762), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_763), .B(n_765), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_763), .B(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
AOI22xp5_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_771), .B1(n_775), .B2(n_776), .Y(n_768) );
AND2x4_ASAP7_75t_L g771 ( .A(n_772), .B(n_773), .Y(n_771) );
NAND2xp5_ASAP7_75t_SL g777 ( .A(n_778), .B(n_780), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
AND2x2_ASAP7_75t_L g784 ( .A(n_785), .B(n_794), .Y(n_784) );
AOI22xp5_ASAP7_75t_SL g785 ( .A1(n_786), .A2(n_787), .B1(n_789), .B2(n_792), .Y(n_785) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVxp67_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
AOI21xp33_ASAP7_75t_L g806 ( .A1(n_797), .A2(n_807), .B(n_811), .Y(n_806) );
INVx1_ASAP7_75t_L g805 ( .A(n_798), .Y(n_805) );
INVx1_ASAP7_75t_L g803 ( .A(n_800), .Y(n_803) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .Y(n_811) );
INVx1_ASAP7_75t_SL g814 ( .A(n_815), .Y(n_814) );
INVx2_ASAP7_75t_SL g815 ( .A(n_816), .Y(n_815) );
INVx2_ASAP7_75t_SL g825 ( .A(n_816), .Y(n_825) );
AND2x2_ASAP7_75t_SL g816 ( .A(n_817), .B(n_818), .Y(n_816) );
NOR2xp33_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .Y(n_822) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
endmodule