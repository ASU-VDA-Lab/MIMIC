module real_jpeg_29460_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_206;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_0),
.A2(n_62),
.B1(n_63),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_0),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_0),
.A2(n_31),
.B1(n_32),
.B2(n_70),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_0),
.A2(n_25),
.B1(n_28),
.B2(n_70),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_1),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_1),
.B(n_80),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_1),
.B(n_62),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g138 ( 
.A1(n_1),
.A2(n_62),
.B(n_134),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_75),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_1),
.A2(n_25),
.B(n_29),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_1),
.B(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_1),
.A2(n_41),
.B1(n_103),
.B2(n_185),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_2),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_3),
.A2(n_25),
.B1(n_28),
.B2(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_4),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_6),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.Y(n_61)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_65),
.Y(n_66)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_6),
.Y(n_133)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_7),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_8),
.A2(n_73),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_8),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_8),
.A2(n_62),
.B1(n_63),
.B2(n_82),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_82),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_8),
.A2(n_25),
.B1(n_28),
.B2(n_82),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_9),
.A2(n_62),
.B1(n_63),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_9),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_9),
.A2(n_68),
.B1(n_73),
.B2(n_83),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_68),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_9),
.A2(n_25),
.B1(n_28),
.B2(n_68),
.Y(n_177)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_11),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_11),
.A2(n_55),
.B1(n_62),
.B2(n_63),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_11),
.A2(n_25),
.B1(n_28),
.B2(n_55),
.Y(n_129)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_13),
.A2(n_25),
.B1(n_28),
.B2(n_39),
.Y(n_49)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_14),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_15),
.A2(n_25),
.B1(n_28),
.B2(n_33),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_122),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_120),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_104),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_20),
.B(n_104),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_84),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_50),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_34),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_24),
.A2(n_36),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_24),
.A2(n_36),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_24),
.A2(n_36),
.B1(n_141),
.B2(n_160),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_24),
.B(n_75),
.Y(n_183)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_25),
.Y(n_28)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_27),
.A2(n_32),
.B(n_75),
.C(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_28),
.B(n_189),
.Y(n_188)
);

AOI32xp33_ASAP7_75t_L g130 ( 
.A1(n_31),
.A2(n_63),
.A3(n_131),
.B1(n_134),
.B2(n_135),
.Y(n_130)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp33_ASAP7_75t_SL g135 ( 
.A(n_32),
.B(n_132),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_53),
.B(n_56),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_36),
.A2(n_142),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_57),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_44),
.B(n_46),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_41),
.A2(n_44),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_41),
.A2(n_171),
.B(n_172),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_41),
.A2(n_116),
.B1(n_177),
.B2(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_42),
.B(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_42),
.A2(n_47),
.B(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_42),
.A2(n_117),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_49),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_58),
.C(n_71),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_51),
.A2(n_52),
.B1(n_58),
.B2(n_59),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_54),
.B(n_57),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_66),
.B1(n_67),
.B2(n_69),
.Y(n_59)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_60),
.A2(n_66),
.B1(n_67),
.B2(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_60),
.A2(n_66),
.B1(n_112),
.B2(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_66),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_63),
.B1(n_77),
.B2(n_78),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_77),
.Y(n_100)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_63),
.A2(n_72),
.B1(n_79),
.B2(n_100),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_66),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_71),
.B(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_76),
.B1(n_80),
.B2(n_81),
.Y(n_71)
);

HAxp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_75),
.CON(n_72),
.SN(n_72)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_73),
.A2(n_77),
.B(n_79),
.C(n_80),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_77),
.Y(n_79)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_75),
.B(n_116),
.Y(n_189)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_98),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_92),
.B2(n_93),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B(n_96),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_101),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_116),
.B(n_118),
.Y(n_115)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_108),
.C(n_110),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_105),
.A2(n_106),
.B1(n_203),
.B2(n_205),
.Y(n_202)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_110),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_113),
.C(n_115),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_115),
.Y(n_147)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_117),
.B(n_129),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_200),
.B(n_206),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_153),
.B(n_199),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_143),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_125),
.B(n_143),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_136),
.C(n_139),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_126),
.A2(n_127),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_130),
.Y(n_150)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_136),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_148),
.B2(n_149),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_144),
.B(n_150),
.C(n_151),
.Y(n_201)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_193),
.B(n_198),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_173),
.B(n_192),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_163),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_156),
.B(n_163),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_161),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_157),
.A2(n_158),
.B1(n_161),
.B2(n_180),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_161),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_170),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_169),
.C(n_170),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_171),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_181),
.B(n_191),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_179),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_175),
.B(n_179),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_186),
.B(n_190),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_183),
.B(n_184),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_194),
.B(n_195),
.Y(n_198)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_201),
.B(n_202),
.Y(n_206)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_203),
.Y(n_205)
);


endmodule