module fake_jpeg_25767_n_79 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_79);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_79;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_29),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_38),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_37),
.B(n_30),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_46),
.Y(n_54)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_32),
.B(n_26),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_1),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_1),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_23),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_48),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

NAND3xp33_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_2),
.C(n_3),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_51),
.A2(n_60),
.B(n_64),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_50),
.B(n_4),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_56),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_61),
.B(n_18),
.Y(n_68)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_58),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_10),
.Y(n_58)
);

NAND3xp33_ASAP7_75t_SL g60 ( 
.A(n_48),
.B(n_11),
.C(n_12),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_15),
.B(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_21),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_54),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_70),
.A2(n_59),
.B1(n_63),
.B2(n_62),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_73),
.C(n_67),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_74),
.B(n_51),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_57),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_66),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_65),
.Y(n_79)
);


endmodule