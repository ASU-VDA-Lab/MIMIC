module fake_jpeg_13242_n_432 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_432);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_432;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_4),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_27),
.B(n_16),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_56),
.B(n_62),
.Y(n_110)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_57),
.Y(n_133)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_59),
.Y(n_154)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_60),
.Y(n_123)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_27),
.B(n_16),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_64),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_65),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_36),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_66),
.B(n_84),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_68),
.Y(n_150)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_69),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_71),
.Y(n_174)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_73),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_75),
.Y(n_163)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_76),
.Y(n_162)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_35),
.B(n_10),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_78),
.B(n_87),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_80),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

INVx2_ASAP7_75t_R g84 ( 
.A(n_35),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_17),
.Y(n_86)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_37),
.B(n_8),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_29),
.B(n_11),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_92),
.Y(n_120)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_90),
.Y(n_148)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

BUFx12f_ASAP7_75t_SL g92 ( 
.A(n_29),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx4_ASAP7_75t_SL g147 ( 
.A(n_93),
.Y(n_147)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_36),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_37),
.B(n_11),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_96),
.B(n_97),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_48),
.B(n_29),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_15),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_24),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_100),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_36),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_106),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_21),
.B(n_12),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_108),
.Y(n_128)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_42),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_87),
.A2(n_50),
.B1(n_51),
.B2(n_30),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_109),
.A2(n_116),
.B1(n_0),
.B2(n_6),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_88),
.C(n_78),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_111),
.B(n_38),
.C(n_26),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_71),
.A2(n_47),
.B1(n_50),
.B2(n_42),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_113),
.A2(n_127),
.B(n_140),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_102),
.A2(n_30),
.B1(n_51),
.B2(n_43),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_119),
.B(n_153),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_76),
.A2(n_47),
.B1(n_42),
.B2(n_29),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_43),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_129),
.B(n_137),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_24),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_77),
.A2(n_54),
.B1(n_52),
.B2(n_40),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_69),
.B(n_22),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_145),
.B(n_146),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_69),
.B(n_22),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_82),
.B(n_21),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_58),
.A2(n_31),
.B1(n_54),
.B2(n_52),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_156),
.A2(n_160),
.B1(n_167),
.B2(n_172),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_99),
.A2(n_28),
.B1(n_46),
.B2(n_38),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_157),
.A2(n_0),
.B1(n_6),
.B2(n_167),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_103),
.B(n_28),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_158),
.B(n_165),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_94),
.A2(n_83),
.B1(n_73),
.B2(n_106),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_74),
.B(n_26),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_63),
.A2(n_40),
.B1(n_33),
.B2(n_31),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_79),
.B(n_55),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_171),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_81),
.B(n_55),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_70),
.A2(n_18),
.B1(n_33),
.B2(n_46),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_160),
.A2(n_85),
.B1(n_100),
.B2(n_101),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_175),
.A2(n_196),
.B1(n_202),
.B2(n_210),
.Y(n_234)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_176),
.Y(n_241)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_123),
.Y(n_177)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_177),
.Y(n_233)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_178),
.Y(n_242)
);

BUFx5_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_180),
.Y(n_260)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_126),
.Y(n_181)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

OR2x2_ASAP7_75t_SL g182 ( 
.A(n_120),
.B(n_15),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_182),
.B(n_186),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_184),
.B(n_219),
.Y(n_280)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_185),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_18),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_118),
.B(n_13),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_187),
.B(n_194),
.Y(n_261)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_125),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_188),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_159),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_189),
.B(n_216),
.Y(n_236)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_163),
.Y(n_190)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_190),
.Y(n_251)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_130),
.Y(n_191)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_191),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_117),
.B(n_36),
.C(n_3),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_192),
.B(n_35),
.C(n_88),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_130),
.Y(n_193)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_193),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_128),
.B(n_0),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_119),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_195),
.B(n_199),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_L g196 ( 
.A1(n_172),
.A2(n_0),
.B1(n_3),
.B2(n_5),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_197),
.Y(n_270)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_122),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_200),
.B(n_204),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

INVx13_ASAP7_75t_L g238 ( 
.A(n_201),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_163),
.Y(n_203)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_203),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_140),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_135),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_205),
.B(n_211),
.Y(n_269)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_147),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_206),
.Y(n_248)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_132),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_207),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_208),
.A2(n_226),
.B1(n_229),
.B2(n_169),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_110),
.A2(n_113),
.B1(n_127),
.B2(n_156),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_136),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_155),
.B(n_133),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_212),
.B(n_213),
.Y(n_278)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_122),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_132),
.Y(n_214)
);

INVx13_ASAP7_75t_L g266 ( 
.A(n_214),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_154),
.B(n_134),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_134),
.B(n_150),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_217),
.B(n_224),
.Y(n_255)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_162),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_218),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_143),
.Y(n_219)
);

O2A1O1Ixp33_ASAP7_75t_SL g220 ( 
.A1(n_148),
.A2(n_141),
.B(n_144),
.C(n_161),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_220),
.A2(n_156),
.B(n_172),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_149),
.A2(n_142),
.B1(n_124),
.B2(n_143),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_222),
.A2(n_201),
.B1(n_191),
.B2(n_193),
.Y(n_244)
);

AO22x2_ASAP7_75t_L g223 ( 
.A1(n_124),
.A2(n_142),
.B1(n_149),
.B2(n_115),
.Y(n_223)
);

AO21x2_ASAP7_75t_L g262 ( 
.A1(n_223),
.A2(n_203),
.B(n_206),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_138),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_150),
.B(n_112),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_225),
.B(n_227),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_162),
.A2(n_138),
.B1(n_114),
.B2(n_121),
.Y(n_226)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_147),
.Y(n_227)
);

OR2x2_ASAP7_75t_SL g228 ( 
.A(n_131),
.B(n_112),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_232),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_115),
.A2(n_166),
.B1(n_114),
.B2(n_174),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_121),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_230),
.Y(n_259)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_131),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_237),
.B(n_244),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_L g240 ( 
.A1(n_221),
.A2(n_169),
.B1(n_204),
.B2(n_175),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_240),
.A2(n_243),
.B1(n_250),
.B2(n_253),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_221),
.A2(n_198),
.B1(n_183),
.B2(n_209),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_186),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_247),
.B(n_254),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_229),
.A2(n_196),
.B1(n_223),
.B2(n_231),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_223),
.A2(n_220),
.B1(n_218),
.B2(n_179),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_176),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_223),
.A2(n_224),
.B1(n_207),
.B2(n_214),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_256),
.A2(n_272),
.B1(n_273),
.B2(n_240),
.Y(n_293)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_262),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_212),
.B(n_182),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_265),
.B(n_267),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_230),
.B(n_232),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_219),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_268),
.B(n_274),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_265),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_208),
.A2(n_195),
.B1(n_221),
.B2(n_204),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_204),
.A2(n_221),
.B1(n_157),
.B2(n_208),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_183),
.B(n_194),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_276),
.A2(n_234),
.B(n_264),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_247),
.C(n_246),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_281),
.B(n_270),
.C(n_277),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_282),
.B(n_285),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_245),
.B(n_274),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_283),
.B(n_308),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_245),
.B(n_252),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_286),
.A2(n_277),
.B(n_257),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_236),
.B(n_261),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_288),
.B(n_295),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_246),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_290),
.Y(n_319)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_241),
.Y(n_292)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_292),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_293),
.A2(n_302),
.B(n_315),
.Y(n_340)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_267),
.Y(n_294)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_294),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_249),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_253),
.A2(n_250),
.B1(n_234),
.B2(n_256),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_296),
.A2(n_309),
.B1(n_289),
.B2(n_293),
.Y(n_338)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_297),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_269),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_298),
.B(n_301),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_276),
.A2(n_254),
.B(n_245),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_299),
.A2(n_311),
.B(n_313),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_249),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_300),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_278),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_255),
.B(n_239),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_242),
.Y(n_303)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_303),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_263),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_305),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_279),
.B(n_242),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_306),
.B(n_310),
.Y(n_324)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_251),
.Y(n_307)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_307),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_271),
.B(n_262),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_262),
.A2(n_239),
.B1(n_259),
.B2(n_244),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_251),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_262),
.B(n_241),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_248),
.B(n_258),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_312),
.B(n_298),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_262),
.A2(n_233),
.B(n_235),
.Y(n_313)
);

AOI21xp33_ASAP7_75t_L g315 ( 
.A1(n_266),
.A2(n_263),
.B(n_260),
.Y(n_315)
);

AOI322xp5_ASAP7_75t_L g317 ( 
.A1(n_286),
.A2(n_266),
.A3(n_238),
.B1(n_257),
.B2(n_235),
.C1(n_233),
.C2(n_270),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_317),
.B(n_332),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_318),
.A2(n_337),
.B(n_311),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_321),
.B(n_328),
.C(n_336),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_312),
.Y(n_325)
);

BUFx12f_ASAP7_75t_L g348 ( 
.A(n_325),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_281),
.B(n_238),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_329),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_302),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_331),
.B(n_308),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_314),
.B(n_294),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_287),
.B(n_304),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_299),
.A2(n_313),
.B(n_311),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_338),
.A2(n_291),
.B1(n_296),
.B2(n_284),
.Y(n_361)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_335),
.Y(n_343)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_343),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_337),
.A2(n_290),
.B(n_302),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_344),
.A2(n_349),
.B(n_353),
.Y(n_375)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_335),
.Y(n_345)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_345),
.Y(n_378)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_339),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_347),
.B(n_351),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_322),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_297),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_352),
.B(n_355),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_326),
.B(n_287),
.C(n_283),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_354),
.B(n_360),
.C(n_321),
.Y(n_369)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_339),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_324),
.B(n_314),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_356),
.B(n_358),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_323),
.A2(n_289),
.B(n_295),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_357),
.A2(n_340),
.B(n_323),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_322),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_336),
.B(n_304),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_359),
.B(n_362),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_326),
.B(n_284),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_361),
.A2(n_327),
.B1(n_318),
.B2(n_309),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_341),
.B(n_288),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_342),
.A2(n_338),
.B1(n_319),
.B2(n_340),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_363),
.A2(n_365),
.B1(n_348),
.B2(n_351),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_364),
.A2(n_316),
.B(n_350),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_357),
.A2(n_330),
.B1(n_327),
.B2(n_291),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_354),
.B(n_349),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_369),
.B(n_373),
.C(n_379),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_346),
.B(n_329),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_370),
.B(n_360),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_346),
.B(n_331),
.C(n_330),
.Y(n_373)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_376),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_361),
.A2(n_341),
.B1(n_334),
.B2(n_333),
.Y(n_377)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_377),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_346),
.B(n_319),
.C(n_325),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_371),
.B(n_362),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_380),
.B(n_389),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_372),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_381),
.B(n_382),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_370),
.B(n_379),
.Y(n_382)
);

NAND4xp25_ASAP7_75t_SL g383 ( 
.A(n_372),
.B(n_301),
.C(n_356),
.D(n_358),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_383),
.B(n_393),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_369),
.B(n_360),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_386),
.B(n_388),
.C(n_391),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_366),
.B(n_316),
.Y(n_389)
);

A2O1A1Ixp33_ASAP7_75t_L g390 ( 
.A1(n_374),
.A2(n_353),
.B(n_352),
.C(n_344),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_390),
.B(n_364),
.Y(n_403)
);

XNOR2x1_ASAP7_75t_L g394 ( 
.A(n_392),
.B(n_365),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_373),
.B(n_359),
.C(n_324),
.Y(n_393)
);

XNOR2x1_ASAP7_75t_L g408 ( 
.A(n_394),
.B(n_399),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_387),
.A2(n_350),
.B1(n_363),
.B2(n_374),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_396),
.B(n_398),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_385),
.Y(n_398)
);

XNOR2x1_ASAP7_75t_L g399 ( 
.A(n_392),
.B(n_367),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_391),
.B(n_285),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_400),
.B(n_348),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_403),
.A2(n_375),
.B(n_393),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_385),
.B(n_348),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_404),
.B(n_405),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_383),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_403),
.A2(n_387),
.B1(n_375),
.B2(n_390),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_406),
.A2(n_388),
.B1(n_378),
.B2(n_368),
.Y(n_417)
);

AO21x1_ASAP7_75t_L g416 ( 
.A1(n_407),
.A2(n_404),
.B(n_394),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_397),
.B(n_395),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_409),
.B(n_410),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_401),
.B(n_348),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_413),
.B(n_348),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_402),
.B(n_399),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_414),
.B(n_402),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_415),
.B(n_417),
.C(n_414),
.Y(n_423)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_416),
.Y(n_422)
);

AOI21x1_ASAP7_75t_L g421 ( 
.A1(n_419),
.A2(n_420),
.B(n_407),
.Y(n_421)
);

NOR2xp67_ASAP7_75t_L g420 ( 
.A(n_406),
.B(n_384),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_421),
.B(n_423),
.Y(n_427)
);

AOI21x1_ASAP7_75t_L g424 ( 
.A1(n_418),
.A2(n_412),
.B(n_411),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_424),
.Y(n_425)
);

AOI322xp5_ASAP7_75t_L g426 ( 
.A1(n_422),
.A2(n_411),
.A3(n_416),
.B1(n_345),
.B2(n_343),
.C1(n_355),
.C2(n_347),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_426),
.A2(n_320),
.B(n_305),
.Y(n_429)
);

OA21x2_ASAP7_75t_SL g428 ( 
.A1(n_425),
.A2(n_415),
.B(n_384),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_428),
.B(n_429),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_430),
.B(n_427),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_431),
.B(n_408),
.Y(n_432)
);


endmodule