module fake_jpeg_25507_n_311 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_311);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_27),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_18),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_45),
.B(n_58),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_51),
.Y(n_79)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_49),
.Y(n_67)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_54),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_19),
.Y(n_54)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_19),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_59),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_18),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_42),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_27),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_60),
.B(n_41),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_42),
.B1(n_32),
.B2(n_40),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_63),
.A2(n_70),
.B1(n_73),
.B2(n_81),
.Y(n_103)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_0),
.B(n_1),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_66),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_43),
.A2(n_28),
.B1(n_30),
.B2(n_40),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_69),
.A2(n_49),
.B1(n_61),
.B2(n_53),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_43),
.A2(n_32),
.B1(n_28),
.B2(n_30),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_72),
.Y(n_100)
);

INVxp33_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_45),
.A2(n_28),
.B1(n_30),
.B2(n_27),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_65),
.Y(n_94)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_87),
.Y(n_109)
);

AOI22x1_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_58),
.B1(n_45),
.B2(n_48),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_89),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_48),
.A2(n_29),
.B1(n_25),
.B2(n_22),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_84),
.A2(n_90),
.B1(n_25),
.B2(n_29),
.Y(n_108)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_41),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_82),
.C(n_70),
.Y(n_97)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_88),
.B(n_52),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_19),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_51),
.A2(n_22),
.B1(n_31),
.B2(n_25),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_92),
.B(n_111),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_93),
.A2(n_73),
.B1(n_67),
.B2(n_85),
.Y(n_134)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_102),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_99),
.C(n_86),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_90),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_98),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_22),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_110),
.Y(n_144)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_107),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_108),
.A2(n_84),
.B1(n_81),
.B2(n_77),
.Y(n_123)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_59),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_62),
.Y(n_112)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

INVxp67_ASAP7_75t_SL g142 ( 
.A(n_114),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_77),
.A2(n_31),
.B1(n_16),
.B2(n_20),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_116),
.A2(n_20),
.B1(n_16),
.B2(n_24),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_71),
.B(n_44),
.Y(n_117)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_89),
.B(n_44),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_79),
.B(n_86),
.C(n_66),
.Y(n_130)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_119),
.Y(n_137)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_124),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_123),
.B(n_103),
.Y(n_156)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_112),
.A2(n_78),
.B(n_88),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_125),
.A2(n_140),
.B(n_130),
.Y(n_170)
);

MAJx2_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_81),
.C(n_79),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_100),
.C(n_92),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_139),
.Y(n_145)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_134),
.A2(n_136),
.B1(n_141),
.B2(n_68),
.Y(n_152)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_96),
.A2(n_86),
.B1(n_87),
.B2(n_76),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_105),
.A2(n_29),
.B(n_31),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_98),
.A2(n_64),
.B1(n_49),
.B2(n_62),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_144),
.B1(n_140),
.B2(n_133),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_129),
.A2(n_103),
.B1(n_111),
.B2(n_113),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_146),
.A2(n_157),
.B1(n_158),
.B2(n_163),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_91),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_154),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_91),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_148),
.B(n_160),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_126),
.B(n_110),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_149),
.B(n_159),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_157),
.Y(n_180)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_99),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_162),
.Y(n_179)
);

OAI32xp33_ASAP7_75t_L g187 ( 
.A1(n_156),
.A2(n_158),
.A3(n_147),
.B1(n_155),
.B2(n_165),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_123),
.A2(n_93),
.B1(n_105),
.B2(n_118),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_127),
.A2(n_109),
.B1(n_100),
.B2(n_104),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_144),
.B(n_108),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_109),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_122),
.A2(n_95),
.B1(n_102),
.B2(n_119),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_165),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_133),
.B(n_95),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_122),
.A2(n_107),
.B1(n_62),
.B2(n_68),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_166),
.A2(n_85),
.B1(n_61),
.B2(n_53),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_120),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_167),
.Y(n_175)
);

OA21x2_ASAP7_75t_L g168 ( 
.A1(n_121),
.A2(n_106),
.B(n_67),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_168),
.A2(n_121),
.B(n_138),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_138),
.B(n_24),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_0),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_170),
.A2(n_142),
.B(n_139),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_171),
.A2(n_173),
.B1(n_177),
.B2(n_180),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_172),
.A2(n_183),
.B(n_185),
.Y(n_212)
);

AOI22x1_ASAP7_75t_L g173 ( 
.A1(n_156),
.A2(n_137),
.B1(n_131),
.B2(n_106),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_170),
.A2(n_135),
.B(n_132),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_192),
.Y(n_205)
);

INVxp33_ASAP7_75t_L g182 ( 
.A(n_169),
.Y(n_182)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_164),
.A2(n_137),
.B1(n_131),
.B2(n_67),
.Y(n_183)
);

XNOR2x1_ASAP7_75t_L g184 ( 
.A(n_145),
.B(n_17),
.Y(n_184)
);

XNOR2x1_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_17),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_146),
.A2(n_154),
.B1(n_166),
.B2(n_152),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_162),
.A2(n_124),
.B(n_26),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_186),
.B(n_26),
.Y(n_210)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

OAI32xp33_ASAP7_75t_L g188 ( 
.A1(n_145),
.A2(n_160),
.A3(n_148),
.B1(n_168),
.B2(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_188),
.Y(n_215)
);

OAI32xp33_ASAP7_75t_L g190 ( 
.A1(n_168),
.A2(n_27),
.A3(n_23),
.B1(n_106),
.B2(n_37),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_37),
.Y(n_203)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_193),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_195),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_150),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_196),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_153),
.C(n_150),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_200),
.C(n_209),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_153),
.C(n_37),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_202),
.B(n_210),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_183),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_50),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_207),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_184),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_191),
.A2(n_61),
.B1(n_46),
.B2(n_34),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_208),
.A2(n_219),
.B1(n_192),
.B2(n_195),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_41),
.C(n_50),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_50),
.C(n_23),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_175),
.C(n_178),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_26),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_216),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_17),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_191),
.A2(n_46),
.B1(n_23),
.B2(n_3),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_176),
.B(n_23),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_173),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_181),
.Y(n_222)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_222),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_181),
.Y(n_224)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_224),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_171),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_228),
.Y(n_242)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_226),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_205),
.Y(n_227)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_227),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_215),
.A2(n_176),
.B1(n_185),
.B2(n_189),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_230),
.B(n_231),
.Y(n_244)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_206),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_232),
.B(n_235),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_186),
.C(n_174),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_236),
.C(n_209),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_202),
.A2(n_211),
.B1(n_201),
.B2(n_173),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_174),
.C(n_189),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_240),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_175),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_238),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_214),
.B(n_194),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_239),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_220),
.B(n_14),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_227),
.A2(n_203),
.B1(n_212),
.B2(n_207),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_245),
.A2(n_23),
.B1(n_2),
.B2(n_3),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_253),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_213),
.C(n_216),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_255),
.C(n_228),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_236),
.A2(n_235),
.B(n_233),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_251),
.A2(n_14),
.B(n_13),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_210),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_193),
.C(n_219),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_266),
.Y(n_275)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_265),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_221),
.C(n_229),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_262),
.C(n_263),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_249),
.A2(n_229),
.B(n_190),
.Y(n_261)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_237),
.C(n_234),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_234),
.C(n_23),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_264),
.A2(n_12),
.B(n_2),
.Y(n_276)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_241),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_13),
.C(n_12),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_1),
.C(n_2),
.Y(n_281)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_268),
.B(n_269),
.Y(n_272)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_256),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_262),
.A2(n_252),
.B(n_243),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_270),
.A2(n_4),
.B(n_5),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_257),
.A2(n_250),
.B1(n_251),
.B2(n_245),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_278),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_248),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_258),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_276),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_267),
.A2(n_247),
.B1(n_253),
.B2(n_12),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_247),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_281),
.C(n_258),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_287),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_283),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_286),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_285),
.A2(n_288),
.B(n_272),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_1),
.C(n_3),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_277),
.A2(n_4),
.B(n_5),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_6),
.C(n_7),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_291),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_6),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_275),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_292),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_273),
.C(n_280),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_295),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_297),
.A2(n_6),
.B(n_8),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_281),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_298),
.A2(n_9),
.B(n_10),
.Y(n_302)
);

NOR3xp33_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_284),
.C(n_270),
.Y(n_300)
);

O2A1O1Ixp33_ASAP7_75t_SL g305 ( 
.A1(n_300),
.A2(n_301),
.B(n_293),
.C(n_299),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_302),
.A2(n_296),
.B(n_10),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_305),
.B(n_306),
.Y(n_307)
);

OAI321xp33_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_304),
.A3(n_296),
.B1(n_303),
.B2(n_295),
.C(n_10),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_9),
.B(n_11),
.Y(n_309)
);

BUFx24_ASAP7_75t_SL g310 ( 
.A(n_309),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_11),
.B(n_308),
.Y(n_311)
);


endmodule