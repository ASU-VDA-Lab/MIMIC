module fake_netlist_6_2746_n_1851 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1851);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1851;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1669;
wire n_1403;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_181),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_115),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_92),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_63),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_130),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_54),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_171),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_140),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_126),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_7),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_119),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_10),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_106),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_2),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_38),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_148),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_13),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_135),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_97),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_88),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_120),
.Y(n_204)
);

BUFx8_ASAP7_75t_SL g205 ( 
.A(n_103),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_153),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_94),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_112),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_122),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_51),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_132),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_111),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_59),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_59),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_19),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_176),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_152),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_161),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_20),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_65),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_21),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_182),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_89),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_75),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_146),
.Y(n_226)
);

BUFx2_ASAP7_75t_SL g227 ( 
.A(n_145),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_149),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_118),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_53),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_53),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_27),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_158),
.Y(n_233)
);

BUFx5_ASAP7_75t_L g234 ( 
.A(n_73),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_174),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_109),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_57),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_7),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_42),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_15),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_179),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_82),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_99),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_147),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_25),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_101),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_169),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_104),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_125),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_134),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_93),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_40),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_151),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_167),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_79),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_31),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_17),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_78),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_155),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_177),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_100),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_175),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_15),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_28),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_44),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_129),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_71),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_156),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_87),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_128),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_56),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_139),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_50),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_10),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_136),
.Y(n_275)
);

BUFx5_ASAP7_75t_L g276 ( 
.A(n_90),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_2),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_16),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_11),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_68),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_34),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_21),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_65),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_4),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_36),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_41),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_1),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_166),
.Y(n_288)
);

BUFx10_ASAP7_75t_L g289 ( 
.A(n_47),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_43),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_98),
.Y(n_291)
);

BUFx10_ASAP7_75t_L g292 ( 
.A(n_144),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_36),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_105),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_57),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_63),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_162),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_25),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_47),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_42),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_127),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_159),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_72),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_157),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_86),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_44),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_116),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_133),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_91),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_124),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_150),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_74),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_62),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_50),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_173),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_170),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_11),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_58),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_138),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_85),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_121),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_95),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_64),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_34),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_27),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_43),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_107),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_18),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_31),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_14),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_14),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_5),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_70),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_55),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_46),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_81),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_66),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_48),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_49),
.Y(n_339)
);

BUFx8_ASAP7_75t_SL g340 ( 
.A(n_0),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_8),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_66),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_131),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_45),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_113),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_16),
.Y(n_346)
);

BUFx10_ASAP7_75t_L g347 ( 
.A(n_46),
.Y(n_347)
);

BUFx10_ASAP7_75t_L g348 ( 
.A(n_28),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_33),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_96),
.Y(n_350)
);

CKINVDCx12_ASAP7_75t_R g351 ( 
.A(n_40),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_67),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_164),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_37),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_52),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_26),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_142),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_172),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_4),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_30),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_114),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_41),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_49),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_160),
.Y(n_364)
);

BUFx10_ASAP7_75t_L g365 ( 
.A(n_45),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_102),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_222),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_340),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_232),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_270),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_191),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_222),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_338),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_222),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_323),
.B(n_1),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_222),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_222),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_222),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_225),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_188),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_294),
.B(n_303),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_222),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_288),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_324),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_214),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_222),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_220),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_236),
.Y(n_388)
);

INVxp33_ASAP7_75t_L g389 ( 
.A(n_197),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_273),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_273),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_237),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_289),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_260),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_205),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_271),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_238),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_183),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_338),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_338),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_273),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_185),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_294),
.B(n_3),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_217),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_245),
.Y(n_405)
);

NOR2xp67_ASAP7_75t_L g406 ( 
.A(n_200),
.B(n_3),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_296),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_296),
.Y(n_408)
);

INVxp33_ASAP7_75t_SL g409 ( 
.A(n_186),
.Y(n_409)
);

NOR2xp67_ASAP7_75t_L g410 ( 
.A(n_213),
.B(n_5),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_329),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_329),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_273),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_257),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_303),
.B(n_6),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_264),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_219),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_352),
.Y(n_418)
);

NOR2xp67_ASAP7_75t_L g419 ( 
.A(n_213),
.B(n_6),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_273),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_223),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_352),
.Y(n_422)
);

INVxp33_ASAP7_75t_L g423 ( 
.A(n_192),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_356),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_274),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_224),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_356),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_198),
.Y(n_428)
);

INVxp33_ASAP7_75t_SL g429 ( 
.A(n_186),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_212),
.B(n_297),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_226),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_278),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_239),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_289),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_240),
.Y(n_435)
);

INVxp67_ASAP7_75t_SL g436 ( 
.A(n_288),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_212),
.B(n_8),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_252),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_263),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_265),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_281),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_229),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_287),
.Y(n_443)
);

INVxp33_ASAP7_75t_L g444 ( 
.A(n_295),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_283),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_299),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_300),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_325),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_233),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_351),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_330),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_242),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_284),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_289),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_363),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_285),
.Y(n_456)
);

INVxp33_ASAP7_75t_L g457 ( 
.A(n_216),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_286),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_243),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_244),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_315),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_305),
.B(n_9),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_246),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_290),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_195),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_293),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_306),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_315),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_313),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_314),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_317),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_379),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_395),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_390),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_398),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_390),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_391),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_371),
.B(n_277),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_391),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_401),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_R g481 ( 
.A(n_402),
.B(n_247),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_413),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_381),
.B(n_235),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_385),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_413),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_420),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_379),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_420),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_379),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_379),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_436),
.B(n_316),
.Y(n_491)
);

BUFx8_ASAP7_75t_L g492 ( 
.A(n_465),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_400),
.B(n_316),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_404),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_373),
.B(n_297),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_417),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_421),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_426),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_388),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_379),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_367),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_369),
.B(n_292),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_372),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_461),
.B(n_231),
.Y(n_504)
);

CKINVDCx16_ASAP7_75t_R g505 ( 
.A(n_384),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_367),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_374),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_376),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_394),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_385),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_465),
.B(n_231),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_377),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_378),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_382),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_386),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_400),
.Y(n_516)
);

INVxp67_ASAP7_75t_SL g517 ( 
.A(n_383),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_428),
.Y(n_518)
);

CKINVDCx16_ASAP7_75t_R g519 ( 
.A(n_393),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_399),
.Y(n_520)
);

INVx6_ASAP7_75t_L g521 ( 
.A(n_383),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_387),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_431),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_369),
.B(n_292),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_433),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_442),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_370),
.B(n_353),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_435),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_449),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_468),
.B(n_282),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_438),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_452),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_430),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_439),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_440),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_437),
.Y(n_536)
);

INVxp67_ASAP7_75t_SL g537 ( 
.A(n_375),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_443),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_459),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_460),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_446),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_463),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_368),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_447),
.Y(n_544)
);

NAND2xp33_ASAP7_75t_L g545 ( 
.A(n_392),
.B(n_195),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_448),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_451),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_368),
.Y(n_548)
);

CKINVDCx16_ASAP7_75t_R g549 ( 
.A(n_450),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_455),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_392),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_407),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_397),
.B(n_292),
.Y(n_553)
);

NAND2xp33_ASAP7_75t_L g554 ( 
.A(n_536),
.B(n_225),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_503),
.Y(n_555)
);

INVx4_ASAP7_75t_SL g556 ( 
.A(n_536),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_537),
.B(n_408),
.Y(n_557)
);

BUFx10_ASAP7_75t_L g558 ( 
.A(n_483),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g559 ( 
.A1(n_533),
.A2(n_415),
.B1(n_403),
.B2(n_380),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_472),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_503),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_521),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_533),
.B(n_397),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_517),
.B(n_409),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_487),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_507),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_507),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_552),
.B(n_411),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_552),
.B(n_412),
.Y(n_569)
);

OR2x6_ASAP7_75t_L g570 ( 
.A(n_521),
.B(n_227),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_482),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_SL g572 ( 
.A(n_505),
.B(n_519),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_521),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_511),
.B(n_491),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_552),
.B(n_418),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_472),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_508),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_482),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_521),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_533),
.B(n_405),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_501),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_533),
.A2(n_462),
.B1(n_282),
.B2(n_419),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_553),
.B(n_429),
.Y(n_583)
);

INVxp33_ASAP7_75t_SL g584 ( 
.A(n_481),
.Y(n_584)
);

OR2x6_ASAP7_75t_L g585 ( 
.A(n_527),
.B(n_406),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_536),
.B(n_405),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_545),
.B(n_429),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_501),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_472),
.Y(n_589)
);

INVx4_ASAP7_75t_L g590 ( 
.A(n_533),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_536),
.B(n_414),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_484),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_502),
.B(n_414),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_536),
.B(n_416),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_536),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_495),
.B(n_396),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_506),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_493),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_524),
.B(n_416),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_506),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_508),
.A2(n_410),
.B1(n_221),
.B2(n_216),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_472),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_512),
.B(n_425),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_519),
.B(n_425),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_510),
.B(n_432),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_522),
.B(n_432),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_485),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_493),
.Y(n_608)
);

BUFx10_ASAP7_75t_L g609 ( 
.A(n_473),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_512),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g611 ( 
.A(n_549),
.B(n_434),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_472),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_485),
.Y(n_613)
);

BUFx4f_ASAP7_75t_L g614 ( 
.A(n_550),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_486),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_514),
.B(n_441),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_472),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_492),
.B(n_445),
.Y(n_618)
);

AO22x2_ASAP7_75t_L g619 ( 
.A1(n_504),
.A2(n_221),
.B1(n_353),
.B2(n_256),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_515),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_492),
.B(n_445),
.Y(n_621)
);

INVx1_ASAP7_75t_SL g622 ( 
.A(n_478),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_490),
.Y(n_623)
);

AND2x6_ASAP7_75t_L g624 ( 
.A(n_513),
.B(n_225),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_513),
.B(n_453),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_515),
.Y(n_626)
);

OAI22xp33_ASAP7_75t_L g627 ( 
.A1(n_549),
.A2(n_389),
.B1(n_230),
.B2(n_359),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_490),
.Y(n_628)
);

BUFx10_ASAP7_75t_L g629 ( 
.A(n_475),
.Y(n_629)
);

NAND3xp33_ASAP7_75t_L g630 ( 
.A(n_530),
.B(n_456),
.C(n_453),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_513),
.B(n_456),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_513),
.B(n_458),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_530),
.B(n_422),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_486),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_493),
.Y(n_635)
);

INVxp33_ASAP7_75t_L g636 ( 
.A(n_478),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_518),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_493),
.A2(n_424),
.B1(n_427),
.B2(n_444),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_551),
.A2(n_466),
.B1(n_470),
.B2(n_469),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_490),
.Y(n_640)
);

NAND2xp33_ASAP7_75t_R g641 ( 
.A(n_494),
.B(n_458),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_490),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_518),
.Y(n_643)
);

NOR2x1p5_ASAP7_75t_L g644 ( 
.A(n_496),
.B(n_464),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_492),
.B(n_464),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_541),
.B(n_466),
.Y(n_646)
);

BUFx10_ASAP7_75t_L g647 ( 
.A(n_497),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_541),
.B(n_467),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_489),
.B(n_467),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_520),
.B(n_457),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_550),
.A2(n_423),
.B1(n_225),
.B2(n_366),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_520),
.B(n_469),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_541),
.B(n_470),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_525),
.Y(n_654)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_538),
.B(n_454),
.Y(n_655)
);

NOR2x1p5_ASAP7_75t_L g656 ( 
.A(n_498),
.B(n_471),
.Y(n_656)
);

NAND2xp33_ASAP7_75t_L g657 ( 
.A(n_550),
.B(n_225),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_541),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_488),
.Y(n_659)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_538),
.B(n_471),
.Y(n_660)
);

INVxp67_ASAP7_75t_L g661 ( 
.A(n_492),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_544),
.B(n_184),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_544),
.B(n_187),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_488),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_499),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_474),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_476),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_550),
.A2(n_366),
.B1(n_308),
.B2(n_311),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_546),
.B(n_307),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_546),
.B(n_318),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_476),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_547),
.A2(n_534),
.B1(n_528),
.B2(n_531),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_547),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_477),
.Y(n_674)
);

INVx1_ASAP7_75t_SL g675 ( 
.A(n_509),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_528),
.B(n_193),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_500),
.B(n_302),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_490),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_523),
.B(n_307),
.Y(n_679)
);

BUFx2_ASAP7_75t_L g680 ( 
.A(n_526),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_531),
.B(n_310),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_590),
.B(n_479),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_591),
.B(n_529),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_573),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_650),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_667),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_590),
.B(n_479),
.Y(n_687)
);

INVx4_ASAP7_75t_L g688 ( 
.A(n_573),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_667),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_579),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_590),
.B(n_480),
.Y(n_691)
);

NAND2x1p5_ASAP7_75t_L g692 ( 
.A(n_595),
.B(n_194),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_574),
.B(n_563),
.Y(n_693)
);

NOR2xp67_ASAP7_75t_L g694 ( 
.A(n_639),
.B(n_630),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_598),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_SL g696 ( 
.A(n_584),
.B(n_583),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_650),
.B(n_532),
.Y(n_697)
);

BUFx8_ASAP7_75t_L g698 ( 
.A(n_680),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_594),
.B(n_558),
.Y(n_699)
);

BUFx2_ASAP7_75t_L g700 ( 
.A(n_680),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_608),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_574),
.B(n_358),
.Y(n_702)
);

NOR3xp33_ASAP7_75t_L g703 ( 
.A(n_587),
.B(n_540),
.C(n_539),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_619),
.A2(n_279),
.B1(n_355),
.B2(n_298),
.Y(n_704)
);

INVxp67_ASAP7_75t_L g705 ( 
.A(n_596),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_580),
.B(n_500),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_671),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_579),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_596),
.B(n_189),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_561),
.B(n_516),
.Y(n_710)
);

NOR3xp33_ASAP7_75t_L g711 ( 
.A(n_605),
.B(n_542),
.C(n_535),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_561),
.B(n_196),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_577),
.B(n_202),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_671),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_603),
.B(n_189),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_625),
.A2(n_632),
.B(n_631),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_619),
.A2(n_577),
.B1(n_559),
.B2(n_569),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_586),
.A2(n_254),
.B1(n_255),
.B2(n_253),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_555),
.B(n_215),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_635),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_556),
.B(n_308),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_674),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_557),
.B(n_534),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_566),
.B(n_567),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_558),
.B(n_190),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_674),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_558),
.B(n_557),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_616),
.B(n_190),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_564),
.B(n_199),
.Y(n_729)
);

INVx2_ASAP7_75t_SL g730 ( 
.A(n_652),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_660),
.B(n_199),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_610),
.B(n_218),
.Y(n_732)
);

AOI22xp5_ASAP7_75t_L g733 ( 
.A1(n_585),
.A2(n_593),
.B1(n_648),
.B2(n_646),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_635),
.Y(n_734)
);

INVxp67_ASAP7_75t_L g735 ( 
.A(n_606),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_581),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_660),
.B(n_201),
.Y(n_737)
);

INVxp67_ASAP7_75t_L g738 ( 
.A(n_611),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_652),
.B(n_201),
.Y(n_739)
);

A2O1A1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_653),
.A2(n_258),
.B(n_267),
.C(n_251),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_584),
.B(n_203),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_585),
.A2(n_269),
.B1(n_248),
.B2(n_241),
.Y(n_742)
);

AND2x4_ASAP7_75t_SL g743 ( 
.A(n_629),
.B(n_543),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_666),
.B(n_228),
.Y(n_744)
);

OR2x6_ASAP7_75t_L g745 ( 
.A(n_661),
.B(n_280),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_673),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_673),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_619),
.A2(n_339),
.B1(n_349),
.B2(n_362),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_581),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_565),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_681),
.B(n_203),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_637),
.Y(n_752)
);

OR2x2_ASAP7_75t_L g753 ( 
.A(n_655),
.B(n_210),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_643),
.Y(n_754)
);

AND2x4_ASAP7_75t_SL g755 ( 
.A(n_629),
.B(n_548),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_556),
.B(n_308),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_588),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_588),
.Y(n_758)
);

OR2x2_ASAP7_75t_L g759 ( 
.A(n_655),
.B(n_210),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_568),
.B(n_304),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_R g761 ( 
.A(n_641),
.B(n_204),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_571),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_654),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_568),
.B(n_357),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_569),
.B(n_249),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_582),
.B(n_204),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_597),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_575),
.B(n_250),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_597),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_585),
.B(n_206),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_607),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_585),
.A2(n_301),
.B1(n_364),
.B2(n_361),
.Y(n_772)
);

OAI21xp33_ASAP7_75t_L g773 ( 
.A1(n_633),
.A2(n_344),
.B(n_360),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_607),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_649),
.B(n_206),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_633),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_627),
.B(n_207),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_613),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_670),
.B(n_207),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_600),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_613),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_600),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_638),
.B(n_347),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_670),
.B(n_208),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_599),
.B(n_208),
.Y(n_785)
);

NOR2xp67_ASAP7_75t_L g786 ( 
.A(n_592),
.B(n_259),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_619),
.A2(n_366),
.B1(n_308),
.B2(n_276),
.Y(n_787)
);

A2O1A1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_620),
.A2(n_320),
.B(n_261),
.C(n_262),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_562),
.B(n_662),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_679),
.B(n_209),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_570),
.A2(n_312),
.B1(n_319),
.B2(n_321),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_662),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_554),
.A2(n_366),
.B1(n_276),
.B2(n_234),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_677),
.B(n_209),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_662),
.B(n_347),
.Y(n_795)
);

INVx4_ASAP7_75t_L g796 ( 
.A(n_658),
.Y(n_796)
);

OR2x2_ASAP7_75t_L g797 ( 
.A(n_622),
.B(n_334),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_615),
.Y(n_798)
);

NOR2xp67_ASAP7_75t_SL g799 ( 
.A(n_612),
.B(n_211),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_626),
.B(n_266),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_663),
.B(n_336),
.Y(n_801)
);

INVx3_ASAP7_75t_L g802 ( 
.A(n_571),
.Y(n_802)
);

OAI22xp5_ASAP7_75t_L g803 ( 
.A1(n_570),
.A2(n_336),
.B1(n_343),
.B2(n_345),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_669),
.B(n_343),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_614),
.A2(n_272),
.B(n_268),
.Y(n_805)
);

OAI221xp5_ASAP7_75t_L g806 ( 
.A1(n_601),
.A2(n_672),
.B1(n_651),
.B2(n_331),
.C(n_326),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_615),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_611),
.B(n_350),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_644),
.B(n_347),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_656),
.B(n_348),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_634),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_604),
.B(n_328),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_570),
.B(n_332),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_634),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_676),
.A2(n_234),
.B1(n_276),
.B2(n_354),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_659),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_730),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_735),
.B(n_665),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_693),
.B(n_676),
.Y(n_819)
);

OR2x6_ASAP7_75t_L g820 ( 
.A(n_700),
.B(n_618),
.Y(n_820)
);

AOI21x1_ASAP7_75t_L g821 ( 
.A1(n_682),
.A2(n_578),
.B(n_664),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_693),
.B(n_570),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_L g823 ( 
.A1(n_787),
.A2(n_621),
.B1(n_645),
.B2(n_668),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_716),
.A2(n_733),
.B(n_709),
.C(n_702),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_705),
.B(n_675),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_696),
.B(n_727),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_736),
.Y(n_827)
);

INVx1_ASAP7_75t_SL g828 ( 
.A(n_697),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_702),
.B(n_738),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_709),
.B(n_629),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_SL g831 ( 
.A(n_694),
.B(n_572),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_686),
.Y(n_832)
);

INVx4_ASAP7_75t_L g833 ( 
.A(n_684),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_736),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_794),
.B(n_560),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_794),
.B(n_560),
.Y(n_836)
);

INVxp67_ASAP7_75t_SL g837 ( 
.A(n_750),
.Y(n_837)
);

OAI21xp5_ASAP7_75t_L g838 ( 
.A1(n_717),
.A2(n_576),
.B(n_642),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_717),
.A2(n_576),
.B(n_642),
.Y(n_839)
);

A2O1A1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_779),
.A2(n_784),
.B(n_737),
.C(n_731),
.Y(n_840)
);

OAI21xp33_ASAP7_75t_L g841 ( 
.A1(n_731),
.A2(n_360),
.B(n_334),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_787),
.A2(n_335),
.B1(n_344),
.B2(n_346),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_704),
.A2(n_354),
.B1(n_346),
.B2(n_342),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_685),
.B(n_647),
.Y(n_844)
);

OAI321xp33_ASAP7_75t_L g845 ( 
.A1(n_704),
.A2(n_348),
.A3(n_365),
.B1(n_337),
.B2(n_341),
.C(n_342),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_715),
.B(n_636),
.Y(n_846)
);

BUFx12f_ASAP7_75t_L g847 ( 
.A(n_698),
.Y(n_847)
);

INVxp67_ASAP7_75t_L g848 ( 
.A(n_737),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_775),
.B(n_576),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_689),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_715),
.A2(n_628),
.B1(n_589),
.B2(n_602),
.Y(n_851)
);

O2A1O1Ixp5_ASAP7_75t_SL g852 ( 
.A1(n_699),
.A2(n_642),
.B(n_628),
.C(n_602),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_775),
.B(n_589),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_779),
.B(n_784),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_752),
.B(n_589),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_792),
.A2(n_333),
.B1(n_309),
.B2(n_275),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_743),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_754),
.B(n_612),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_729),
.B(n_797),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_760),
.A2(n_657),
.B(n_624),
.Y(n_860)
);

NOR2x1_ASAP7_75t_L g861 ( 
.A(n_683),
.B(n_684),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_707),
.Y(n_862)
);

OAI21xp5_ASAP7_75t_L g863 ( 
.A1(n_764),
.A2(n_624),
.B(n_291),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_707),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_749),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_789),
.Y(n_866)
);

AO22x1_ASAP7_75t_L g867 ( 
.A1(n_790),
.A2(n_636),
.B1(n_337),
.B2(n_335),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_763),
.B(n_678),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_695),
.A2(n_322),
.B1(n_327),
.B2(n_624),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_776),
.B(n_647),
.Y(n_870)
);

INVx4_ASAP7_75t_L g871 ( 
.A(n_690),
.Y(n_871)
);

INVx6_ASAP7_75t_L g872 ( 
.A(n_809),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_783),
.B(n_647),
.Y(n_873)
);

O2A1O1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_728),
.A2(n_307),
.B(n_341),
.C(n_365),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_690),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_714),
.A2(n_624),
.B(n_640),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_749),
.Y(n_877)
);

AO21x1_ASAP7_75t_L g878 ( 
.A1(n_692),
.A2(n_234),
.B(n_276),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_708),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_748),
.A2(n_815),
.B1(n_793),
.B2(n_785),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_714),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_722),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_747),
.B(n_609),
.Y(n_883)
);

O2A1O1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_788),
.A2(n_624),
.B(n_12),
.C(n_13),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_757),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_757),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_708),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_722),
.Y(n_888)
);

A2O1A1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_785),
.A2(n_623),
.B(n_617),
.C(n_565),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_726),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_747),
.B(n_609),
.Y(n_891)
);

NOR3xp33_ASAP7_75t_L g892 ( 
.A(n_790),
.B(n_609),
.C(n_12),
.Y(n_892)
);

BUFx12f_ASAP7_75t_L g893 ( 
.A(n_745),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_724),
.A2(n_276),
.B(n_234),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_789),
.A2(n_276),
.B(n_234),
.Y(n_895)
);

NOR2xp67_ASAP7_75t_L g896 ( 
.A(n_772),
.B(n_69),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_726),
.B(n_276),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_744),
.A2(n_234),
.B(n_180),
.Y(n_898)
);

INVx4_ASAP7_75t_L g899 ( 
.A(n_796),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_765),
.B(n_234),
.Y(n_900)
);

OAI321xp33_ASAP7_75t_L g901 ( 
.A1(n_748),
.A2(n_9),
.A3(n_17),
.B1(n_18),
.B2(n_19),
.C(n_22),
.Y(n_901)
);

A2O1A1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_812),
.A2(n_770),
.B(n_804),
.C(n_813),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_761),
.B(n_234),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_812),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_768),
.B(n_23),
.Y(n_905)
);

AO21x1_ASAP7_75t_L g906 ( 
.A1(n_692),
.A2(n_24),
.B(n_26),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_770),
.A2(n_29),
.B(n_30),
.C(n_32),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_758),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_798),
.B(n_80),
.Y(n_909)
);

AOI21x1_ASAP7_75t_L g910 ( 
.A1(n_710),
.A2(n_756),
.B(n_721),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_725),
.B(n_32),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_798),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_758),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_807),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_800),
.A2(n_83),
.B(n_178),
.Y(n_915)
);

O2A1O1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_712),
.A2(n_33),
.B(n_35),
.C(n_37),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_767),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_688),
.Y(n_918)
);

BUFx2_ASAP7_75t_L g919 ( 
.A(n_761),
.Y(n_919)
);

BUFx12f_ASAP7_75t_L g920 ( 
.A(n_745),
.Y(n_920)
);

BUFx12f_ASAP7_75t_L g921 ( 
.A(n_745),
.Y(n_921)
);

A2O1A1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_804),
.A2(n_35),
.B(n_38),
.C(n_39),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_807),
.B(n_84),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_746),
.B(n_39),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_753),
.Y(n_925)
);

NOR3xp33_ASAP7_75t_L g926 ( 
.A(n_741),
.B(n_48),
.C(n_52),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_777),
.B(n_54),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_813),
.A2(n_55),
.B(n_56),
.C(n_58),
.Y(n_928)
);

A2O1A1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_701),
.A2(n_734),
.B(n_720),
.C(n_814),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_688),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_795),
.B(n_117),
.Y(n_931)
);

NAND3xp33_ASAP7_75t_L g932 ( 
.A(n_711),
.B(n_60),
.C(n_61),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_816),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_808),
.B(n_61),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_771),
.A2(n_123),
.B(n_163),
.Y(n_935)
);

O2A1O1Ixp5_ASAP7_75t_L g936 ( 
.A1(n_751),
.A2(n_110),
.B(n_154),
.C(n_143),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_810),
.B(n_77),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_774),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_762),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_778),
.A2(n_108),
.B(n_141),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_767),
.A2(n_76),
.B(n_137),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_781),
.B(n_62),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_811),
.B(n_64),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_769),
.A2(n_782),
.B(n_780),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_742),
.B(n_67),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_739),
.B(n_759),
.Y(n_946)
);

OAI21x1_ASAP7_75t_L g947 ( 
.A1(n_802),
.A2(n_782),
.B(n_756),
.Y(n_947)
);

OAI22xp5_ASAP7_75t_L g948 ( 
.A1(n_815),
.A2(n_793),
.B1(n_713),
.B2(n_806),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_719),
.A2(n_732),
.B1(n_766),
.B2(n_791),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_786),
.B(n_773),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_801),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_718),
.B(n_703),
.Y(n_952)
);

OAI21xp33_ASAP7_75t_L g953 ( 
.A1(n_803),
.A2(n_740),
.B(n_743),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_805),
.B(n_799),
.Y(n_954)
);

INVx4_ASAP7_75t_L g955 ( 
.A(n_755),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_755),
.B(n_705),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_706),
.A2(n_590),
.B(n_595),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_705),
.B(n_702),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_686),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_686),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_736),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_706),
.A2(n_590),
.B(n_595),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_693),
.B(n_723),
.Y(n_963)
);

AOI21x1_ASAP7_75t_L g964 ( 
.A1(n_682),
.A2(n_691),
.B(n_687),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_693),
.B(n_723),
.Y(n_965)
);

A2O1A1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_693),
.A2(n_716),
.B(n_733),
.C(n_709),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_684),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_956),
.Y(n_968)
);

NAND2x1p5_ASAP7_75t_L g969 ( 
.A(n_930),
.B(n_918),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_963),
.B(n_965),
.Y(n_970)
);

AOI221xp5_ASAP7_75t_SL g971 ( 
.A1(n_880),
.A2(n_840),
.B1(n_902),
.B2(n_854),
.C(n_927),
.Y(n_971)
);

OAI21x1_ASAP7_75t_L g972 ( 
.A1(n_947),
.A2(n_944),
.B(n_821),
.Y(n_972)
);

AOI21x1_ASAP7_75t_L g973 ( 
.A1(n_849),
.A2(n_853),
.B(n_836),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_958),
.B(n_828),
.Y(n_974)
);

OAI22x1_ASAP7_75t_L g975 ( 
.A1(n_846),
.A2(n_848),
.B1(n_911),
.B2(n_829),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_966),
.B(n_824),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_832),
.Y(n_977)
);

AOI21x1_ASAP7_75t_L g978 ( 
.A1(n_835),
.A2(n_964),
.B(n_900),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_918),
.Y(n_979)
);

AOI21x1_ASAP7_75t_L g980 ( 
.A1(n_957),
.A2(n_962),
.B(n_954),
.Y(n_980)
);

AO21x1_ASAP7_75t_L g981 ( 
.A1(n_898),
.A2(n_880),
.B(n_823),
.Y(n_981)
);

AO31x2_ASAP7_75t_L g982 ( 
.A1(n_889),
.A2(n_878),
.A3(n_948),
.B(n_906),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_948),
.A2(n_819),
.B1(n_823),
.B2(n_822),
.Y(n_983)
);

AO21x2_ASAP7_75t_L g984 ( 
.A1(n_863),
.A2(n_898),
.B(n_860),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_828),
.B(n_873),
.Y(n_985)
);

CKINVDCx8_ASAP7_75t_R g986 ( 
.A(n_919),
.Y(n_986)
);

NAND2x1p5_ASAP7_75t_L g987 ( 
.A(n_930),
.B(n_918),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_857),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_850),
.Y(n_989)
);

AO221x1_ASAP7_75t_L g990 ( 
.A1(n_843),
.A2(n_842),
.B1(n_949),
.B2(n_845),
.C(n_901),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_862),
.B(n_864),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_830),
.B(n_831),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_847),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_852),
.A2(n_839),
.B(n_838),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_881),
.B(n_882),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_888),
.B(n_890),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_912),
.B(n_914),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_925),
.B(n_818),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_825),
.B(n_831),
.Y(n_999)
);

AOI21x1_ASAP7_75t_L g1000 ( 
.A1(n_910),
.A2(n_923),
.B(n_909),
.Y(n_1000)
);

OA22x2_ASAP7_75t_L g1001 ( 
.A1(n_843),
.A2(n_842),
.B1(n_820),
.B2(n_951),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_959),
.B(n_960),
.Y(n_1002)
);

NOR2x1_ASAP7_75t_SL g1003 ( 
.A(n_933),
.B(n_899),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_905),
.B(n_938),
.Y(n_1004)
);

INVx2_ASAP7_75t_SL g1005 ( 
.A(n_817),
.Y(n_1005)
);

CKINVDCx8_ASAP7_75t_R g1006 ( 
.A(n_875),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_827),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_934),
.A2(n_946),
.B(n_859),
.C(n_826),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_834),
.B(n_865),
.Y(n_1009)
);

INVx1_ASAP7_75t_SL g1010 ( 
.A(n_870),
.Y(n_1010)
);

AO31x2_ASAP7_75t_L g1011 ( 
.A1(n_929),
.A2(n_904),
.A3(n_923),
.B(n_909),
.Y(n_1011)
);

AOI21xp33_ASAP7_75t_L g1012 ( 
.A1(n_952),
.A2(n_901),
.B(n_841),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_877),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_885),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_886),
.B(n_908),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_931),
.A2(n_839),
.B1(n_922),
.B2(n_928),
.Y(n_1016)
);

BUFx12f_ASAP7_75t_L g1017 ( 
.A(n_955),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_913),
.B(n_917),
.Y(n_1018)
);

BUFx3_ASAP7_75t_L g1019 ( 
.A(n_955),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_937),
.B(n_950),
.Y(n_1020)
);

OR2x6_ASAP7_75t_L g1021 ( 
.A(n_820),
.B(n_893),
.Y(n_1021)
);

AOI21x1_ASAP7_75t_L g1022 ( 
.A1(n_897),
.A2(n_858),
.B(n_868),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_961),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_933),
.B(n_866),
.Y(n_1024)
);

AOI21x1_ASAP7_75t_L g1025 ( 
.A1(n_855),
.A2(n_943),
.B(n_942),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_933),
.B(n_866),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_939),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_939),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_931),
.B(n_937),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_876),
.A2(n_895),
.B(n_851),
.Y(n_1030)
);

OA21x2_ASAP7_75t_L g1031 ( 
.A1(n_941),
.A2(n_894),
.B(n_936),
.Y(n_1031)
);

OAI21xp33_ASAP7_75t_L g1032 ( 
.A1(n_926),
.A2(n_892),
.B(n_924),
.Y(n_1032)
);

AOI21x1_ASAP7_75t_L g1033 ( 
.A1(n_903),
.A2(n_861),
.B(n_915),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_875),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_837),
.A2(n_953),
.B(n_884),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_879),
.B(n_967),
.Y(n_1036)
);

O2A1O1Ixp5_ASAP7_75t_L g1037 ( 
.A1(n_883),
.A2(n_891),
.B(n_945),
.C(n_940),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_967),
.Y(n_1038)
);

OAI22x1_ASAP7_75t_L g1039 ( 
.A1(n_932),
.A2(n_845),
.B1(n_844),
.B2(n_833),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_879),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_872),
.A2(n_896),
.B1(n_856),
.B2(n_820),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_907),
.A2(n_869),
.B(n_935),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_887),
.B(n_967),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_887),
.Y(n_1044)
);

AOI21xp33_ASAP7_75t_L g1045 ( 
.A1(n_874),
.A2(n_916),
.B(n_899),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_833),
.A2(n_871),
.B(n_867),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_872),
.A2(n_871),
.B(n_920),
.C(n_921),
.Y(n_1047)
);

OR2x6_ASAP7_75t_L g1048 ( 
.A(n_955),
.B(n_857),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_918),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_958),
.B(n_705),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_963),
.B(n_965),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_947),
.A2(n_944),
.B(n_821),
.Y(n_1052)
);

AOI21x1_ASAP7_75t_L g1053 ( 
.A1(n_821),
.A2(n_853),
.B(n_849),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_875),
.B(n_967),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_963),
.B(n_965),
.Y(n_1055)
);

AO21x1_ASAP7_75t_L g1056 ( 
.A1(n_854),
.A2(n_898),
.B(n_880),
.Y(n_1056)
);

INVx4_ASAP7_75t_L g1057 ( 
.A(n_918),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_958),
.B(n_705),
.Y(n_1058)
);

AND2x6_ASAP7_75t_L g1059 ( 
.A(n_931),
.B(n_937),
.Y(n_1059)
);

AO31x2_ASAP7_75t_L g1060 ( 
.A1(n_889),
.A2(n_878),
.A3(n_966),
.B(n_824),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_947),
.A2(n_944),
.B(n_821),
.Y(n_1061)
);

AO31x2_ASAP7_75t_L g1062 ( 
.A1(n_889),
.A2(n_878),
.A3(n_966),
.B(n_824),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_880),
.A2(n_840),
.B1(n_854),
.B2(n_963),
.Y(n_1063)
);

INVx2_ASAP7_75t_SL g1064 ( 
.A(n_817),
.Y(n_1064)
);

AOI21x1_ASAP7_75t_L g1065 ( 
.A1(n_821),
.A2(n_853),
.B(n_849),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_963),
.B(n_965),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_947),
.A2(n_944),
.B(n_821),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_947),
.A2(n_944),
.B(n_821),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_832),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_875),
.B(n_967),
.Y(n_1070)
);

AO31x2_ASAP7_75t_L g1071 ( 
.A1(n_889),
.A2(n_878),
.A3(n_966),
.B(n_824),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_966),
.A2(n_840),
.B(n_824),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_847),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_L g1074 ( 
.A1(n_947),
.A2(n_944),
.B(n_821),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_854),
.A2(n_840),
.B1(n_846),
.B2(n_831),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_854),
.B(n_848),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_963),
.B(n_965),
.Y(n_1077)
);

AND2x6_ASAP7_75t_L g1078 ( 
.A(n_931),
.B(n_937),
.Y(n_1078)
);

AOI21xp33_ASAP7_75t_L g1079 ( 
.A1(n_854),
.A2(n_880),
.B(n_840),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_854),
.B(n_848),
.Y(n_1080)
);

INVx3_ASAP7_75t_SL g1081 ( 
.A(n_955),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_827),
.Y(n_1082)
);

AOI21x1_ASAP7_75t_L g1083 ( 
.A1(n_821),
.A2(n_853),
.B(n_849),
.Y(n_1083)
);

AO31x2_ASAP7_75t_L g1084 ( 
.A1(n_889),
.A2(n_878),
.A3(n_966),
.B(n_824),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_847),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_947),
.A2(n_944),
.B(n_821),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_848),
.B(n_735),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_848),
.B(n_735),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_947),
.A2(n_944),
.B(n_821),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_963),
.B(n_965),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_854),
.B(n_848),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_958),
.B(n_705),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_956),
.Y(n_1093)
);

AO21x1_ASAP7_75t_L g1094 ( 
.A1(n_854),
.A2(n_898),
.B(n_880),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_827),
.Y(n_1095)
);

BUFx2_ASAP7_75t_L g1096 ( 
.A(n_956),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_958),
.B(n_705),
.Y(n_1097)
);

HAxp5_ASAP7_75t_L g1098 ( 
.A(n_1087),
.B(n_1088),
.CON(n_1098),
.SN(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1007),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_968),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_977),
.Y(n_1101)
);

INVx4_ASAP7_75t_L g1102 ( 
.A(n_979),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_989),
.Y(n_1103)
);

OR2x2_ASAP7_75t_L g1104 ( 
.A(n_974),
.B(n_1050),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1069),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_1054),
.B(n_1070),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_1006),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_1075),
.A2(n_1077),
.B1(n_970),
.B2(n_1051),
.Y(n_1108)
);

AND2x6_ASAP7_75t_L g1109 ( 
.A(n_979),
.B(n_1049),
.Y(n_1109)
);

BUFx5_ASAP7_75t_L g1110 ( 
.A(n_1027),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_1093),
.Y(n_1111)
);

BUFx10_ASAP7_75t_L g1112 ( 
.A(n_1054),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1058),
.B(n_1092),
.Y(n_1113)
);

INVx6_ASAP7_75t_L g1114 ( 
.A(n_1017),
.Y(n_1114)
);

INVxp67_ASAP7_75t_L g1115 ( 
.A(n_998),
.Y(n_1115)
);

INVx1_ASAP7_75t_SL g1116 ( 
.A(n_985),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_979),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_999),
.A2(n_971),
.B1(n_1063),
.B2(n_990),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_L g1119 ( 
.A1(n_1001),
.A2(n_1012),
.B1(n_981),
.B2(n_1056),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_991),
.Y(n_1120)
);

HB1xp67_ASAP7_75t_L g1121 ( 
.A(n_1005),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_SL g1122 ( 
.A(n_1012),
.B(n_1008),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_988),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_1096),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_991),
.Y(n_1125)
);

BUFx12f_ASAP7_75t_L g1126 ( 
.A(n_1073),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1097),
.B(n_1020),
.Y(n_1127)
);

INVx5_ASAP7_75t_L g1128 ( 
.A(n_1049),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_1064),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_995),
.Y(n_1130)
);

NAND3xp33_ASAP7_75t_L g1131 ( 
.A(n_1079),
.B(n_1072),
.C(n_1063),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_1044),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_995),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_1076),
.B(n_1080),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_970),
.A2(n_1055),
.B1(n_1066),
.B2(n_1090),
.Y(n_1135)
);

OR2x6_ASAP7_75t_L g1136 ( 
.A(n_1048),
.B(n_1021),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1082),
.Y(n_1137)
);

HB1xp67_ASAP7_75t_L g1138 ( 
.A(n_1010),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_996),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1051),
.B(n_1055),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1066),
.A2(n_1077),
.B1(n_1090),
.B2(n_1016),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1001),
.A2(n_1094),
.B1(n_1079),
.B2(n_1032),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_996),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_997),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_1010),
.Y(n_1145)
);

CKINVDCx8_ASAP7_75t_R g1146 ( 
.A(n_1085),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_1034),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_1070),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_997),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1091),
.B(n_1004),
.Y(n_1150)
);

NAND2x1p5_ASAP7_75t_L g1151 ( 
.A(n_1057),
.B(n_1049),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1016),
.A2(n_976),
.B1(n_1072),
.B2(n_1029),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1059),
.B(n_1078),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_1034),
.Y(n_1154)
);

BUFx12f_ASAP7_75t_L g1155 ( 
.A(n_993),
.Y(n_1155)
);

INVxp67_ASAP7_75t_SL g1156 ( 
.A(n_969),
.Y(n_1156)
);

BUFx12f_ASAP7_75t_L g1157 ( 
.A(n_1034),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1004),
.B(n_976),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_1036),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_983),
.B(n_1059),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1048),
.B(n_1038),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1059),
.B(n_1078),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1002),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_986),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_975),
.B(n_992),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1036),
.B(n_1043),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_1021),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_983),
.B(n_1059),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1078),
.B(n_1002),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1081),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_1029),
.B(n_1041),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1078),
.B(n_1024),
.Y(n_1172)
);

NAND3xp33_ASAP7_75t_L g1173 ( 
.A(n_1042),
.B(n_1035),
.C(n_1045),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1042),
.A2(n_1037),
.B(n_1045),
.C(n_1046),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1013),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1014),
.Y(n_1176)
);

AOI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_984),
.A2(n_1039),
.B1(n_1021),
.B2(n_1023),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_1019),
.Y(n_1178)
);

OR2x2_ASAP7_75t_SL g1179 ( 
.A(n_1043),
.B(n_1040),
.Y(n_1179)
);

OA21x2_ASAP7_75t_L g1180 ( 
.A1(n_972),
.A2(n_1074),
.B(n_1068),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1024),
.B(n_1026),
.Y(n_1181)
);

OR2x6_ASAP7_75t_L g1182 ( 
.A(n_1046),
.B(n_1047),
.Y(n_1182)
);

INVx4_ASAP7_75t_L g1183 ( 
.A(n_969),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_1026),
.B(n_1028),
.Y(n_1184)
);

NAND3xp33_ASAP7_75t_L g1185 ( 
.A(n_994),
.B(n_1031),
.C(n_1095),
.Y(n_1185)
);

AND2x2_ASAP7_75t_SL g1186 ( 
.A(n_1031),
.B(n_1009),
.Y(n_1186)
);

AOI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1009),
.A2(n_1015),
.B1(n_1018),
.B2(n_994),
.Y(n_1187)
);

INVx4_ASAP7_75t_L g1188 ( 
.A(n_987),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_987),
.Y(n_1189)
);

OA21x2_ASAP7_75t_L g1190 ( 
.A1(n_1052),
.A2(n_1089),
.B(n_1086),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1015),
.B(n_1018),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_1025),
.B(n_1033),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1084),
.B(n_1060),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1003),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_973),
.A2(n_1022),
.B1(n_978),
.B2(n_1000),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_982),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1060),
.B(n_1084),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1060),
.B(n_1084),
.Y(n_1198)
);

OR2x2_ASAP7_75t_L g1199 ( 
.A(n_1011),
.B(n_982),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_982),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_1062),
.Y(n_1201)
);

INVx3_ASAP7_75t_SL g1202 ( 
.A(n_1011),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1030),
.B(n_1083),
.Y(n_1203)
);

INVx5_ASAP7_75t_L g1204 ( 
.A(n_1062),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1011),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_SL g1206 ( 
.A1(n_1071),
.A2(n_1062),
.B1(n_1065),
.B2(n_1053),
.Y(n_1206)
);

OR2x2_ASAP7_75t_L g1207 ( 
.A(n_1071),
.B(n_1061),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_1071),
.B(n_980),
.Y(n_1208)
);

OAI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1067),
.A2(n_854),
.B1(n_696),
.B2(n_1075),
.Y(n_1209)
);

OR2x2_ASAP7_75t_L g1210 ( 
.A(n_974),
.B(n_705),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1007),
.Y(n_1211)
);

NAND2xp33_ASAP7_75t_L g1212 ( 
.A(n_1059),
.B(n_840),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_970),
.B(n_1051),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_974),
.B(n_958),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_999),
.B(n_828),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_974),
.B(n_958),
.Y(n_1216)
);

OR2x2_ASAP7_75t_L g1217 ( 
.A(n_974),
.B(n_705),
.Y(n_1217)
);

BUFx3_ASAP7_75t_L g1218 ( 
.A(n_1006),
.Y(n_1218)
);

BUFx2_ASAP7_75t_L g1219 ( 
.A(n_968),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_974),
.B(n_958),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_970),
.B(n_1051),
.Y(n_1221)
);

AOI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1075),
.A2(n_854),
.B1(n_880),
.B2(n_999),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_SL g1223 ( 
.A1(n_976),
.A2(n_966),
.B(n_824),
.Y(n_1223)
);

INVxp67_ASAP7_75t_L g1224 ( 
.A(n_998),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1054),
.B(n_1070),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_1006),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_970),
.B(n_1051),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_970),
.B(n_1051),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_970),
.B(n_1051),
.Y(n_1229)
);

NAND2x1p5_ASAP7_75t_L g1230 ( 
.A(n_1057),
.B(n_979),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1075),
.A2(n_880),
.B1(n_840),
.B2(n_854),
.Y(n_1231)
);

AOI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1075),
.A2(n_854),
.B1(n_880),
.B2(n_999),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_977),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_974),
.B(n_958),
.Y(n_1234)
);

INVx3_ASAP7_75t_L g1235 ( 
.A(n_979),
.Y(n_1235)
);

NOR2x1_ASAP7_75t_L g1236 ( 
.A(n_1057),
.B(n_680),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_1054),
.B(n_1070),
.Y(n_1237)
);

NOR2x1_ASAP7_75t_SL g1238 ( 
.A(n_992),
.B(n_918),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_SL g1239 ( 
.A1(n_1072),
.A2(n_846),
.B(n_587),
.C(n_593),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1231),
.A2(n_1131),
.B1(n_1122),
.B2(n_1232),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1101),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1103),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1105),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_1126),
.Y(n_1244)
);

BUFx2_ASAP7_75t_R g1245 ( 
.A(n_1146),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1221),
.B(n_1140),
.Y(n_1246)
);

INVx6_ASAP7_75t_L g1247 ( 
.A(n_1107),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1113),
.B(n_1127),
.Y(n_1248)
);

HB1xp67_ASAP7_75t_L g1249 ( 
.A(n_1204),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1222),
.A2(n_1232),
.B(n_1231),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1233),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_SL g1252 ( 
.A1(n_1122),
.A2(n_1131),
.B1(n_1152),
.B2(n_1173),
.Y(n_1252)
);

AOI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1171),
.A2(n_1222),
.B1(n_1165),
.B2(n_1215),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1175),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_1204),
.Y(n_1255)
);

INVx2_ASAP7_75t_SL g1256 ( 
.A(n_1107),
.Y(n_1256)
);

INVx3_ASAP7_75t_L g1257 ( 
.A(n_1183),
.Y(n_1257)
);

INVx5_ASAP7_75t_L g1258 ( 
.A(n_1109),
.Y(n_1258)
);

INVx1_ASAP7_75t_SL g1259 ( 
.A(n_1100),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_1111),
.Y(n_1260)
);

AOI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1203),
.A2(n_1192),
.B(n_1195),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1176),
.Y(n_1262)
);

BUFx10_ASAP7_75t_L g1263 ( 
.A(n_1107),
.Y(n_1263)
);

BUFx12f_ASAP7_75t_L g1264 ( 
.A(n_1226),
.Y(n_1264)
);

BUFx10_ASAP7_75t_L g1265 ( 
.A(n_1226),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1173),
.A2(n_1152),
.B1(n_1142),
.B2(n_1118),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1099),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_SL g1268 ( 
.A1(n_1141),
.A2(n_1212),
.B1(n_1108),
.B2(n_1135),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1140),
.B(n_1213),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1118),
.A2(n_1141),
.B1(n_1108),
.B2(n_1135),
.Y(n_1270)
);

INVx2_ASAP7_75t_SL g1271 ( 
.A(n_1226),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1191),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_1123),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_SL g1274 ( 
.A1(n_1213),
.A2(n_1228),
.B1(n_1227),
.B2(n_1229),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1128),
.Y(n_1275)
);

AO21x1_ASAP7_75t_L g1276 ( 
.A1(n_1209),
.A2(n_1160),
.B(n_1168),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1119),
.A2(n_1227),
.B1(n_1228),
.B2(n_1229),
.Y(n_1277)
);

BUFx2_ASAP7_75t_R g1278 ( 
.A(n_1218),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_SL g1279 ( 
.A1(n_1134),
.A2(n_1116),
.B1(n_1214),
.B2(n_1216),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1157),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_1170),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_SL g1282 ( 
.A1(n_1116),
.A2(n_1234),
.B1(n_1220),
.B2(n_1160),
.Y(n_1282)
);

INVx2_ASAP7_75t_SL g1283 ( 
.A(n_1114),
.Y(n_1283)
);

CKINVDCx6p67_ASAP7_75t_R g1284 ( 
.A(n_1155),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1150),
.A2(n_1158),
.B1(n_1168),
.B2(n_1104),
.Y(n_1285)
);

CKINVDCx6p67_ASAP7_75t_R g1286 ( 
.A(n_1164),
.Y(n_1286)
);

INVx1_ASAP7_75t_SL g1287 ( 
.A(n_1124),
.Y(n_1287)
);

AOI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1136),
.A2(n_1115),
.B1(n_1224),
.B2(n_1236),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1150),
.A2(n_1158),
.B1(n_1125),
.B2(n_1144),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1137),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1120),
.A2(n_1139),
.B1(n_1143),
.B2(n_1163),
.Y(n_1291)
);

OR2x2_ASAP7_75t_L g1292 ( 
.A(n_1210),
.B(n_1217),
.Y(n_1292)
);

INVx2_ASAP7_75t_SL g1293 ( 
.A(n_1114),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1130),
.A2(n_1133),
.B1(n_1149),
.B2(n_1145),
.Y(n_1294)
);

AOI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1136),
.A2(n_1167),
.B1(n_1182),
.B2(n_1178),
.Y(n_1295)
);

AOI21xp33_ASAP7_75t_SL g1296 ( 
.A1(n_1136),
.A2(n_1129),
.B(n_1121),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1138),
.A2(n_1182),
.B1(n_1196),
.B2(n_1211),
.Y(n_1297)
);

CKINVDCx11_ASAP7_75t_R g1298 ( 
.A(n_1112),
.Y(n_1298)
);

BUFx6f_ASAP7_75t_L g1299 ( 
.A(n_1128),
.Y(n_1299)
);

BUFx2_ASAP7_75t_R g1300 ( 
.A(n_1153),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1204),
.Y(n_1301)
);

AO21x1_ASAP7_75t_SL g1302 ( 
.A1(n_1200),
.A2(n_1193),
.B(n_1197),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_1106),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1181),
.Y(n_1304)
);

HB1xp67_ASAP7_75t_L g1305 ( 
.A(n_1181),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1166),
.B(n_1239),
.Y(n_1306)
);

BUFx8_ASAP7_75t_L g1307 ( 
.A(n_1219),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_SL g1308 ( 
.A1(n_1098),
.A2(n_1238),
.B1(n_1201),
.B2(n_1223),
.Y(n_1308)
);

BUFx2_ASAP7_75t_R g1309 ( 
.A(n_1162),
.Y(n_1309)
);

OA21x2_ASAP7_75t_L g1310 ( 
.A1(n_1174),
.A2(n_1185),
.B(n_1205),
.Y(n_1310)
);

AND2x4_ASAP7_75t_L g1311 ( 
.A(n_1225),
.B(n_1237),
.Y(n_1311)
);

INVx11_ASAP7_75t_L g1312 ( 
.A(n_1109),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1166),
.B(n_1159),
.Y(n_1313)
);

CKINVDCx11_ASAP7_75t_R g1314 ( 
.A(n_1112),
.Y(n_1314)
);

NAND2x1p5_ASAP7_75t_L g1315 ( 
.A(n_1188),
.B(n_1161),
.Y(n_1315)
);

BUFx8_ASAP7_75t_L g1316 ( 
.A(n_1132),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_SL g1317 ( 
.A1(n_1177),
.A2(n_1169),
.B(n_1172),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1179),
.A2(n_1177),
.B1(n_1169),
.B2(n_1172),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1207),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1237),
.B(n_1148),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1208),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_1147),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1117),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1202),
.A2(n_1206),
.B1(n_1199),
.B2(n_1184),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1187),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1189),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1206),
.A2(n_1198),
.B1(n_1186),
.B2(n_1194),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1156),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1154),
.B(n_1235),
.Y(n_1329)
);

INVx3_ASAP7_75t_L g1330 ( 
.A(n_1102),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1110),
.Y(n_1331)
);

CKINVDCx20_ASAP7_75t_R g1332 ( 
.A(n_1117),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1117),
.B(n_1230),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1109),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1110),
.Y(n_1335)
);

BUFx2_ASAP7_75t_SL g1336 ( 
.A(n_1109),
.Y(n_1336)
);

INVx6_ASAP7_75t_L g1337 ( 
.A(n_1151),
.Y(n_1337)
);

AND2x4_ASAP7_75t_L g1338 ( 
.A(n_1151),
.B(n_1230),
.Y(n_1338)
);

NAND2x1p5_ASAP7_75t_L g1339 ( 
.A(n_1180),
.B(n_1190),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1101),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_SL g1341 ( 
.A1(n_1122),
.A2(n_990),
.B1(n_880),
.B2(n_999),
.Y(n_1341)
);

OR2x6_ASAP7_75t_L g1342 ( 
.A(n_1136),
.B(n_1182),
.Y(n_1342)
);

INVx11_ASAP7_75t_L g1343 ( 
.A(n_1157),
.Y(n_1343)
);

INVx1_ASAP7_75t_SL g1344 ( 
.A(n_1113),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1101),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1113),
.B(n_1127),
.Y(n_1346)
);

AO21x1_ASAP7_75t_L g1347 ( 
.A1(n_1122),
.A2(n_854),
.B(n_1231),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_SL g1348 ( 
.A1(n_1122),
.A2(n_990),
.B1(n_880),
.B2(n_999),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1101),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1101),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1221),
.B(n_1140),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_1146),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1204),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1113),
.B(n_1127),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1101),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1101),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1122),
.A2(n_990),
.B1(n_880),
.B2(n_999),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1215),
.B(n_854),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1101),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1204),
.Y(n_1360)
);

BUFx2_ASAP7_75t_R g1361 ( 
.A(n_1146),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1101),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1101),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1101),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1100),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1101),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1231),
.A2(n_990),
.B1(n_854),
.B2(n_880),
.Y(n_1367)
);

INVx3_ASAP7_75t_L g1368 ( 
.A(n_1183),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1342),
.B(n_1321),
.Y(n_1369)
);

INVx2_ASAP7_75t_SL g1370 ( 
.A(n_1337),
.Y(n_1370)
);

BUFx12f_ASAP7_75t_L g1371 ( 
.A(n_1263),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1250),
.B(n_1319),
.Y(n_1372)
);

AO21x1_ASAP7_75t_SL g1373 ( 
.A1(n_1270),
.A2(n_1240),
.B(n_1266),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1339),
.Y(n_1374)
);

INVx4_ASAP7_75t_SL g1375 ( 
.A(n_1342),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1246),
.B(n_1351),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_1342),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1325),
.Y(n_1378)
);

BUFx4f_ASAP7_75t_L g1379 ( 
.A(n_1315),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1310),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1240),
.B(n_1252),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1252),
.B(n_1272),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1310),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1310),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1306),
.B(n_1270),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1272),
.B(n_1268),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1269),
.B(n_1358),
.Y(n_1387)
);

INVxp67_ASAP7_75t_L g1388 ( 
.A(n_1248),
.Y(n_1388)
);

OR2x6_ASAP7_75t_L g1389 ( 
.A(n_1317),
.B(n_1318),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1358),
.B(n_1304),
.Y(n_1390)
);

OAI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1268),
.A2(n_1348),
.B(n_1341),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1261),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1266),
.B(n_1305),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1331),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1335),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1249),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1305),
.Y(n_1397)
);

OR2x6_ASAP7_75t_L g1398 ( 
.A(n_1276),
.B(n_1347),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1285),
.B(n_1253),
.Y(n_1399)
);

INVx1_ASAP7_75t_SL g1400 ( 
.A(n_1313),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1341),
.B(n_1348),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1357),
.B(n_1274),
.Y(n_1402)
);

BUFx12f_ASAP7_75t_L g1403 ( 
.A(n_1263),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1328),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1241),
.Y(n_1405)
);

INVx3_ASAP7_75t_L g1406 ( 
.A(n_1258),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1242),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1243),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1251),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1357),
.B(n_1274),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1340),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1345),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1277),
.B(n_1285),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1349),
.Y(n_1414)
);

INVx3_ASAP7_75t_L g1415 ( 
.A(n_1258),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1302),
.B(n_1327),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1282),
.B(n_1279),
.Y(n_1417)
);

AO21x2_ASAP7_75t_L g1418 ( 
.A1(n_1255),
.A2(n_1301),
.B(n_1360),
.Y(n_1418)
);

AND2x4_ASAP7_75t_SL g1419 ( 
.A(n_1353),
.B(n_1360),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1282),
.B(n_1279),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1350),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1355),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1346),
.B(n_1354),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1356),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1359),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1362),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1258),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1363),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1364),
.Y(n_1429)
);

AO21x2_ASAP7_75t_L g1430 ( 
.A1(n_1366),
.A2(n_1262),
.B(n_1254),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1267),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1326),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1277),
.B(n_1292),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1260),
.Y(n_1434)
);

BUFx4f_ASAP7_75t_SL g1435 ( 
.A(n_1352),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1290),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1316),
.Y(n_1437)
);

AO21x2_ASAP7_75t_L g1438 ( 
.A1(n_1296),
.A2(n_1295),
.B(n_1288),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_1365),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1367),
.B(n_1289),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1289),
.B(n_1324),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1291),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1316),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1344),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1291),
.Y(n_1445)
);

AO21x2_ASAP7_75t_L g1446 ( 
.A1(n_1324),
.A2(n_1308),
.B(n_1297),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1308),
.B(n_1294),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1294),
.Y(n_1448)
);

NOR2x1_ASAP7_75t_L g1449 ( 
.A(n_1257),
.B(n_1368),
.Y(n_1449)
);

INVx2_ASAP7_75t_SL g1450 ( 
.A(n_1337),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1259),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1287),
.B(n_1278),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1303),
.B(n_1311),
.Y(n_1453)
);

NAND3xp33_ASAP7_75t_L g1454 ( 
.A(n_1307),
.B(n_1320),
.C(n_1314),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1336),
.Y(n_1455)
);

INVx1_ASAP7_75t_SL g1456 ( 
.A(n_1337),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1338),
.Y(n_1457)
);

OAI211xp5_ASAP7_75t_L g1458 ( 
.A1(n_1298),
.A2(n_1314),
.B(n_1320),
.C(n_1322),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1311),
.B(n_1303),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1275),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1333),
.B(n_1329),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1430),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1418),
.B(n_1397),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1430),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1430),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1407),
.Y(n_1466)
);

INVx2_ASAP7_75t_SL g1467 ( 
.A(n_1419),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1418),
.Y(n_1468)
);

AOI222xp33_ASAP7_75t_L g1469 ( 
.A1(n_1391),
.A2(n_1264),
.B1(n_1307),
.B2(n_1281),
.C1(n_1283),
.C2(n_1293),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1376),
.B(n_1281),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1407),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1418),
.B(n_1256),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1391),
.A2(n_1286),
.B1(n_1298),
.B2(n_1273),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1387),
.B(n_1271),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1407),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1372),
.B(n_1323),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1390),
.B(n_1273),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1418),
.B(n_1280),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1382),
.B(n_1323),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1382),
.B(n_1323),
.Y(n_1480)
);

INVxp67_ASAP7_75t_L g1481 ( 
.A(n_1451),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1412),
.B(n_1414),
.Y(n_1482)
);

INVx4_ASAP7_75t_L g1483 ( 
.A(n_1406),
.Y(n_1483)
);

INVx3_ASAP7_75t_L g1484 ( 
.A(n_1374),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1380),
.B(n_1280),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1414),
.B(n_1247),
.Y(n_1486)
);

AOI222xp33_ASAP7_75t_L g1487 ( 
.A1(n_1381),
.A2(n_1247),
.B1(n_1244),
.B2(n_1265),
.C1(n_1332),
.C2(n_1334),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1421),
.B(n_1309),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1396),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1421),
.B(n_1300),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1400),
.B(n_1330),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1375),
.B(n_1299),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1373),
.A2(n_1284),
.B1(n_1265),
.B2(n_1299),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1400),
.B(n_1299),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1433),
.B(n_1299),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1435),
.B(n_1245),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1375),
.B(n_1312),
.Y(n_1497)
);

AOI221xp5_ASAP7_75t_L g1498 ( 
.A1(n_1381),
.A2(n_1343),
.B1(n_1361),
.B2(n_1401),
.C(n_1402),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1422),
.B(n_1426),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1426),
.B(n_1428),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1428),
.B(n_1394),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1383),
.B(n_1384),
.Y(n_1502)
);

OAI33xp33_ASAP7_75t_L g1503 ( 
.A1(n_1388),
.A2(n_1411),
.A3(n_1429),
.B1(n_1425),
.B2(n_1405),
.B3(n_1424),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1394),
.B(n_1395),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1395),
.B(n_1386),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1405),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1444),
.B(n_1385),
.Y(n_1507)
);

NOR2x1_ASAP7_75t_L g1508 ( 
.A(n_1449),
.B(n_1398),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1385),
.B(n_1402),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1408),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1410),
.B(n_1434),
.Y(n_1511)
);

INVxp67_ASAP7_75t_L g1512 ( 
.A(n_1439),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1396),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1386),
.B(n_1417),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1417),
.B(n_1420),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1410),
.B(n_1393),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1498),
.A2(n_1373),
.B1(n_1401),
.B2(n_1446),
.Y(n_1517)
);

OAI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1473),
.A2(n_1399),
.B1(n_1413),
.B2(n_1454),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1466),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1506),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1505),
.B(n_1416),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1505),
.B(n_1416),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1506),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1501),
.B(n_1374),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_SL g1525 ( 
.A1(n_1515),
.A2(n_1447),
.B1(n_1446),
.B2(n_1441),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1489),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1493),
.A2(n_1399),
.B1(n_1454),
.B2(n_1447),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1507),
.B(n_1393),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1515),
.B(n_1404),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_SL g1530 ( 
.A(n_1469),
.B(n_1379),
.Y(n_1530)
);

OAI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1469),
.A2(n_1508),
.B(n_1478),
.Y(n_1531)
);

NAND3xp33_ASAP7_75t_L g1532 ( 
.A(n_1487),
.B(n_1398),
.C(n_1441),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1510),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1509),
.B(n_1432),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_1496),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1516),
.B(n_1420),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1504),
.B(n_1446),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_1470),
.B(n_1379),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1463),
.B(n_1383),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1511),
.A2(n_1398),
.B1(n_1389),
.B2(n_1379),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1477),
.B(n_1458),
.Y(n_1541)
);

NAND3xp33_ASAP7_75t_L g1542 ( 
.A(n_1481),
.B(n_1398),
.C(n_1448),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1514),
.B(n_1512),
.Y(n_1543)
);

OAI21xp33_ASAP7_75t_L g1544 ( 
.A1(n_1495),
.A2(n_1398),
.B(n_1440),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1482),
.B(n_1446),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1482),
.B(n_1389),
.Y(n_1546)
);

NAND4xp25_ASAP7_75t_SL g1547 ( 
.A(n_1508),
.B(n_1440),
.C(n_1455),
.D(n_1456),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1476),
.B(n_1378),
.Y(n_1548)
);

OAI221xp5_ASAP7_75t_SL g1549 ( 
.A1(n_1478),
.A2(n_1389),
.B1(n_1448),
.B2(n_1442),
.C(n_1445),
.Y(n_1549)
);

OAI221xp5_ASAP7_75t_SL g1550 ( 
.A1(n_1474),
.A2(n_1389),
.B1(n_1445),
.B2(n_1442),
.C(n_1439),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1476),
.B(n_1409),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1486),
.B(n_1409),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1499),
.B(n_1389),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1486),
.B(n_1411),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1488),
.A2(n_1438),
.B1(n_1377),
.B2(n_1369),
.Y(n_1555)
);

NAND4xp25_ASAP7_75t_L g1556 ( 
.A(n_1491),
.B(n_1452),
.C(n_1423),
.D(n_1443),
.Y(n_1556)
);

OA21x2_ASAP7_75t_L g1557 ( 
.A1(n_1462),
.A2(n_1384),
.B(n_1392),
.Y(n_1557)
);

OAI21xp5_ASAP7_75t_SL g1558 ( 
.A1(n_1497),
.A2(n_1369),
.B(n_1455),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1513),
.B(n_1424),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1499),
.B(n_1369),
.Y(n_1560)
);

AOI221xp5_ASAP7_75t_L g1561 ( 
.A1(n_1503),
.A2(n_1423),
.B1(n_1425),
.B2(n_1429),
.C(n_1436),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1488),
.A2(n_1379),
.B1(n_1377),
.B2(n_1443),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1500),
.B(n_1375),
.Y(n_1563)
);

NOR3xp33_ASAP7_75t_L g1564 ( 
.A(n_1485),
.B(n_1456),
.C(n_1427),
.Y(n_1564)
);

NAND4xp25_ASAP7_75t_SL g1565 ( 
.A(n_1490),
.B(n_1459),
.C(n_1449),
.D(n_1461),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_L g1566 ( 
.A(n_1494),
.B(n_1437),
.Y(n_1566)
);

AOI211xp5_ASAP7_75t_SL g1567 ( 
.A1(n_1472),
.A2(n_1415),
.B(n_1427),
.C(n_1406),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1484),
.B(n_1479),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_L g1569 ( 
.A(n_1490),
.B(n_1437),
.Y(n_1569)
);

OAI221xp5_ASAP7_75t_SL g1570 ( 
.A1(n_1485),
.A2(n_1377),
.B1(n_1437),
.B2(n_1443),
.C(n_1457),
.Y(n_1570)
);

NAND3xp33_ASAP7_75t_L g1571 ( 
.A(n_1472),
.B(n_1431),
.C(n_1436),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_SL g1572 ( 
.A(n_1497),
.B(n_1370),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1557),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1520),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1539),
.B(n_1463),
.Y(n_1575)
);

NAND2x1p5_ASAP7_75t_L g1576 ( 
.A(n_1530),
.B(n_1483),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1520),
.Y(n_1577)
);

BUFx2_ASAP7_75t_SL g1578 ( 
.A(n_1526),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1568),
.B(n_1468),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1528),
.B(n_1462),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1523),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1539),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1537),
.B(n_1468),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1521),
.B(n_1484),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1523),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1537),
.B(n_1502),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1521),
.B(n_1479),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1533),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1522),
.B(n_1480),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1533),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1545),
.B(n_1464),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1545),
.B(n_1464),
.Y(n_1592)
);

AND2x4_ASAP7_75t_SL g1593 ( 
.A(n_1564),
.B(n_1497),
.Y(n_1593)
);

INVx2_ASAP7_75t_SL g1594 ( 
.A(n_1519),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1536),
.B(n_1465),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1557),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1571),
.B(n_1559),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1571),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1557),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1522),
.B(n_1480),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1546),
.B(n_1466),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1553),
.B(n_1471),
.Y(n_1602)
);

NOR2x1_ASAP7_75t_R g1603 ( 
.A(n_1535),
.B(n_1371),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1553),
.B(n_1471),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1524),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1534),
.B(n_1465),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1560),
.B(n_1475),
.Y(n_1607)
);

AND2x4_ASAP7_75t_L g1608 ( 
.A(n_1563),
.B(n_1483),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_L g1609 ( 
.A(n_1535),
.B(n_1461),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1574),
.Y(n_1610)
);

INVxp67_ASAP7_75t_L g1611 ( 
.A(n_1597),
.Y(n_1611)
);

INVxp67_ASAP7_75t_SL g1612 ( 
.A(n_1598),
.Y(n_1612)
);

A2O1A1Ixp33_ASAP7_75t_L g1613 ( 
.A1(n_1593),
.A2(n_1532),
.B(n_1544),
.C(n_1525),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1597),
.B(n_1551),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1595),
.B(n_1529),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1574),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1603),
.B(n_1541),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1582),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1579),
.B(n_1531),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1577),
.Y(n_1620)
);

AND2x4_ASAP7_75t_SL g1621 ( 
.A(n_1608),
.B(n_1497),
.Y(n_1621)
);

BUFx2_ASAP7_75t_L g1622 ( 
.A(n_1576),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1603),
.B(n_1569),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1591),
.B(n_1552),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1595),
.B(n_1554),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1577),
.Y(n_1626)
);

INVx1_ASAP7_75t_SL g1627 ( 
.A(n_1578),
.Y(n_1627)
);

INVxp67_ASAP7_75t_L g1628 ( 
.A(n_1578),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1581),
.Y(n_1629)
);

NOR2xp67_ASAP7_75t_SL g1630 ( 
.A(n_1598),
.B(n_1532),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1593),
.B(n_1567),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1573),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1581),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1585),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1585),
.Y(n_1635)
);

AND2x4_ASAP7_75t_SL g1636 ( 
.A(n_1608),
.B(n_1492),
.Y(n_1636)
);

BUFx2_ASAP7_75t_L g1637 ( 
.A(n_1576),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1580),
.B(n_1544),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1588),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1593),
.B(n_1563),
.Y(n_1640)
);

NAND2x1p5_ASAP7_75t_L g1641 ( 
.A(n_1594),
.B(n_1467),
.Y(n_1641)
);

AOI32xp33_ASAP7_75t_L g1642 ( 
.A1(n_1587),
.A2(n_1517),
.A3(n_1527),
.B1(n_1518),
.B2(n_1540),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1580),
.B(n_1587),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1584),
.B(n_1543),
.Y(n_1644)
);

BUFx2_ASAP7_75t_L g1645 ( 
.A(n_1576),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1588),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1590),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1573),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1584),
.B(n_1558),
.Y(n_1649)
);

AOI32xp33_ASAP7_75t_L g1650 ( 
.A1(n_1589),
.A2(n_1555),
.A3(n_1562),
.B1(n_1566),
.B2(n_1548),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1591),
.B(n_1542),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1611),
.B(n_1589),
.Y(n_1652)
);

NOR2xp33_ASAP7_75t_SL g1653 ( 
.A(n_1630),
.B(n_1570),
.Y(n_1653)
);

INVx1_ASAP7_75t_SL g1654 ( 
.A(n_1627),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1631),
.B(n_1608),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1632),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1610),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1614),
.B(n_1600),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1610),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1634),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1632),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1634),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1651),
.B(n_1592),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1631),
.B(n_1608),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1621),
.B(n_1600),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1651),
.B(n_1592),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1621),
.B(n_1601),
.Y(n_1667)
);

INVx2_ASAP7_75t_SL g1668 ( 
.A(n_1636),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1636),
.B(n_1601),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1619),
.B(n_1602),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1618),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1612),
.B(n_1643),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1648),
.Y(n_1673)
);

AND3x2_ASAP7_75t_L g1674 ( 
.A(n_1617),
.B(n_1609),
.C(n_1605),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1638),
.B(n_1602),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1616),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1630),
.A2(n_1565),
.B1(n_1547),
.B2(n_1556),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1619),
.B(n_1649),
.Y(n_1678)
);

INVxp67_ASAP7_75t_L g1679 ( 
.A(n_1623),
.Y(n_1679)
);

INVx1_ASAP7_75t_SL g1680 ( 
.A(n_1622),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1649),
.B(n_1622),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1628),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1620),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1650),
.B(n_1604),
.Y(n_1684)
);

OAI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1613),
.A2(n_1542),
.B(n_1556),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1626),
.Y(n_1686)
);

AOI211xp5_ASAP7_75t_L g1687 ( 
.A1(n_1613),
.A2(n_1550),
.B(n_1549),
.C(n_1538),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1648),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1637),
.B(n_1604),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1624),
.B(n_1583),
.Y(n_1690)
);

NAND2xp33_ASAP7_75t_SL g1691 ( 
.A(n_1640),
.B(n_1572),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1629),
.Y(n_1692)
);

OAI32xp33_ASAP7_75t_L g1693 ( 
.A1(n_1641),
.A2(n_1583),
.A3(n_1606),
.B1(n_1586),
.B2(n_1599),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1615),
.B(n_1606),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1624),
.B(n_1575),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1633),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1625),
.B(n_1607),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1656),
.Y(n_1698)
);

BUFx3_ASAP7_75t_L g1699 ( 
.A(n_1654),
.Y(n_1699)
);

INVx1_ASAP7_75t_SL g1700 ( 
.A(n_1680),
.Y(n_1700)
);

CKINVDCx20_ASAP7_75t_R g1701 ( 
.A(n_1679),
.Y(n_1701)
);

INVx1_ASAP7_75t_SL g1702 ( 
.A(n_1680),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1656),
.Y(n_1703)
);

HB1xp67_ASAP7_75t_L g1704 ( 
.A(n_1671),
.Y(n_1704)
);

INVx1_ASAP7_75t_SL g1705 ( 
.A(n_1674),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1657),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1682),
.B(n_1635),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1656),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1653),
.B(n_1684),
.Y(n_1709)
);

BUFx3_ASAP7_75t_L g1710 ( 
.A(n_1681),
.Y(n_1710)
);

INVx1_ASAP7_75t_SL g1711 ( 
.A(n_1681),
.Y(n_1711)
);

INVx1_ASAP7_75t_SL g1712 ( 
.A(n_1678),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_1678),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1672),
.B(n_1639),
.Y(n_1714)
);

INVxp67_ASAP7_75t_L g1715 ( 
.A(n_1653),
.Y(n_1715)
);

OAI21xp33_ASAP7_75t_SL g1716 ( 
.A1(n_1685),
.A2(n_1642),
.B(n_1640),
.Y(n_1716)
);

OA21x2_ASAP7_75t_L g1717 ( 
.A1(n_1661),
.A2(n_1596),
.B(n_1573),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1672),
.B(n_1646),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1655),
.B(n_1637),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1657),
.Y(n_1720)
);

CKINVDCx16_ASAP7_75t_R g1721 ( 
.A(n_1691),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1668),
.B(n_1655),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1664),
.B(n_1670),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1659),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1659),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1660),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1660),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1661),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1662),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1694),
.B(n_1647),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1661),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1664),
.B(n_1670),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1662),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1668),
.B(n_1645),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1676),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1676),
.Y(n_1736)
);

NOR4xp25_ASAP7_75t_L g1737 ( 
.A(n_1716),
.B(n_1677),
.C(n_1663),
.D(n_1666),
.Y(n_1737)
);

INVx1_ASAP7_75t_SL g1738 ( 
.A(n_1699),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1710),
.Y(n_1739)
);

OAI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1721),
.A2(n_1687),
.B1(n_1652),
.B2(n_1675),
.Y(n_1740)
);

INVxp67_ASAP7_75t_SL g1741 ( 
.A(n_1699),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1723),
.B(n_1665),
.Y(n_1742)
);

AOI222xp33_ASAP7_75t_L g1743 ( 
.A1(n_1716),
.A2(n_1693),
.B1(n_1645),
.B2(n_1687),
.C1(n_1689),
.C2(n_1658),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1713),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1723),
.B(n_1665),
.Y(n_1745)
);

OAI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1721),
.A2(n_1667),
.B1(n_1669),
.B2(n_1697),
.Y(n_1746)
);

OAI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1705),
.A2(n_1667),
.B1(n_1669),
.B2(n_1666),
.Y(n_1747)
);

INVx1_ASAP7_75t_SL g1748 ( 
.A(n_1699),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_SL g1749 ( 
.A(n_1701),
.B(n_1693),
.Y(n_1749)
);

O2A1O1Ixp33_ASAP7_75t_L g1750 ( 
.A1(n_1715),
.A2(n_1663),
.B(n_1696),
.C(n_1692),
.Y(n_1750)
);

O2A1O1Ixp5_ASAP7_75t_L g1751 ( 
.A1(n_1709),
.A2(n_1696),
.B(n_1683),
.C(n_1692),
.Y(n_1751)
);

NOR2xp67_ASAP7_75t_L g1752 ( 
.A(n_1704),
.B(n_1683),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1706),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1711),
.B(n_1689),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1711),
.B(n_1686),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1705),
.B(n_1695),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_1700),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1706),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1710),
.B(n_1686),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1710),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1732),
.B(n_1719),
.Y(n_1761)
);

AOI21xp5_ASAP7_75t_L g1762 ( 
.A1(n_1712),
.A2(n_1690),
.B(n_1695),
.Y(n_1762)
);

BUFx2_ASAP7_75t_L g1763 ( 
.A(n_1722),
.Y(n_1763)
);

INVx1_ASAP7_75t_SL g1764 ( 
.A(n_1712),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1720),
.Y(n_1765)
);

BUFx3_ASAP7_75t_L g1766 ( 
.A(n_1757),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1741),
.B(n_1700),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_SL g1768 ( 
.A(n_1737),
.B(n_1702),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1763),
.Y(n_1769)
);

AOI221x1_ASAP7_75t_SL g1770 ( 
.A1(n_1740),
.A2(n_1707),
.B1(n_1722),
.B2(n_1736),
.C(n_1735),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_L g1771 ( 
.A(n_1738),
.B(n_1702),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1763),
.Y(n_1772)
);

NAND3xp33_ASAP7_75t_L g1773 ( 
.A(n_1743),
.B(n_1707),
.C(n_1734),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1748),
.B(n_1730),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1744),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1757),
.B(n_1722),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1764),
.B(n_1754),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1744),
.Y(n_1778)
);

INVx1_ASAP7_75t_SL g1779 ( 
.A(n_1761),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1756),
.B(n_1732),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1761),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1739),
.B(n_1722),
.Y(n_1782)
);

AND2x4_ASAP7_75t_L g1783 ( 
.A(n_1752),
.B(n_1719),
.Y(n_1783)
);

HB1xp67_ASAP7_75t_L g1784 ( 
.A(n_1752),
.Y(n_1784)
);

OAI221xp5_ASAP7_75t_L g1785 ( 
.A1(n_1749),
.A2(n_1718),
.B1(n_1714),
.B2(n_1734),
.C(n_1730),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1742),
.B(n_1714),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1742),
.B(n_1718),
.Y(n_1787)
);

AOI21xp33_ASAP7_75t_SL g1788 ( 
.A1(n_1747),
.A2(n_1736),
.B(n_1735),
.Y(n_1788)
);

NAND4xp25_ASAP7_75t_L g1789 ( 
.A(n_1770),
.B(n_1776),
.C(n_1768),
.D(n_1766),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1768),
.A2(n_1746),
.B1(n_1739),
.B2(n_1760),
.Y(n_1790)
);

OAI211xp5_ASAP7_75t_L g1791 ( 
.A1(n_1773),
.A2(n_1750),
.B(n_1760),
.C(n_1759),
.Y(n_1791)
);

AOI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1785),
.A2(n_1751),
.B(n_1755),
.Y(n_1792)
);

OAI221xp5_ASAP7_75t_L g1793 ( 
.A1(n_1780),
.A2(n_1762),
.B1(n_1745),
.B2(n_1758),
.C(n_1753),
.Y(n_1793)
);

OAI21xp33_ASAP7_75t_L g1794 ( 
.A1(n_1776),
.A2(n_1745),
.B(n_1753),
.Y(n_1794)
);

AOI21xp5_ASAP7_75t_L g1795 ( 
.A1(n_1784),
.A2(n_1765),
.B(n_1758),
.Y(n_1795)
);

NOR2x1_ASAP7_75t_L g1796 ( 
.A(n_1766),
.B(n_1765),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1771),
.B(n_1720),
.Y(n_1797)
);

AOI21xp33_ASAP7_75t_SL g1798 ( 
.A1(n_1771),
.A2(n_1725),
.B(n_1724),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1769),
.Y(n_1799)
);

AOI221xp5_ASAP7_75t_L g1800 ( 
.A1(n_1788),
.A2(n_1733),
.B1(n_1724),
.B2(n_1729),
.C(n_1725),
.Y(n_1800)
);

OAI221xp5_ASAP7_75t_L g1801 ( 
.A1(n_1767),
.A2(n_1733),
.B1(n_1726),
.B2(n_1729),
.C(n_1727),
.Y(n_1801)
);

NAND3xp33_ASAP7_75t_L g1802 ( 
.A(n_1777),
.B(n_1727),
.C(n_1726),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1790),
.B(n_1783),
.Y(n_1803)
);

OAI22xp5_ASAP7_75t_SL g1804 ( 
.A1(n_1797),
.A2(n_1772),
.B1(n_1779),
.B2(n_1778),
.Y(n_1804)
);

OAI211xp5_ASAP7_75t_SL g1805 ( 
.A1(n_1791),
.A2(n_1782),
.B(n_1774),
.C(n_1775),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1792),
.A2(n_1783),
.B(n_1781),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1796),
.Y(n_1807)
);

NOR3xp33_ASAP7_75t_L g1808 ( 
.A(n_1789),
.B(n_1781),
.C(n_1787),
.Y(n_1808)
);

AOI211xp5_ASAP7_75t_L g1809 ( 
.A1(n_1798),
.A2(n_1783),
.B(n_1787),
.C(n_1786),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1799),
.Y(n_1810)
);

NAND3xp33_ASAP7_75t_SL g1811 ( 
.A(n_1794),
.B(n_1786),
.C(n_1703),
.Y(n_1811)
);

OA22x2_ASAP7_75t_L g1812 ( 
.A1(n_1793),
.A2(n_1731),
.B1(n_1728),
.B2(n_1708),
.Y(n_1812)
);

AOI21xp5_ASAP7_75t_L g1813 ( 
.A1(n_1795),
.A2(n_1703),
.B(n_1698),
.Y(n_1813)
);

NOR3xp33_ASAP7_75t_SL g1814 ( 
.A(n_1801),
.B(n_1403),
.C(n_1371),
.Y(n_1814)
);

NOR2x1_ASAP7_75t_L g1815 ( 
.A(n_1802),
.B(n_1698),
.Y(n_1815)
);

NAND3xp33_ASAP7_75t_L g1816 ( 
.A(n_1808),
.B(n_1800),
.C(n_1703),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1806),
.B(n_1690),
.Y(n_1817)
);

OAI221xp5_ASAP7_75t_L g1818 ( 
.A1(n_1805),
.A2(n_1731),
.B1(n_1728),
.B2(n_1708),
.C(n_1698),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1815),
.Y(n_1819)
);

NAND5xp2_ASAP7_75t_L g1820 ( 
.A(n_1809),
.B(n_1641),
.C(n_1561),
.D(n_1453),
.E(n_1403),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1807),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1811),
.Y(n_1822)
);

AOI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1822),
.A2(n_1803),
.B1(n_1804),
.B2(n_1814),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1819),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1817),
.B(n_1810),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1821),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1816),
.Y(n_1827)
);

INVxp67_ASAP7_75t_L g1828 ( 
.A(n_1818),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_SL g1829 ( 
.A(n_1820),
.B(n_1812),
.Y(n_1829)
);

O2A1O1Ixp33_ASAP7_75t_L g1830 ( 
.A1(n_1827),
.A2(n_1828),
.B(n_1824),
.C(n_1825),
.Y(n_1830)
);

NAND4xp25_ASAP7_75t_L g1831 ( 
.A(n_1823),
.B(n_1813),
.C(n_1708),
.D(n_1731),
.Y(n_1831)
);

OR5x1_ASAP7_75t_L g1832 ( 
.A(n_1829),
.B(n_1826),
.C(n_1728),
.D(n_1717),
.E(n_1688),
.Y(n_1832)
);

INVxp33_ASAP7_75t_SL g1833 ( 
.A(n_1823),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1824),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1827),
.B(n_1673),
.Y(n_1835)
);

NAND5xp2_ASAP7_75t_L g1836 ( 
.A(n_1833),
.B(n_1830),
.C(n_1831),
.D(n_1832),
.E(n_1834),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1835),
.B(n_1673),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1835),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1833),
.B(n_1673),
.Y(n_1839)
);

AO22x2_ASAP7_75t_L g1840 ( 
.A1(n_1838),
.A2(n_1688),
.B1(n_1594),
.B2(n_1599),
.Y(n_1840)
);

NAND4xp75_ASAP7_75t_L g1841 ( 
.A(n_1840),
.B(n_1839),
.C(n_1837),
.D(n_1836),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1841),
.B(n_1688),
.Y(n_1842)
);

NOR2x1_ASAP7_75t_L g1843 ( 
.A(n_1841),
.B(n_1717),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1843),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1842),
.B(n_1717),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1844),
.B(n_1644),
.Y(n_1846)
);

NOR2xp33_ASAP7_75t_L g1847 ( 
.A(n_1845),
.B(n_1371),
.Y(n_1847)
);

XOR2xp5_ASAP7_75t_L g1848 ( 
.A(n_1846),
.B(n_1403),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1848),
.Y(n_1849)
);

OAI221xp5_ASAP7_75t_R g1850 ( 
.A1(n_1849),
.A2(n_1847),
.B1(n_1717),
.B2(n_1641),
.C(n_1594),
.Y(n_1850)
);

AOI211xp5_ASAP7_75t_L g1851 ( 
.A1(n_1850),
.A2(n_1370),
.B(n_1450),
.C(n_1460),
.Y(n_1851)
);


endmodule