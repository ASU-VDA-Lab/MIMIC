module fake_jpeg_4998_n_337 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_48),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_15),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_45),
.Y(n_68)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_49),
.Y(n_85)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_51),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_27),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_53),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_26),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_54),
.Y(n_79)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_14),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_26),
.B(n_1),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_56),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_16),
.Y(n_56)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_45),
.A2(n_23),
.B1(n_32),
.B2(n_18),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_59),
.A2(n_60),
.B(n_61),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_23),
.B1(n_32),
.B2(n_18),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_46),
.A2(n_16),
.B1(n_25),
.B2(n_33),
.Y(n_61)
);

NAND2x1_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_28),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_10),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_25),
.B1(n_33),
.B2(n_22),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_42),
.A2(n_34),
.B1(n_31),
.B2(n_24),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_70),
.A2(n_73),
.B1(n_74),
.B2(n_80),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_42),
.A2(n_53),
.B1(n_50),
.B2(n_39),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_50),
.A2(n_34),
.B1(n_31),
.B2(n_24),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_49),
.A2(n_22),
.B1(n_21),
.B2(n_28),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_75),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_49),
.A2(n_28),
.B1(n_21),
.B2(n_30),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_77),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_28),
.B1(n_21),
.B2(n_30),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_78),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_43),
.A2(n_21),
.B1(n_31),
.B2(n_24),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_53),
.A2(n_34),
.B1(n_20),
.B2(n_3),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_89),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_43),
.A2(n_20),
.B1(n_2),
.B2(n_3),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_54),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_11),
.Y(n_117)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_88),
.Y(n_108)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_56),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_99),
.Y(n_126)
);

CKINVDCx6p67_ASAP7_75t_R g92 ( 
.A(n_38),
.Y(n_92)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_92),
.Y(n_138)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_47),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_94),
.B1(n_97),
.B2(n_11),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_37),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_37),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_93),
.B1(n_100),
.B2(n_98),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_51),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g123 ( 
.A(n_98),
.Y(n_123)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_39),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_39),
.Y(n_102)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_103),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_63),
.B(n_7),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_106),
.B(n_110),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_65),
.B(n_93),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_107),
.B(n_112),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_63),
.B(n_9),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_64),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_111),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_117),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_65),
.A2(n_11),
.B1(n_93),
.B2(n_91),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_118),
.A2(n_96),
.B1(n_101),
.B2(n_104),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_76),
.B(n_11),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_124),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_121),
.A2(n_67),
.B1(n_58),
.B2(n_84),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_63),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_64),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_105),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_139),
.B(n_155),
.Y(n_196)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_136),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_145),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_111),
.B(n_79),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_166),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_107),
.A2(n_68),
.B(n_102),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_142),
.A2(n_173),
.B(n_112),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_128),
.A2(n_99),
.B1(n_66),
.B2(n_86),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_143),
.A2(n_148),
.B(n_150),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_107),
.A2(n_97),
.B(n_79),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_154),
.Y(n_185)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_67),
.B1(n_90),
.B2(n_70),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_146),
.A2(n_162),
.B1(n_163),
.B2(n_122),
.Y(n_195)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_149),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_107),
.A2(n_66),
.B1(n_71),
.B2(n_87),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_71),
.Y(n_150)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_151),
.B(n_160),
.Y(n_193)
);

AND2x6_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_92),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_88),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_156),
.B(n_158),
.Y(n_198)
);

OAI21xp33_ASAP7_75t_SL g183 ( 
.A1(n_157),
.A2(n_165),
.B(n_125),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_119),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_108),
.Y(n_160)
);

AND2x6_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_92),
.Y(n_161)
);

A2O1A1O1Ixp25_ASAP7_75t_L g210 ( 
.A1(n_161),
.A2(n_133),
.B(n_135),
.C(n_137),
.D(n_116),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_113),
.A2(n_74),
.B1(n_73),
.B2(n_81),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_131),
.A2(n_62),
.B1(n_85),
.B2(n_92),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_164),
.A2(n_174),
.B1(n_134),
.B2(n_106),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_127),
.A2(n_72),
.B1(n_96),
.B2(n_57),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_57),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_168),
.B(n_170),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_120),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_169),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_126),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_112),
.B(n_115),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_144),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_127),
.B(n_132),
.C(n_130),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_118),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_135),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_177),
.B(n_152),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_156),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_178),
.Y(n_217)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_180),
.Y(n_220)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_183),
.A2(n_184),
.B1(n_160),
.B2(n_149),
.Y(n_230)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_186),
.B(n_190),
.Y(n_216)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_110),
.A3(n_134),
.B1(n_117),
.B2(n_125),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_173),
.Y(n_228)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_192),
.B(n_199),
.Y(n_233)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_151),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_195),
.A2(n_212),
.B1(n_167),
.B2(n_153),
.Y(n_223)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_197),
.Y(n_215)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_141),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_176),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_202),
.B(n_205),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_147),
.B(n_122),
.Y(n_203)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_203),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_174),
.A2(n_137),
.B1(n_109),
.B2(n_125),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_204),
.A2(n_176),
.B1(n_175),
.B2(n_172),
.Y(n_235)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_206),
.B(n_172),
.Y(n_241)
);

INVxp33_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_150),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_159),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_213),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_153),
.A2(n_109),
.B1(n_133),
.B2(n_135),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_171),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_163),
.Y(n_214)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_214),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_142),
.C(n_166),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_229),
.C(n_206),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_223),
.A2(n_231),
.B1(n_180),
.B2(n_184),
.Y(n_252)
);

NAND2xp33_ASAP7_75t_SL g226 ( 
.A(n_196),
.B(n_167),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_226),
.A2(n_186),
.B1(n_213),
.B2(n_199),
.Y(n_247)
);

OAI32xp33_ASAP7_75t_L g227 ( 
.A1(n_182),
.A2(n_167),
.A3(n_148),
.B1(n_150),
.B2(n_143),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_227),
.B(n_228),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_192),
.A2(n_201),
.B1(n_209),
.B2(n_181),
.Y(n_231)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_235),
.Y(n_244)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

INVx13_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_152),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_211),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_243),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_195),
.A2(n_116),
.B1(n_147),
.B2(n_145),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_242),
.A2(n_204),
.B1(n_178),
.B2(n_193),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_179),
.B(n_140),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_185),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_245),
.B(n_249),
.C(n_250),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_263),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_247),
.A2(n_257),
.B(n_233),
.Y(n_275)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_237),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_248),
.B(n_255),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_185),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_252),
.A2(n_262),
.B1(n_212),
.B2(n_240),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_202),
.Y(n_253)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_254),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_222),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_236),
.B(n_190),
.Y(n_256)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_238),
.A2(n_177),
.B(n_198),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_234),
.B(n_191),
.Y(n_259)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_259),
.Y(n_285)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_216),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_201),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_243),
.Y(n_268)
);

INVx13_ASAP7_75t_L g265 ( 
.A(n_218),
.Y(n_265)
);

OA22x2_ASAP7_75t_L g271 ( 
.A1(n_265),
.A2(n_200),
.B1(n_188),
.B2(n_225),
.Y(n_271)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_235),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_266),
.A2(n_267),
.B1(n_223),
.B2(n_217),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_242),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_SL g288 ( 
.A(n_268),
.B(n_271),
.C(n_275),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_251),
.A2(n_220),
.B1(n_221),
.B2(n_232),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_269),
.A2(n_278),
.B1(n_281),
.B2(n_283),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_227),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_277),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_229),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_251),
.A2(n_221),
.B1(n_232),
.B2(n_224),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_279),
.A2(n_266),
.B(n_280),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_244),
.A2(n_238),
.B1(n_224),
.B2(n_210),
.Y(n_280)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_280),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_244),
.A2(n_239),
.B1(n_189),
.B2(n_218),
.Y(n_283)
);

BUFx12_ASAP7_75t_L g286 ( 
.A(n_271),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_298),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_284),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_291),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_271),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_258),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_268),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_293),
.A2(n_269),
.B1(n_278),
.B2(n_272),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_245),
.C(n_249),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_296),
.C(n_299),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_250),
.C(n_257),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_253),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_297),
.B(n_265),
.Y(n_309)
);

NOR3xp33_ASAP7_75t_SL g298 ( 
.A(n_275),
.B(n_258),
.C(n_247),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_246),
.Y(n_299)
);

FAx1_ASAP7_75t_SL g317 ( 
.A(n_301),
.B(n_294),
.CI(n_298),
.CON(n_317),
.SN(n_317)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_303),
.C(n_306),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_270),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_290),
.A2(n_255),
.B1(n_262),
.B2(n_274),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_308),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_264),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_294),
.A2(n_279),
.B1(n_248),
.B2(n_263),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_311),
.C(n_299),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_271),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_295),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_293),
.A2(n_285),
.B1(n_273),
.B2(n_215),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_307),
.B(n_260),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_314),
.Y(n_325)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_315),
.Y(n_323)
);

AND2x6_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_288),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_316),
.A2(n_300),
.B1(n_307),
.B2(n_306),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_317),
.B(n_286),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_304),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_318),
.A2(n_319),
.B1(n_286),
.B2(n_194),
.Y(n_327)
);

MAJx2_ASAP7_75t_L g319 ( 
.A(n_303),
.B(n_288),
.C(n_296),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_320),
.B(n_302),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_305),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_321),
.A2(n_316),
.B(n_318),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_324),
.C(n_317),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_326),
.B(n_327),
.Y(n_328)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_329),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_323),
.A2(n_313),
.B(n_319),
.Y(n_330)
);

AOI322xp5_ASAP7_75t_L g332 ( 
.A1(n_330),
.A2(n_331),
.A3(n_323),
.B1(n_324),
.B2(n_325),
.C1(n_321),
.C2(n_254),
.Y(n_332)
);

AO21x1_ASAP7_75t_L g334 ( 
.A1(n_332),
.A2(n_328),
.B(n_260),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_334),
.B(n_333),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_208),
.Y(n_337)
);


endmodule