module fake_jpeg_2506_n_503 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_503);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_503;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx4f_ASAP7_75t_SL g45 ( 
.A(n_1),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_10),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_57),
.Y(n_143)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_59),
.B(n_61),
.Y(n_122)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_60),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_26),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_62),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_18),
.B(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_63),
.B(n_65),
.Y(n_135)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_64),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_18),
.B(n_17),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_26),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_66),
.B(n_68),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_17),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_69),
.B(n_70),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_13),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_71),
.B(n_81),
.Y(n_147)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_73),
.Y(n_193)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_74),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_75),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_78),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_80),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_41),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_83),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_27),
.B(n_12),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_84),
.B(n_86),
.Y(n_168)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_85),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_27),
.B(n_13),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

INVx6_ASAP7_75t_SL g88 ( 
.A(n_45),
.Y(n_88)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_89),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_42),
.B(n_12),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_90),
.B(n_98),
.Y(n_172)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_91),
.Y(n_179)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_92),
.Y(n_184)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_94),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_38),
.B(n_9),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_95),
.B(n_96),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_9),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_97),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_50),
.B(n_0),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_99),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_32),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_100),
.Y(n_148)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_24),
.Y(n_101)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_2),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_102),
.B(n_105),
.Y(n_192)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_25),
.B(n_2),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_28),
.B(n_2),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_106),
.B(n_111),
.Y(n_199)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_107),
.Y(n_173)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_28),
.Y(n_108)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_32),
.Y(n_110)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_110),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_23),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_32),
.Y(n_112)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_112),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_23),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_113),
.B(n_114),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_43),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_23),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_115),
.B(n_117),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_39),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_46),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_43),
.Y(n_120)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_49),
.Y(n_121)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_121),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_88),
.A2(n_56),
.B1(n_46),
.B2(n_30),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g202 ( 
.A1(n_127),
.A2(n_140),
.B1(n_194),
.B2(n_195),
.Y(n_202)
);

BUFx10_ASAP7_75t_L g134 ( 
.A(n_64),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g212 ( 
.A(n_134),
.Y(n_212)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_67),
.Y(n_136)
);

INVx3_ASAP7_75t_SL g227 ( 
.A(n_136),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_90),
.A2(n_51),
.B1(n_30),
.B2(n_19),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_75),
.A2(n_51),
.B1(n_30),
.B2(n_19),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_144),
.A2(n_150),
.B1(n_160),
.B2(n_57),
.Y(n_211)
);

AO22x1_ASAP7_75t_SL g145 ( 
.A1(n_102),
.A2(n_51),
.B1(n_19),
.B2(n_49),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_145),
.B(n_110),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_77),
.A2(n_21),
.B1(n_47),
.B2(n_40),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_101),
.A2(n_52),
.B1(n_21),
.B2(n_29),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_154),
.A2(n_144),
.B1(n_150),
.B2(n_167),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_79),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_156),
.B(n_161),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_103),
.A2(n_29),
.B1(n_47),
.B2(n_40),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_114),
.B(n_52),
.Y(n_161)
);

AOI21xp33_ASAP7_75t_L g163 ( 
.A1(n_120),
.A2(n_36),
.B(n_35),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_163),
.B(n_180),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_104),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_174),
.Y(n_232)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_64),
.Y(n_175)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_175),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_116),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_176),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_119),
.B(n_39),
.Y(n_180)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_89),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_183),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_121),
.B(n_36),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_185),
.B(n_197),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_58),
.B(n_39),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_186),
.B(n_187),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_78),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_82),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_190),
.B(n_196),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_100),
.A2(n_35),
.B1(n_33),
.B2(n_4),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_92),
.A2(n_33),
.B1(n_3),
.B2(n_4),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_97),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_73),
.B(n_2),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_109),
.Y(n_198)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_198),
.Y(n_241)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_74),
.Y(n_200)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_200),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_201),
.A2(n_85),
.B(n_118),
.Y(n_203)
);

OA21x2_ASAP7_75t_L g283 ( 
.A1(n_203),
.A2(n_224),
.B(n_225),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_201),
.A2(n_107),
.B1(n_99),
.B2(n_93),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_204),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_146),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_205),
.B(n_206),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_137),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_181),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_207),
.B(n_209),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

INVxp67_ASAP7_75t_SL g289 ( 
.A(n_208),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_5),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_126),
.Y(n_210)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_210),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_211),
.B(n_217),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_6),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_213),
.B(n_221),
.Y(n_281)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_171),
.Y(n_214)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_214),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_154),
.A2(n_60),
.B1(n_62),
.B2(n_33),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_215),
.A2(n_203),
.B1(n_218),
.B2(n_240),
.Y(n_274)
);

OAI32xp33_ASAP7_75t_L g217 ( 
.A1(n_172),
.A2(n_192),
.A3(n_169),
.B1(n_145),
.B2(n_168),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_218),
.A2(n_261),
.B1(n_256),
.B2(n_227),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_166),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_219),
.B(n_220),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_147),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_172),
.B(n_6),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_147),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_222),
.B(n_223),
.Y(n_277)
);

A2O1A1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_135),
.A2(n_112),
.B(n_76),
.C(n_8),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_127),
.A2(n_6),
.B(n_7),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_160),
.A2(n_6),
.B(n_7),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_135),
.A2(n_168),
.B(n_122),
.C(n_180),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_226),
.B(n_213),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_165),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_228),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_191),
.A2(n_7),
.B1(n_9),
.B2(n_139),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_230),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_125),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_231),
.Y(n_291)
);

BUFx12f_ASAP7_75t_L g233 ( 
.A(n_134),
.Y(n_233)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_233),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_152),
.A2(n_186),
.B1(n_148),
.B2(n_177),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_234),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_132),
.A2(n_182),
.B1(n_188),
.B2(n_128),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_236),
.B(n_240),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_189),
.A2(n_159),
.B1(n_178),
.B2(n_184),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_238),
.Y(n_316)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_133),
.Y(n_239)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_239),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_194),
.A2(n_195),
.B(n_140),
.Y(n_246)
);

NAND2x1_ASAP7_75t_SL g302 ( 
.A(n_246),
.B(n_256),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_124),
.B(n_151),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_247),
.B(n_248),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_179),
.B(n_129),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_141),
.Y(n_249)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_249),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_164),
.B(n_159),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_250),
.B(n_253),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_170),
.B(n_173),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_251),
.B(n_260),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_130),
.A2(n_149),
.B1(n_123),
.B2(n_162),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_252),
.A2(n_255),
.B1(n_258),
.B2(n_259),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_178),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_184),
.Y(n_254)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_254),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_131),
.A2(n_162),
.B1(n_182),
.B2(n_166),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_158),
.B(n_143),
.Y(n_256)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_131),
.Y(n_257)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_257),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_157),
.A2(n_142),
.B1(n_155),
.B2(n_138),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_142),
.A2(n_181),
.B1(n_144),
.B2(n_140),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_153),
.B(n_134),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_160),
.A2(n_150),
.B1(n_144),
.B2(n_163),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_175),
.Y(n_262)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_262),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_181),
.B(n_169),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_205),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_131),
.Y(n_265)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_265),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_144),
.A2(n_140),
.B1(n_160),
.B2(n_150),
.Y(n_266)
);

AO21x2_ASAP7_75t_L g299 ( 
.A1(n_266),
.A2(n_225),
.B(n_251),
.Y(n_299)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_171),
.Y(n_267)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_267),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_229),
.B(n_207),
.C(n_222),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_269),
.B(n_212),
.C(n_281),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_274),
.A2(n_296),
.B1(n_301),
.B2(n_202),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_280),
.B(n_290),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_244),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_286),
.B(n_315),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_216),
.B(n_221),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_292),
.B(n_281),
.C(n_269),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_218),
.A2(n_246),
.B1(n_266),
.B2(n_217),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_239),
.Y(n_297)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_297),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_299),
.A2(n_245),
.B1(n_243),
.B2(n_241),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_224),
.A2(n_202),
.B1(n_237),
.B2(n_236),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_202),
.A2(n_256),
.B1(n_260),
.B2(n_223),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_304),
.Y(n_318)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_249),
.Y(n_306)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_306),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_209),
.B(n_242),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_307),
.B(n_313),
.Y(n_337)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_257),
.Y(n_308)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_308),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_309),
.A2(n_212),
.B(n_233),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_202),
.A2(n_254),
.B1(n_210),
.B2(n_243),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_312),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_214),
.B(n_267),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_227),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_231),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_317),
.A2(n_325),
.B1(n_329),
.B2(n_344),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_320),
.A2(n_323),
.B1(n_327),
.B2(n_333),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_299),
.A2(n_206),
.B1(n_245),
.B2(n_226),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_313),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_324),
.B(n_328),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_299),
.A2(n_279),
.B1(n_298),
.B2(n_309),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_294),
.B(n_235),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_326),
.B(n_330),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_299),
.A2(n_232),
.B1(n_265),
.B2(n_235),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_292),
.B(n_262),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_299),
.A2(n_232),
.B1(n_263),
.B2(n_233),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_307),
.B(n_280),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_271),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_331),
.B(n_334),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_332),
.A2(n_342),
.B(n_305),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_279),
.A2(n_212),
.B1(n_233),
.B2(n_263),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_284),
.B(n_212),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_271),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_335),
.B(n_343),
.Y(n_367)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_268),
.Y(n_340)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_340),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_341),
.B(n_293),
.C(n_295),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_302),
.A2(n_277),
.B(n_283),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_282),
.B(n_273),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_279),
.A2(n_296),
.B1(n_274),
.B2(n_301),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_298),
.A2(n_300),
.B1(n_283),
.B2(n_284),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_345),
.A2(n_300),
.B1(n_270),
.B2(n_305),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_285),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_346),
.Y(n_366)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_272),
.Y(n_347)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_347),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_348),
.B(n_341),
.Y(n_355)
);

OAI21xp33_ASAP7_75t_L g349 ( 
.A1(n_283),
.A2(n_276),
.B(n_270),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_349),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_291),
.B(n_287),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_350),
.B(n_314),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_302),
.B(n_288),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_351),
.B(n_289),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_354),
.A2(n_380),
.B1(n_327),
.B2(n_320),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_355),
.B(n_381),
.C(n_341),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_348),
.B(n_278),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_356),
.B(n_362),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_358),
.A2(n_359),
.B(n_365),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_318),
.A2(n_275),
.B(n_316),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_332),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_364),
.B(n_369),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_325),
.A2(n_316),
.B(n_275),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_336),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_368),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_338),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_370),
.B(n_334),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_350),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_371),
.B(n_335),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_342),
.A2(n_291),
.B(n_310),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_373),
.A2(n_379),
.B(n_339),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_338),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_375),
.B(n_343),
.Y(n_392)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_319),
.Y(n_376)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_376),
.Y(n_404)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_336),
.Y(n_377)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_377),
.Y(n_398)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_319),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_378),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_344),
.A2(n_293),
.B(n_311),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_317),
.A2(n_295),
.B1(n_308),
.B2(n_303),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_353),
.A2(n_345),
.B1(n_329),
.B2(n_324),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_382),
.A2(n_401),
.B1(n_378),
.B2(n_376),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_367),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_383),
.B(n_395),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_384),
.B(n_385),
.C(n_388),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_355),
.B(n_351),
.C(n_337),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_356),
.B(n_351),
.C(n_337),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_389),
.A2(n_394),
.B(n_402),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g421 ( 
.A(n_390),
.B(n_392),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_374),
.A2(n_323),
.B(n_333),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_369),
.B(n_321),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_397),
.B(n_403),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g399 ( 
.A(n_362),
.B(n_321),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_363),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_381),
.B(n_360),
.C(n_357),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_400),
.B(n_405),
.C(n_406),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_374),
.A2(n_358),
.B(n_373),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_375),
.B(n_330),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_SL g405 ( 
.A(n_357),
.B(n_328),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_367),
.B(n_363),
.Y(n_406)
);

OAI22xp33_ASAP7_75t_SL g407 ( 
.A1(n_361),
.A2(n_331),
.B1(n_326),
.B2(n_322),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_407),
.A2(n_380),
.B1(n_364),
.B2(n_370),
.Y(n_417)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_404),
.Y(n_408)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_408),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_396),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_409),
.B(n_411),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_396),
.Y(n_411)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_404),
.Y(n_413)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_413),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_383),
.A2(n_361),
.B1(n_379),
.B2(n_365),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_414),
.A2(n_427),
.B1(n_428),
.B2(n_429),
.Y(n_432)
);

MAJx2_ASAP7_75t_L g434 ( 
.A(n_415),
.B(n_393),
.C(n_399),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_417),
.Y(n_437)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_406),
.Y(n_418)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_418),
.Y(n_447)
);

BUFx24_ASAP7_75t_SL g419 ( 
.A(n_392),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_419),
.B(n_424),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_395),
.B(n_352),
.Y(n_420)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_420),
.Y(n_433)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_386),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_384),
.B(n_366),
.C(n_347),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_425),
.B(n_416),
.C(n_423),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_382),
.B(n_352),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_426),
.Y(n_443)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_386),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_398),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_398),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_430),
.A2(n_401),
.B1(n_394),
.B2(n_390),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_434),
.B(n_439),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_435),
.A2(n_448),
.B1(n_414),
.B2(n_420),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_436),
.B(n_441),
.C(n_444),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_426),
.A2(n_402),
.B1(n_400),
.B2(n_389),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_438),
.A2(n_417),
.B1(n_412),
.B2(n_424),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_416),
.B(n_385),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_425),
.B(n_388),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_440),
.B(n_436),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_423),
.B(n_393),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_418),
.B(n_405),
.C(n_387),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_430),
.A2(n_387),
.B1(n_359),
.B2(n_391),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_449),
.B(n_454),
.Y(n_463)
);

BUFx12_ASAP7_75t_L g450 ( 
.A(n_443),
.Y(n_450)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_450),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_451),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_431),
.B(n_410),
.Y(n_454)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_442),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_455),
.B(n_456),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_439),
.B(n_412),
.C(n_415),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_446),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_457),
.A2(n_459),
.B1(n_461),
.B2(n_422),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_437),
.A2(n_427),
.B(n_421),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_458),
.B(n_460),
.Y(n_471)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_433),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_433),
.B(n_410),
.Y(n_460)
);

BUFx12_ASAP7_75t_L g461 ( 
.A(n_432),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_462),
.A2(n_432),
.B1(n_437),
.B2(n_421),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_456),
.B(n_440),
.C(n_441),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_464),
.B(n_465),
.C(n_469),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_453),
.B(n_447),
.C(n_438),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_453),
.B(n_444),
.C(n_409),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_470),
.B(n_461),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_452),
.B(n_435),
.C(n_448),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_472),
.B(n_434),
.C(n_461),
.Y(n_482)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_473),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_463),
.B(n_457),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_474),
.B(n_476),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_468),
.A2(n_462),
.B1(n_454),
.B2(n_458),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_467),
.B(n_455),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_477),
.B(n_480),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_471),
.A2(n_460),
.B(n_459),
.Y(n_478)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_478),
.B(n_481),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_469),
.B(n_452),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_482),
.B(n_464),
.C(n_466),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_479),
.B(n_480),
.C(n_465),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_485),
.B(n_486),
.Y(n_492)
);

INVx6_ASAP7_75t_L g486 ( 
.A(n_479),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_475),
.A2(n_468),
.B(n_472),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_488),
.B(n_478),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_489),
.B(n_482),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_490),
.B(n_483),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_486),
.B(n_481),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_491),
.A2(n_493),
.B1(n_494),
.B2(n_483),
.Y(n_496)
);

BUFx4f_ASAP7_75t_SL g494 ( 
.A(n_485),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_492),
.B(n_484),
.C(n_487),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_495),
.Y(n_498)
);

OAI321xp33_ASAP7_75t_L g499 ( 
.A1(n_496),
.A2(n_497),
.A3(n_450),
.B1(n_429),
.B2(n_445),
.C(n_413),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_499),
.B(n_408),
.C(n_372),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_500),
.A2(n_498),
.B(n_372),
.Y(n_501)
);

OAI21x1_ASAP7_75t_L g502 ( 
.A1(n_501),
.A2(n_391),
.B(n_322),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_502),
.B(n_340),
.Y(n_503)
);


endmodule