module fake_netlist_5_987_n_901 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_901);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_901;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_316;
wire n_855;
wire n_389;
wire n_843;
wire n_785;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_452;
wire n_885;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_841;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_859;
wire n_864;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_854;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_820;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_448;
wire n_259;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_804;
wire n_867;
wire n_537;
wire n_587;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_782;
wire n_325;
wire n_449;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_894;
wire n_271;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_654;
wire n_370;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_255;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_849;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_432;
wire n_395;
wire n_553;
wire n_727;
wire n_839;
wire n_311;
wire n_813;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_277;
wire n_338;
wire n_477;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_557;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_679;
wire n_237;
wire n_513;
wire n_425;
wire n_407;
wire n_527;
wire n_647;
wire n_710;
wire n_707;
wire n_832;
wire n_695;
wire n_795;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_799;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_759;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_143),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_184),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_199),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_50),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_126),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_155),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_120),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_62),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_172),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_42),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_188),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_142),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_12),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_18),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_200),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_88),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_100),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_178),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_46),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_22),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_80),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_56),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_74),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_131),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_2),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_105),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_124),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_154),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_32),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_85),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_34),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_107),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_82),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_122),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_41),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_86),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_79),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_29),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_161),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_10),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_44),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_160),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_69),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_173),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_175),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_87),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_110),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_180),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_19),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_198),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_63),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_47),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_170),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_187),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_83),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_99),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_45),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_5),
.Y(n_263)
);

INVxp33_ASAP7_75t_SL g264 ( 
.A(n_26),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_102),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_148),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_129),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_6),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_158),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_7),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_156),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_133),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_151),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_15),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_191),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_192),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_70),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_157),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_182),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_163),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_186),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_38),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_169),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_211),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_274),
.Y(n_285)
);

INVxp67_ASAP7_75t_SL g286 ( 
.A(n_246),
.Y(n_286)
);

INVxp67_ASAP7_75t_SL g287 ( 
.A(n_220),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

INVxp67_ASAP7_75t_SL g289 ( 
.A(n_220),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_233),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_218),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_225),
.Y(n_292)
);

INVxp67_ASAP7_75t_SL g293 ( 
.A(n_206),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_204),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_232),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_205),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_217),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_208),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_209),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_207),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_216),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_221),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_213),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_283),
.Y(n_304)
);

INVxp33_ASAP7_75t_SL g305 ( 
.A(n_263),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_223),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_226),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_254),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_227),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_214),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_228),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_224),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_235),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_239),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_230),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_242),
.Y(n_316)
);

NOR2xp67_ASAP7_75t_L g317 ( 
.A(n_212),
.B(n_0),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_245),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_268),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_270),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_242),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_264),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_252),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_252),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_247),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_232),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_233),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_256),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_240),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_248),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_215),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_249),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_253),
.B(n_0),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_219),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_265),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_271),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_287),
.B(n_256),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_300),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_325),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_325),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_289),
.B(n_232),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_285),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_326),
.B(n_237),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_318),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_291),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_294),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_301),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_307),
.B(n_269),
.Y(n_348)
);

NAND2xp33_ASAP7_75t_R g349 ( 
.A(n_291),
.B(n_229),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_297),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_296),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_302),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_306),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_309),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_298),
.B(n_212),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_R g356 ( 
.A(n_290),
.B(n_231),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_311),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_313),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_329),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_312),
.Y(n_360)
);

OA21x2_ASAP7_75t_L g361 ( 
.A1(n_330),
.A2(n_260),
.B(n_275),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_284),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_336),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_288),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_293),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_299),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_303),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_335),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_314),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_332),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_333),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_317),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_310),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_331),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_295),
.Y(n_375)
);

AND2x4_ASAP7_75t_L g376 ( 
.A(n_286),
.B(n_260),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_331),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_308),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_295),
.B(n_276),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_334),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_312),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_320),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_315),
.Y(n_383)
);

NAND2xp33_ASAP7_75t_L g384 ( 
.A(n_320),
.B(n_210),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_334),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_292),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_319),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_322),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_322),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_323),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_352),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_386),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_386),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_390),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_354),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_359),
.Y(n_396)
);

BUFx10_ASAP7_75t_L g397 ( 
.A(n_343),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_355),
.B(n_305),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_358),
.Y(n_399)
);

OR2x2_ASAP7_75t_L g400 ( 
.A(n_370),
.B(n_323),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_342),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_370),
.Y(n_402)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_339),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_376),
.B(n_210),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_361),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_342),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_350),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_L g408 ( 
.A1(n_371),
.A2(n_305),
.B1(n_278),
.B2(n_282),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_350),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_358),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_376),
.B(n_210),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_337),
.B(n_234),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_375),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_388),
.B(n_324),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_357),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_383),
.B(n_328),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_387),
.B(n_327),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_337),
.B(n_324),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_358),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_358),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_371),
.B(n_236),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_357),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_376),
.B(n_210),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_361),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_358),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_341),
.B(n_304),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_341),
.B(n_321),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_362),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_363),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_361),
.Y(n_430)
);

BUFx4f_ASAP7_75t_L g431 ( 
.A(n_389),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_L g432 ( 
.A1(n_361),
.A2(n_222),
.B1(n_281),
.B2(n_280),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_346),
.Y(n_433)
);

INVxp67_ASAP7_75t_SL g434 ( 
.A(n_363),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_363),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_363),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_363),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_338),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_364),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_365),
.B(n_238),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_368),
.B(n_369),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_346),
.B(n_316),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_385),
.A2(n_279),
.B1(n_277),
.B2(n_273),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_364),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_338),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_338),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_351),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_347),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_347),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_347),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_353),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_385),
.B(n_222),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_379),
.B(n_241),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_385),
.B(n_222),
.Y(n_454)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_353),
.Y(n_455)
);

AND2x6_ASAP7_75t_L g456 ( 
.A(n_379),
.B(n_222),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_388),
.B(n_243),
.Y(n_457)
);

OR2x2_ASAP7_75t_L g458 ( 
.A(n_344),
.B(n_244),
.Y(n_458)
);

OR2x6_ASAP7_75t_L g459 ( 
.A(n_345),
.B(n_1),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_353),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_351),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_398),
.B(n_374),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_405),
.B(n_424),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_424),
.B(n_379),
.Y(n_464)
);

OAI22xp33_ASAP7_75t_L g465 ( 
.A1(n_400),
.A2(n_377),
.B1(n_374),
.B2(n_380),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_431),
.B(n_366),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_398),
.B(n_377),
.Y(n_467)
);

AO22x1_ASAP7_75t_L g468 ( 
.A1(n_418),
.A2(n_380),
.B1(n_382),
.B2(n_381),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_402),
.B(n_366),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_441),
.A2(n_349),
.B1(n_360),
.B2(n_373),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_450),
.B(n_367),
.Y(n_471)
);

NAND3xp33_ASAP7_75t_L g472 ( 
.A(n_408),
.B(n_421),
.C(n_441),
.Y(n_472)
);

NAND2x1_ASAP7_75t_L g473 ( 
.A(n_430),
.B(n_372),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_407),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_397),
.B(n_367),
.Y(n_475)
);

OAI22xp33_ASAP7_75t_L g476 ( 
.A1(n_412),
.A2(n_373),
.B1(n_339),
.B2(n_340),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_450),
.B(n_384),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_431),
.B(n_340),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_409),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_455),
.B(n_348),
.Y(n_480)
);

NOR3x1_ASAP7_75t_L g481 ( 
.A(n_394),
.B(n_378),
.C(n_1),
.Y(n_481)
);

INVx4_ASAP7_75t_L g482 ( 
.A(n_448),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_397),
.B(n_356),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_415),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_455),
.B(n_432),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_426),
.B(n_378),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_430),
.B(n_250),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_427),
.Y(n_488)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_448),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_397),
.B(n_251),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_391),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_408),
.B(n_255),
.Y(n_492)
);

AND2x4_ASAP7_75t_SL g493 ( 
.A(n_401),
.B(n_257),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_432),
.B(n_258),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g495 ( 
.A1(n_404),
.A2(n_272),
.B1(n_267),
.B2(n_266),
.Y(n_495)
);

A2O1A1Ixp33_ASAP7_75t_SL g496 ( 
.A1(n_399),
.A2(n_262),
.B(n_261),
.C(n_259),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_406),
.B(n_28),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_446),
.B(n_30),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_449),
.B(n_438),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_414),
.B(n_2),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_395),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_448),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_396),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_403),
.B(n_3),
.Y(n_504)
);

NAND3xp33_ASAP7_75t_SL g505 ( 
.A(n_416),
.B(n_3),
.C(n_4),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_457),
.A2(n_101),
.B1(n_202),
.B2(n_201),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_457),
.B(n_4),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_440),
.A2(n_98),
.B1(n_196),
.B2(n_195),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_453),
.A2(n_97),
.B1(n_194),
.B2(n_193),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_438),
.B(n_31),
.Y(n_510)
);

AOI22xp33_ASAP7_75t_L g511 ( 
.A1(n_404),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_445),
.B(n_33),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_415),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_445),
.B(n_35),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_451),
.B(n_36),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_413),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_459),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_416),
.A2(n_106),
.B1(n_190),
.B2(n_189),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_413),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_451),
.B(n_37),
.Y(n_520)
);

INVx2_ASAP7_75t_SL g521 ( 
.A(n_458),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_448),
.B(n_39),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_422),
.Y(n_523)
);

NAND2x1_ASAP7_75t_L g524 ( 
.A(n_399),
.B(n_40),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_460),
.B(n_43),
.Y(n_525)
);

NAND3xp33_ASAP7_75t_L g526 ( 
.A(n_443),
.B(n_8),
.C(n_9),
.Y(n_526)
);

NAND2xp33_ASAP7_75t_L g527 ( 
.A(n_456),
.B(n_460),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_417),
.A2(n_111),
.B1(n_185),
.B2(n_183),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_460),
.B(n_48),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_460),
.B(n_49),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_417),
.A2(n_452),
.B1(n_454),
.B2(n_423),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_433),
.B(n_11),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_422),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_447),
.B(n_11),
.Y(n_534)
);

INVx5_ASAP7_75t_L g535 ( 
.A(n_482),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_516),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_513),
.Y(n_537)
);

INVx1_ASAP7_75t_SL g538 ( 
.A(n_486),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_523),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_533),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_463),
.B(n_411),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_484),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_474),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_502),
.Y(n_544)
);

INVx5_ASAP7_75t_L g545 ( 
.A(n_482),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_479),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_463),
.B(n_411),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_497),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_472),
.B(n_464),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_497),
.Y(n_550)
);

BUFx12f_ASAP7_75t_SL g551 ( 
.A(n_504),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_499),
.Y(n_552)
);

NOR3xp33_ASAP7_75t_SL g553 ( 
.A(n_505),
.B(n_461),
.C(n_452),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_R g554 ( 
.A(n_462),
.B(n_442),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_470),
.B(n_392),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_464),
.B(n_423),
.Y(n_556)
);

BUFx6f_ASAP7_75t_SL g557 ( 
.A(n_521),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_488),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_491),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_485),
.B(n_454),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_501),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_503),
.Y(n_562)
);

INVx6_ASAP7_75t_L g563 ( 
.A(n_500),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_519),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_467),
.B(n_393),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_524),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_507),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_471),
.B(n_493),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_473),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_502),
.Y(n_570)
);

NAND2xp33_ASAP7_75t_L g571 ( 
.A(n_480),
.B(n_456),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_487),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_477),
.Y(n_573)
);

NOR3xp33_ASAP7_75t_SL g574 ( 
.A(n_517),
.B(n_444),
.C(n_439),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_475),
.B(n_428),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_494),
.A2(n_456),
.B1(n_410),
.B2(n_437),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_469),
.B(n_459),
.Y(n_577)
);

NOR3xp33_ASAP7_75t_SL g578 ( 
.A(n_517),
.B(n_459),
.C(n_435),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_466),
.B(n_419),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g580 ( 
.A(n_532),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_489),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_487),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_529),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_R g584 ( 
.A(n_527),
.B(n_529),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_531),
.B(n_434),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_465),
.B(n_419),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_478),
.B(n_429),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_476),
.B(n_495),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_468),
.B(n_429),
.Y(n_589)
);

NOR2xp67_ASAP7_75t_L g590 ( 
.A(n_483),
.B(n_420),
.Y(n_590)
);

NAND2xp33_ASAP7_75t_SL g591 ( 
.A(n_490),
.B(n_425),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_530),
.Y(n_592)
);

INVx5_ASAP7_75t_L g593 ( 
.A(n_496),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_530),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_567),
.A2(n_528),
.B1(n_518),
.B2(n_511),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_565),
.B(n_492),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_567),
.B(n_534),
.Y(n_597)
);

AO31x2_ASAP7_75t_L g598 ( 
.A1(n_585),
.A2(n_525),
.A3(n_522),
.B(n_498),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_543),
.Y(n_599)
);

OR2x6_ASAP7_75t_L g600 ( 
.A(n_558),
.B(n_526),
.Y(n_600)
);

NAND2x1p5_ASAP7_75t_L g601 ( 
.A(n_535),
.B(n_436),
.Y(n_601)
);

INVx5_ASAP7_75t_L g602 ( 
.A(n_535),
.Y(n_602)
);

AO31x2_ASAP7_75t_L g603 ( 
.A1(n_585),
.A2(n_520),
.A3(n_515),
.B(n_514),
.Y(n_603)
);

OAI21x1_ASAP7_75t_L g604 ( 
.A1(n_583),
.A2(n_512),
.B(n_510),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_552),
.B(n_573),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_546),
.Y(n_606)
);

OAI21x1_ASAP7_75t_L g607 ( 
.A1(n_592),
.A2(n_594),
.B(n_549),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_582),
.B(n_456),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_538),
.B(n_481),
.Y(n_609)
);

OAI21xp5_ASAP7_75t_L g610 ( 
.A1(n_549),
.A2(n_506),
.B(n_509),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_572),
.B(n_456),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_538),
.B(n_436),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_535),
.B(n_508),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_L g614 ( 
.A1(n_560),
.A2(n_112),
.B(n_181),
.Y(n_614)
);

OAI21x1_ASAP7_75t_L g615 ( 
.A1(n_556),
.A2(n_570),
.B(n_544),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_535),
.A2(n_109),
.B(n_177),
.Y(n_616)
);

OAI21x1_ASAP7_75t_L g617 ( 
.A1(n_560),
.A2(n_108),
.B(n_176),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_563),
.Y(n_618)
);

OAI21xp5_ASAP7_75t_L g619 ( 
.A1(n_541),
.A2(n_104),
.B(n_174),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_544),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_570),
.Y(n_621)
);

OA21x2_ASAP7_75t_L g622 ( 
.A1(n_541),
.A2(n_103),
.B(n_171),
.Y(n_622)
);

OAI21x1_ASAP7_75t_L g623 ( 
.A1(n_556),
.A2(n_96),
.B(n_168),
.Y(n_623)
);

OAI21xp5_ASAP7_75t_L g624 ( 
.A1(n_547),
.A2(n_95),
.B(n_167),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_575),
.B(n_554),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_542),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_548),
.B(n_12),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_L g628 ( 
.A1(n_547),
.A2(n_94),
.B(n_166),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_548),
.B(n_13),
.Y(n_629)
);

NAND2x1p5_ASAP7_75t_L g630 ( 
.A(n_545),
.B(n_51),
.Y(n_630)
);

BUFx12f_ASAP7_75t_L g631 ( 
.A(n_536),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_548),
.B(n_13),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_580),
.B(n_14),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_550),
.Y(n_634)
);

INVx5_ASAP7_75t_L g635 ( 
.A(n_545),
.Y(n_635)
);

OA21x2_ASAP7_75t_L g636 ( 
.A1(n_576),
.A2(n_113),
.B(n_165),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_550),
.B(n_14),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_537),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_545),
.B(n_52),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_557),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_561),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_550),
.B(n_15),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_599),
.Y(n_643)
);

NAND3xp33_ASAP7_75t_SL g644 ( 
.A(n_596),
.B(n_588),
.C(n_578),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_634),
.B(n_559),
.Y(n_645)
);

AO21x2_ASAP7_75t_L g646 ( 
.A1(n_610),
.A2(n_584),
.B(n_571),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_602),
.A2(n_635),
.B(n_545),
.Y(n_647)
);

AOI21xp33_ASAP7_75t_L g648 ( 
.A1(n_596),
.A2(n_580),
.B(n_555),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_606),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_625),
.B(n_577),
.Y(n_650)
);

AOI21x1_ASAP7_75t_L g651 ( 
.A1(n_613),
.A2(n_590),
.B(n_586),
.Y(n_651)
);

OA21x2_ASAP7_75t_L g652 ( 
.A1(n_607),
.A2(n_539),
.B(n_540),
.Y(n_652)
);

OAI21x1_ASAP7_75t_L g653 ( 
.A1(n_615),
.A2(n_569),
.B(n_587),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_631),
.Y(n_654)
);

OAI21x1_ASAP7_75t_L g655 ( 
.A1(n_607),
.A2(n_581),
.B(n_589),
.Y(n_655)
);

OAI21xp5_ASAP7_75t_L g656 ( 
.A1(n_595),
.A2(n_553),
.B(n_579),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_605),
.B(n_578),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_634),
.B(n_562),
.Y(n_658)
);

OA21x2_ASAP7_75t_L g659 ( 
.A1(n_617),
.A2(n_574),
.B(n_553),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_609),
.B(n_577),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_638),
.Y(n_661)
);

NOR2xp67_ASAP7_75t_L g662 ( 
.A(n_618),
.B(n_568),
.Y(n_662)
);

OAI21x1_ASAP7_75t_L g663 ( 
.A1(n_604),
.A2(n_593),
.B(n_564),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_631),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_600),
.Y(n_665)
);

OAI21x1_ASAP7_75t_L g666 ( 
.A1(n_604),
.A2(n_593),
.B(n_566),
.Y(n_666)
);

A2O1A1Ixp33_ASAP7_75t_L g667 ( 
.A1(n_619),
.A2(n_624),
.B(n_628),
.C(n_614),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_602),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_640),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_638),
.B(n_641),
.Y(n_670)
);

NAND2x1p5_ASAP7_75t_L g671 ( 
.A(n_602),
.B(n_579),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_626),
.Y(n_672)
);

OAI21x1_ASAP7_75t_L g673 ( 
.A1(n_617),
.A2(n_593),
.B(n_566),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_626),
.Y(n_674)
);

NAND2xp33_ASAP7_75t_L g675 ( 
.A(n_602),
.B(n_574),
.Y(n_675)
);

OAI21x1_ASAP7_75t_L g676 ( 
.A1(n_623),
.A2(n_593),
.B(n_566),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_597),
.B(n_568),
.Y(n_677)
);

OA21x2_ASAP7_75t_L g678 ( 
.A1(n_623),
.A2(n_591),
.B(n_563),
.Y(n_678)
);

OAI21x1_ASAP7_75t_L g679 ( 
.A1(n_613),
.A2(n_563),
.B(n_551),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_635),
.Y(n_680)
);

OAI21x1_ASAP7_75t_SL g681 ( 
.A1(n_616),
.A2(n_557),
.B(n_116),
.Y(n_681)
);

CKINVDCx11_ASAP7_75t_R g682 ( 
.A(n_600),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_600),
.A2(n_536),
.B1(n_17),
.B2(n_18),
.Y(n_683)
);

OAI21x1_ASAP7_75t_L g684 ( 
.A1(n_636),
.A2(n_536),
.B(n_115),
.Y(n_684)
);

OAI22xp5_ASAP7_75t_L g685 ( 
.A1(n_635),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_644),
.A2(n_633),
.B1(n_627),
.B2(n_637),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_654),
.Y(n_687)
);

OAI211xp5_ASAP7_75t_SL g688 ( 
.A1(n_648),
.A2(n_642),
.B(n_632),
.C(n_629),
.Y(n_688)
);

AOI221xp5_ASAP7_75t_L g689 ( 
.A1(n_667),
.A2(n_640),
.B1(n_639),
.B2(n_612),
.C(n_608),
.Y(n_689)
);

AO31x2_ASAP7_75t_L g690 ( 
.A1(n_667),
.A2(n_611),
.A3(n_603),
.B(n_598),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_643),
.Y(n_691)
);

CKINVDCx11_ASAP7_75t_R g692 ( 
.A(n_664),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_677),
.B(n_620),
.Y(n_693)
);

BUFx2_ASAP7_75t_L g694 ( 
.A(n_660),
.Y(n_694)
);

BUFx2_ASAP7_75t_L g695 ( 
.A(n_650),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_668),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_656),
.B(n_635),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_649),
.Y(n_698)
);

AOI222xp33_ASAP7_75t_L g699 ( 
.A1(n_683),
.A2(n_639),
.B1(n_621),
.B2(n_620),
.C1(n_22),
.C2(n_23),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_657),
.A2(n_636),
.B1(n_621),
.B2(n_630),
.Y(n_700)
);

OR2x6_ASAP7_75t_L g701 ( 
.A(n_679),
.B(n_630),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_657),
.B(n_598),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_661),
.Y(n_703)
);

AO21x2_ASAP7_75t_L g704 ( 
.A1(n_676),
.A2(n_598),
.B(n_603),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_661),
.B(n_598),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_665),
.A2(n_636),
.B1(n_622),
.B2(n_601),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_670),
.B(n_622),
.Y(n_707)
);

AO21x2_ASAP7_75t_L g708 ( 
.A1(n_676),
.A2(n_603),
.B(n_622),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_682),
.A2(n_601),
.B1(n_603),
.B2(n_21),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_670),
.B(n_16),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_646),
.A2(n_675),
.B(n_666),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_SL g712 ( 
.A1(n_685),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_712)
);

OAI211xp5_ASAP7_75t_SL g713 ( 
.A1(n_682),
.A2(n_20),
.B(n_24),
.C(n_25),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_670),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_675),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_658),
.B(n_27),
.Y(n_716)
);

CKINVDCx6p67_ASAP7_75t_R g717 ( 
.A(n_664),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_658),
.Y(n_718)
);

INVx5_ASAP7_75t_L g719 ( 
.A(n_668),
.Y(n_719)
);

AO31x2_ASAP7_75t_L g720 ( 
.A1(n_672),
.A2(n_27),
.A3(n_203),
.B(n_54),
.Y(n_720)
);

INVx6_ASAP7_75t_L g721 ( 
.A(n_669),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_674),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_652),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_652),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_652),
.Y(n_725)
);

INVx6_ASAP7_75t_L g726 ( 
.A(n_669),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_679),
.A2(n_53),
.B1(n_55),
.B2(n_57),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_SL g728 ( 
.A1(n_659),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_645),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_658),
.B(n_61),
.Y(n_730)
);

INVx4_ASAP7_75t_L g731 ( 
.A(n_668),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_646),
.B(n_164),
.Y(n_732)
);

CKINVDCx8_ASAP7_75t_R g733 ( 
.A(n_645),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_645),
.B(n_64),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_686),
.A2(n_662),
.B1(n_654),
.B2(n_671),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_733),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_693),
.B(n_659),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_721),
.Y(n_738)
);

AO21x2_ASAP7_75t_L g739 ( 
.A1(n_711),
.A2(n_673),
.B(n_663),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_695),
.B(n_651),
.Y(n_740)
);

BUFx2_ASAP7_75t_L g741 ( 
.A(n_718),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_714),
.B(n_680),
.Y(n_742)
);

INVx4_ASAP7_75t_L g743 ( 
.A(n_721),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_699),
.A2(n_659),
.B1(n_681),
.B2(n_671),
.Y(n_744)
);

OAI221xp5_ASAP7_75t_L g745 ( 
.A1(n_715),
.A2(n_678),
.B1(n_680),
.B2(n_647),
.C(n_655),
.Y(n_745)
);

HB1xp67_ASAP7_75t_L g746 ( 
.A(n_691),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_715),
.A2(n_709),
.B1(n_694),
.B2(n_712),
.Y(n_747)
);

OAI21x1_ASAP7_75t_L g748 ( 
.A1(n_711),
.A2(n_663),
.B(n_673),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_699),
.A2(n_655),
.B1(n_684),
.B2(n_653),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_713),
.A2(n_684),
.B1(n_653),
.B2(n_678),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_688),
.A2(n_678),
.B1(n_680),
.B2(n_666),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_716),
.B(n_65),
.Y(n_752)
);

AOI221xp5_ASAP7_75t_L g753 ( 
.A1(n_688),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.C(n_71),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_726),
.Y(n_754)
);

INVx1_ASAP7_75t_SL g755 ( 
.A(n_726),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_697),
.A2(n_72),
.B1(n_73),
.B2(n_75),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_689),
.A2(n_162),
.B1(n_77),
.B2(n_78),
.Y(n_757)
);

OA21x2_ASAP7_75t_L g758 ( 
.A1(n_702),
.A2(n_723),
.B(n_724),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_L g759 ( 
.A1(n_700),
.A2(n_76),
.B1(n_81),
.B2(n_84),
.Y(n_759)
);

NAND2x1_ASAP7_75t_L g760 ( 
.A(n_701),
.B(n_89),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_689),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_698),
.Y(n_762)
);

AOI221xp5_ASAP7_75t_L g763 ( 
.A1(n_702),
.A2(n_93),
.B1(n_114),
.B2(n_117),
.C(n_118),
.Y(n_763)
);

HB1xp67_ASAP7_75t_L g764 ( 
.A(n_722),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_728),
.A2(n_159),
.B1(n_121),
.B2(n_123),
.Y(n_765)
);

BUFx4f_ASAP7_75t_SL g766 ( 
.A(n_717),
.Y(n_766)
);

BUFx4f_ASAP7_75t_SL g767 ( 
.A(n_687),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_729),
.A2(n_710),
.B1(n_732),
.B2(n_734),
.Y(n_768)
);

OAI21xp5_ASAP7_75t_L g769 ( 
.A1(n_732),
.A2(n_119),
.B(n_125),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_710),
.B(n_127),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_703),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_758),
.Y(n_772)
);

OA21x2_ASAP7_75t_L g773 ( 
.A1(n_748),
.A2(n_725),
.B(n_706),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_737),
.B(n_704),
.Y(n_774)
);

INVx3_ASAP7_75t_L g775 ( 
.A(n_758),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_758),
.B(n_707),
.Y(n_776)
);

AND2x4_ASAP7_75t_L g777 ( 
.A(n_762),
.B(n_701),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_746),
.B(n_705),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_771),
.B(n_764),
.Y(n_779)
);

AO31x2_ASAP7_75t_L g780 ( 
.A1(n_740),
.A2(n_708),
.A3(n_704),
.B(n_731),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_768),
.B(n_690),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_739),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_738),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_738),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_739),
.Y(n_785)
);

BUFx2_ASAP7_75t_L g786 ( 
.A(n_741),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_755),
.B(n_692),
.Y(n_787)
);

OR2x2_ASAP7_75t_L g788 ( 
.A(n_749),
.B(n_690),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_736),
.B(n_730),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_745),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_749),
.B(n_690),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_742),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_742),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_747),
.A2(n_701),
.B1(n_727),
.B2(n_687),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_751),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_760),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_751),
.B(n_720),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_738),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_770),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_750),
.B(n_720),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_750),
.B(n_708),
.Y(n_801)
);

OAI31xp33_ASAP7_75t_L g802 ( 
.A1(n_790),
.A2(n_735),
.A3(n_761),
.B(n_757),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_772),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_772),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_772),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_776),
.B(n_720),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_779),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_779),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_787),
.B(n_743),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_R g810 ( 
.A(n_789),
.B(n_766),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_775),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_776),
.B(n_744),
.Y(n_812)
);

BUFx2_ASAP7_75t_L g813 ( 
.A(n_777),
.Y(n_813)
);

OAI221xp5_ASAP7_75t_L g814 ( 
.A1(n_790),
.A2(n_761),
.B1(n_757),
.B2(n_769),
.C(n_765),
.Y(n_814)
);

AOI322xp5_ASAP7_75t_L g815 ( 
.A1(n_790),
.A2(n_753),
.A3(n_765),
.B1(n_763),
.B2(n_736),
.C1(n_752),
.C2(n_738),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_781),
.B(n_754),
.Y(n_816)
);

AOI221xp5_ASAP7_75t_L g817 ( 
.A1(n_800),
.A2(n_756),
.B1(n_759),
.B2(n_687),
.C(n_754),
.Y(n_817)
);

OAI22xp33_ASAP7_75t_L g818 ( 
.A1(n_796),
.A2(n_766),
.B1(n_743),
.B2(n_767),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_799),
.B(n_754),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_807),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_819),
.B(n_786),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_803),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_816),
.B(n_786),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_808),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_805),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_813),
.B(n_777),
.Y(n_826)
);

OR2x2_ASAP7_75t_L g827 ( 
.A(n_812),
.B(n_813),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_816),
.B(n_777),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_805),
.Y(n_829)
);

INVxp67_ASAP7_75t_L g830 ( 
.A(n_806),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_825),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_830),
.B(n_806),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_829),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_820),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_824),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_832),
.B(n_826),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_834),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_835),
.B(n_821),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_833),
.B(n_809),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_838),
.A2(n_814),
.B1(n_830),
.B2(n_827),
.Y(n_840)
);

OAI21xp5_ASAP7_75t_L g841 ( 
.A1(n_837),
.A2(n_815),
.B(n_802),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_839),
.B(n_831),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_842),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_841),
.Y(n_844)
);

NOR3xp33_ASAP7_75t_L g845 ( 
.A(n_840),
.B(n_818),
.C(n_817),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_843),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_844),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_845),
.Y(n_848)
);

NAND2xp33_ASAP7_75t_R g849 ( 
.A(n_844),
.B(n_810),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_848),
.B(n_836),
.Y(n_850)
);

NOR3xp33_ASAP7_75t_L g851 ( 
.A(n_847),
.B(n_846),
.C(n_849),
.Y(n_851)
);

NAND3xp33_ASAP7_75t_L g852 ( 
.A(n_849),
.B(n_754),
.C(n_794),
.Y(n_852)
);

AOI221x1_ASAP7_75t_L g853 ( 
.A1(n_848),
.A2(n_821),
.B1(n_832),
.B2(n_782),
.C(n_826),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_846),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_848),
.A2(n_823),
.B1(n_812),
.B2(n_767),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_848),
.A2(n_799),
.B(n_783),
.Y(n_856)
);

O2A1O1Ixp33_ASAP7_75t_SL g857 ( 
.A1(n_850),
.A2(n_784),
.B(n_783),
.C(n_798),
.Y(n_857)
);

NAND4xp25_ASAP7_75t_L g858 ( 
.A(n_851),
.B(n_799),
.C(n_795),
.D(n_800),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_SL g859 ( 
.A1(n_854),
.A2(n_796),
.B(n_784),
.Y(n_859)
);

OAI211xp5_ASAP7_75t_L g860 ( 
.A1(n_853),
.A2(n_852),
.B(n_856),
.C(n_855),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_851),
.A2(n_796),
.B1(n_795),
.B2(n_777),
.Y(n_861)
);

AOI221xp5_ASAP7_75t_L g862 ( 
.A1(n_851),
.A2(n_801),
.B1(n_797),
.B2(n_791),
.C(n_811),
.Y(n_862)
);

OA22x2_ASAP7_75t_L g863 ( 
.A1(n_853),
.A2(n_828),
.B1(n_811),
.B2(n_822),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_860),
.A2(n_796),
.B(n_822),
.Y(n_864)
);

OAI211xp5_ASAP7_75t_SL g865 ( 
.A1(n_861),
.A2(n_788),
.B(n_782),
.C(n_778),
.Y(n_865)
);

OA22x2_ASAP7_75t_L g866 ( 
.A1(n_859),
.A2(n_804),
.B1(n_803),
.B2(n_801),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_858),
.Y(n_867)
);

O2A1O1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_857),
.A2(n_797),
.B(n_788),
.C(n_801),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_862),
.B(n_804),
.Y(n_869)
);

AOI321xp33_ASAP7_75t_L g870 ( 
.A1(n_863),
.A2(n_801),
.A3(n_791),
.B1(n_781),
.B2(n_778),
.C(n_785),
.Y(n_870)
);

AOI21xp33_ASAP7_75t_SL g871 ( 
.A1(n_860),
.A2(n_128),
.B(n_130),
.Y(n_871)
);

NOR2x1_ASAP7_75t_L g872 ( 
.A(n_867),
.B(n_731),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_864),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_871),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_869),
.Y(n_875)
);

NAND4xp75_ASAP7_75t_L g876 ( 
.A(n_870),
.B(n_785),
.C(n_773),
.D(n_135),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_866),
.Y(n_877)
);

AOI221xp5_ASAP7_75t_SL g878 ( 
.A1(n_868),
.A2(n_865),
.B1(n_796),
.B2(n_785),
.C(n_775),
.Y(n_878)
);

NOR2x1_ASAP7_75t_L g879 ( 
.A(n_867),
.B(n_796),
.Y(n_879)
);

NAND2x1p5_ASAP7_75t_L g880 ( 
.A(n_867),
.B(n_719),
.Y(n_880)
);

OAI221xp5_ASAP7_75t_L g881 ( 
.A1(n_874),
.A2(n_774),
.B1(n_719),
.B2(n_696),
.C(n_775),
.Y(n_881)
);

NAND4xp25_ASAP7_75t_L g882 ( 
.A(n_872),
.B(n_774),
.C(n_792),
.D(n_696),
.Y(n_882)
);

NAND3xp33_ASAP7_75t_L g883 ( 
.A(n_873),
.B(n_719),
.C(n_775),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_877),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_L g885 ( 
.A1(n_880),
.A2(n_793),
.B1(n_792),
.B2(n_773),
.Y(n_885)
);

NOR2xp67_ASAP7_75t_L g886 ( 
.A(n_875),
.B(n_132),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_884),
.Y(n_887)
);

AOI221xp5_ASAP7_75t_L g888 ( 
.A1(n_881),
.A2(n_883),
.B1(n_882),
.B2(n_885),
.C(n_878),
.Y(n_888)
);

NOR3x1_ASAP7_75t_L g889 ( 
.A(n_886),
.B(n_876),
.C(n_879),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_884),
.Y(n_890)
);

INVx5_ASAP7_75t_L g891 ( 
.A(n_886),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_891),
.B(n_780),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_887),
.Y(n_893)
);

NAND2x1_ASAP7_75t_SL g894 ( 
.A(n_890),
.B(n_889),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_894),
.A2(n_893),
.B(n_891),
.Y(n_895)
);

OR3x1_ASAP7_75t_L g896 ( 
.A(n_895),
.B(n_888),
.C(n_892),
.Y(n_896)
);

AOI21xp33_ASAP7_75t_SL g897 ( 
.A1(n_896),
.A2(n_134),
.B(n_136),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_SL g898 ( 
.A1(n_897),
.A2(n_793),
.B1(n_773),
.B2(n_139),
.Y(n_898)
);

AOI222xp33_ASAP7_75t_L g899 ( 
.A1(n_898),
.A2(n_137),
.B1(n_138),
.B2(n_140),
.C1(n_141),
.C2(n_144),
.Y(n_899)
);

AOI221xp5_ASAP7_75t_L g900 ( 
.A1(n_899),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.C(n_149),
.Y(n_900)
);

AOI211xp5_ASAP7_75t_L g901 ( 
.A1(n_900),
.A2(n_150),
.B(n_152),
.C(n_153),
.Y(n_901)
);


endmodule