module fake_netlist_6_2261_n_1787 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1787);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1787;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1737;
wire n_236;
wire n_653;
wire n_1464;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_80),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_30),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_89),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_62),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_154),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_140),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_74),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_96),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_64),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_43),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_97),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_16),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_144),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_43),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_6),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_42),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_126),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_114),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_63),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_106),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_31),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_77),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_98),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_105),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_23),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_41),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_26),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_122),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_88),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_27),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_39),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_93),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_100),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_18),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_19),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_38),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_85),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_149),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_6),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_65),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_156),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_145),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_110),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_87),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_0),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_21),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_84),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_3),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_9),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_127),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_102),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_42),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_86),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_139),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_8),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_135),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_107),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_91),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_26),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_157),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_11),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_3),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_37),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_61),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_108),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_148),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_9),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_101),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_72),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_28),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_81),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_160),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_109),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_153),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_125),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_128),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_7),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_14),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_40),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_17),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_24),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_44),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_50),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_15),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_83),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_60),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_124),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_51),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_7),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_155),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_150),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_120),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_14),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_16),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_4),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_90),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_152),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_121),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_67),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_10),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_24),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_68),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_0),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_94),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_25),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_36),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_33),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_10),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_66),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_39),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_92),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_30),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_18),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_4),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_36),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_38),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_95),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_13),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_50),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_2),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_104),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_133),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_40),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_49),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_112),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_59),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g287 ( 
.A(n_75),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_56),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_2),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_8),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_142),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_143),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_71),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_123),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_78),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_129),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_34),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_137),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_51),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_34),
.Y(n_300)
);

INVx4_ASAP7_75t_R g301 ( 
.A(n_147),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_138),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_111),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_131),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_12),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_52),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_103),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_47),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_69),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_11),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_48),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_99),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_13),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_1),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_22),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_76),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_79),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_32),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_17),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_195),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_198),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_161),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_167),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_231),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_195),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_231),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_195),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_169),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_223),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_223),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_173),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_223),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_224),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_177),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_180),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_182),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_242),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_184),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_243),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_243),
.Y(n_340)
);

BUFx2_ASAP7_75t_SL g341 ( 
.A(n_232),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_188),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_189),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_243),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_248),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_192),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_197),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_248),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_242),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_181),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_200),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_289),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_181),
.Y(n_353)
);

OR2x2_ASAP7_75t_L g354 ( 
.A(n_205),
.B(n_1),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_176),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_289),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_236),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_202),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_164),
.B(n_5),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_205),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_304),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_171),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_168),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_168),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_208),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_208),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_174),
.Y(n_367)
);

NOR2xp67_ASAP7_75t_L g368 ( 
.A(n_176),
.B(n_5),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_174),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_238),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_238),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_241),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_241),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_265),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_285),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_164),
.B(n_12),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_285),
.Y(n_377)
);

INVxp33_ASAP7_75t_L g378 ( 
.A(n_265),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_273),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_166),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_203),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_207),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_273),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_283),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_165),
.B(n_15),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_210),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_283),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_288),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_268),
.Y(n_389)
);

NOR2xp67_ASAP7_75t_L g390 ( 
.A(n_240),
.B(n_19),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_288),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_240),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_290),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_268),
.Y(n_394)
);

INVxp33_ASAP7_75t_SL g395 ( 
.A(n_172),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_320),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_389),
.A2(n_162),
.B1(n_170),
.B2(n_194),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_320),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_325),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_325),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_329),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_329),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_330),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_330),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_332),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_332),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_339),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_339),
.Y(n_408)
);

NAND2xp33_ASAP7_75t_L g409 ( 
.A(n_354),
.B(n_272),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_340),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_340),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_344),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_367),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_344),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_327),
.B(n_171),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_345),
.Y(n_416)
);

AND2x2_ASAP7_75t_SL g417 ( 
.A(n_359),
.B(n_235),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_345),
.Y(n_418)
);

AND2x6_ASAP7_75t_L g419 ( 
.A(n_376),
.B(n_235),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_348),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_348),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_352),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_352),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_356),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_356),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_327),
.Y(n_426)
);

BUFx8_ASAP7_75t_L g427 ( 
.A(n_369),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_360),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_362),
.B(n_171),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_360),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_350),
.B(n_269),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_350),
.B(n_213),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_365),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_365),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_366),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_366),
.Y(n_436)
);

AND2x6_ASAP7_75t_L g437 ( 
.A(n_385),
.B(n_235),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_353),
.B(n_269),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_371),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_353),
.B(n_269),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_370),
.B(n_214),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_371),
.Y(n_442)
);

OR2x6_ASAP7_75t_L g443 ( 
.A(n_341),
.B(n_296),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_349),
.A2(n_261),
.B1(n_278),
.B2(n_255),
.Y(n_444)
);

AND3x1_ASAP7_75t_L g445 ( 
.A(n_394),
.B(n_272),
.C(n_290),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_370),
.B(n_324),
.Y(n_446)
);

OAI21x1_ASAP7_75t_L g447 ( 
.A1(n_354),
.A2(n_201),
.B(n_178),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_372),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_326),
.B(n_296),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_372),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_373),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_373),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_374),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_374),
.B(n_296),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_379),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_379),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_383),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_383),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_369),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_384),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_384),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_387),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_337),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_387),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_388),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_388),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_391),
.B(n_165),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_446),
.B(n_322),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_417),
.A2(n_349),
.B1(n_368),
.B2(n_390),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_433),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_427),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_446),
.B(n_323),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_426),
.B(n_395),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g474 ( 
.A(n_415),
.Y(n_474)
);

INVx2_ASAP7_75t_SL g475 ( 
.A(n_415),
.Y(n_475)
);

BUFx4f_ASAP7_75t_L g476 ( 
.A(n_417),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_430),
.Y(n_477)
);

INVxp67_ASAP7_75t_SL g478 ( 
.A(n_426),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_426),
.B(n_328),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_398),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_398),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_450),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_398),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_398),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_450),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_431),
.B(n_391),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_399),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_433),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_399),
.Y(n_489)
);

AND2x6_ASAP7_75t_L g490 ( 
.A(n_415),
.B(n_235),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_399),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_446),
.B(n_331),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_463),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_399),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_427),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_415),
.Y(n_496)
);

CKINVDCx16_ASAP7_75t_R g497 ( 
.A(n_443),
.Y(n_497)
);

OAI22x1_ASAP7_75t_L g498 ( 
.A1(n_463),
.A2(n_459),
.B1(n_413),
.B2(n_444),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_400),
.Y(n_499)
);

AND2x6_ASAP7_75t_L g500 ( 
.A(n_415),
.B(n_235),
.Y(n_500)
);

AND2x2_ASAP7_75t_SL g501 ( 
.A(n_417),
.B(n_178),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_400),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_450),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_427),
.Y(n_504)
);

AND2x6_ASAP7_75t_L g505 ( 
.A(n_415),
.B(n_235),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_432),
.B(n_334),
.Y(n_506)
);

AND3x2_ASAP7_75t_L g507 ( 
.A(n_459),
.B(n_225),
.C(n_201),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_430),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_432),
.B(n_335),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_445),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_451),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_400),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_429),
.Y(n_513)
);

INVx4_ASAP7_75t_L g514 ( 
.A(n_430),
.Y(n_514)
);

INVx1_ASAP7_75t_SL g515 ( 
.A(n_449),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_429),
.B(n_179),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_429),
.B(n_336),
.Y(n_517)
);

INVx2_ASAP7_75t_SL g518 ( 
.A(n_429),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_441),
.B(n_338),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_441),
.B(n_389),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_429),
.B(n_342),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_429),
.B(n_343),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_438),
.B(n_346),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_438),
.B(n_347),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_445),
.B(n_351),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_439),
.Y(n_526)
);

OAI22xp33_ASAP7_75t_L g527 ( 
.A1(n_443),
.A2(n_368),
.B1(n_390),
.B2(n_378),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_430),
.Y(n_528)
);

INVx6_ASAP7_75t_L g529 ( 
.A(n_438),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_438),
.B(n_358),
.Y(n_530)
);

CKINVDCx6p67_ASAP7_75t_R g531 ( 
.A(n_443),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_438),
.B(n_381),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_438),
.B(n_382),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_430),
.Y(n_534)
);

INVxp33_ASAP7_75t_L g535 ( 
.A(n_397),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_431),
.B(n_393),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_439),
.Y(n_537)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_430),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_431),
.B(n_386),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_R g540 ( 
.A(n_409),
.B(n_321),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_417),
.B(n_380),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_419),
.A2(n_300),
.B1(n_314),
.B2(n_306),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_442),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_400),
.Y(n_544)
);

INVx6_ASAP7_75t_L g545 ( 
.A(n_467),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_442),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_427),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_430),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_419),
.A2(n_300),
.B1(n_314),
.B2(n_306),
.Y(n_549)
);

BUFx10_ASAP7_75t_L g550 ( 
.A(n_443),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_440),
.B(n_163),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_402),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_449),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_449),
.B(n_363),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_427),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_447),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_447),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_466),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_440),
.B(n_364),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_440),
.B(n_277),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_427),
.B(n_375),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_451),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_402),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_467),
.B(n_393),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_419),
.B(n_216),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_451),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_430),
.Y(n_567)
);

OR2x2_ASAP7_75t_L g568 ( 
.A(n_413),
.B(n_341),
.Y(n_568)
);

OR2x6_ASAP7_75t_L g569 ( 
.A(n_443),
.B(n_299),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_419),
.A2(n_299),
.B1(n_305),
.B2(n_315),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_452),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g572 ( 
.A(n_444),
.B(n_355),
.Y(n_572)
);

AO22x2_ASAP7_75t_L g573 ( 
.A1(n_467),
.A2(n_305),
.B1(n_315),
.B2(n_317),
.Y(n_573)
);

OR2x6_ASAP7_75t_L g574 ( 
.A(n_443),
.B(n_179),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_430),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_452),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_447),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_452),
.Y(n_578)
);

INVx8_ASAP7_75t_L g579 ( 
.A(n_443),
.Y(n_579)
);

NAND2xp33_ASAP7_75t_L g580 ( 
.A(n_419),
.B(n_225),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_407),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_447),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_402),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_453),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_454),
.B(n_355),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_454),
.Y(n_586)
);

AND2x6_ASAP7_75t_L g587 ( 
.A(n_454),
.B(n_245),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_SL g588 ( 
.A1(n_409),
.A2(n_377),
.B1(n_361),
.B2(n_357),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_419),
.B(n_437),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_402),
.Y(n_590)
);

OR2x2_ASAP7_75t_L g591 ( 
.A(n_443),
.B(n_392),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_466),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_453),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_404),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_453),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_456),
.B(n_392),
.Y(n_596)
);

BUFx4f_ASAP7_75t_L g597 ( 
.A(n_419),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_419),
.A2(n_333),
.B1(n_312),
.B2(n_309),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_418),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_418),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_404),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_419),
.B(n_217),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_456),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_456),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_460),
.B(n_462),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_460),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_419),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_419),
.A2(n_245),
.B1(n_282),
.B2(n_316),
.Y(n_608)
);

INVx6_ASAP7_75t_L g609 ( 
.A(n_407),
.Y(n_609)
);

AO21x2_ASAP7_75t_L g610 ( 
.A1(n_460),
.A2(n_317),
.B(n_316),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_462),
.B(n_183),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_462),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_404),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_419),
.A2(n_282),
.B1(n_211),
.B2(n_204),
.Y(n_614)
);

INVx5_ASAP7_75t_L g615 ( 
.A(n_437),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_464),
.Y(n_616)
);

INVx4_ASAP7_75t_L g617 ( 
.A(n_407),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_464),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_496),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_496),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_506),
.B(n_437),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_585),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_539),
.B(n_175),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_501),
.B(n_437),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_501),
.B(n_437),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_545),
.B(n_437),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_476),
.A2(n_437),
.B1(n_234),
.B2(n_193),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_515),
.B(n_464),
.Y(n_628)
);

INVx5_ASAP7_75t_L g629 ( 
.A(n_490),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_479),
.B(n_185),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_545),
.B(n_437),
.Y(n_631)
);

INVxp33_ASAP7_75t_L g632 ( 
.A(n_493),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_545),
.B(n_437),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_545),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_480),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_L g636 ( 
.A1(n_476),
.A2(n_437),
.B(n_193),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_568),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_585),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_481),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_553),
.B(n_218),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_553),
.B(n_186),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_513),
.Y(n_642)
);

NOR2xp67_ASAP7_75t_L g643 ( 
.A(n_471),
.B(n_416),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_473),
.B(n_187),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_586),
.B(n_437),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_586),
.B(n_437),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_520),
.B(n_190),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_520),
.B(n_191),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_592),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_529),
.Y(n_650)
);

O2A1O1Ixp33_ASAP7_75t_L g651 ( 
.A1(n_551),
.A2(n_465),
.B(n_461),
.C(n_458),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_592),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_564),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_486),
.B(n_416),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_513),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_541),
.A2(n_251),
.B1(n_226),
.B2(n_228),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_474),
.B(n_424),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_486),
.B(n_416),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_474),
.B(n_424),
.Y(n_659)
);

INVx8_ASAP7_75t_L g660 ( 
.A(n_579),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_475),
.B(n_478),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_475),
.B(n_424),
.Y(n_662)
);

OAI21xp33_ASAP7_75t_L g663 ( 
.A1(n_469),
.A2(n_199),
.B(n_196),
.Y(n_663)
);

BUFx6f_ASAP7_75t_SL g664 ( 
.A(n_611),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_518),
.B(n_424),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_481),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_468),
.B(n_206),
.Y(n_667)
);

AND2x6_ASAP7_75t_L g668 ( 
.A(n_556),
.B(n_183),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_577),
.Y(n_669)
);

NOR3xp33_ASAP7_75t_L g670 ( 
.A(n_559),
.B(n_397),
.C(n_211),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_518),
.B(n_424),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_470),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_523),
.B(n_424),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_488),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_472),
.B(n_209),
.Y(n_675)
);

INVx8_ASAP7_75t_L g676 ( 
.A(n_579),
.Y(n_676)
);

NAND2xp33_ASAP7_75t_SL g677 ( 
.A(n_540),
.B(n_212),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_492),
.B(n_215),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_529),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_483),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_564),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_536),
.B(n_428),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_560),
.B(n_219),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_524),
.B(n_221),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_484),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_484),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_533),
.B(n_517),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_536),
.B(n_420),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_487),
.Y(n_689)
);

INVxp67_ASAP7_75t_L g690 ( 
.A(n_596),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_595),
.B(n_428),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_591),
.B(n_250),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_595),
.B(n_428),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_487),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_611),
.B(n_204),
.Y(n_695)
);

BUFx5_ASAP7_75t_L g696 ( 
.A(n_556),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_611),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_476),
.A2(n_258),
.B1(n_252),
.B2(n_256),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_605),
.B(n_428),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_529),
.B(n_434),
.Y(n_700)
);

INVxp67_ASAP7_75t_L g701 ( 
.A(n_591),
.Y(n_701)
);

BUFx4f_ASAP7_75t_L g702 ( 
.A(n_568),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_529),
.B(n_434),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_482),
.B(n_434),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_521),
.B(n_222),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_482),
.B(n_434),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_526),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_489),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_527),
.B(n_257),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_485),
.B(n_435),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_485),
.B(n_435),
.Y(n_711)
);

INVx8_ASAP7_75t_L g712 ( 
.A(n_579),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_503),
.B(n_435),
.Y(n_713)
);

NOR2xp67_ASAP7_75t_L g714 ( 
.A(n_471),
.B(n_420),
.Y(n_714)
);

O2A1O1Ixp33_ASAP7_75t_L g715 ( 
.A1(n_530),
.A2(n_532),
.B(n_580),
.C(n_511),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_L g716 ( 
.A1(n_497),
.A2(n_293),
.B1(n_229),
.B2(n_233),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_537),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_522),
.B(n_227),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_531),
.A2(n_293),
.B1(n_229),
.B2(n_233),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_503),
.B(n_435),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_577),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_R g722 ( 
.A(n_495),
.B(n_259),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_554),
.B(n_420),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_597),
.B(n_262),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_573),
.A2(n_220),
.B1(n_234),
.B2(n_246),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_511),
.B(n_436),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_597),
.B(n_264),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_598),
.B(n_271),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_489),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_509),
.B(n_291),
.Y(n_730)
);

NAND3xp33_ASAP7_75t_L g731 ( 
.A(n_525),
.B(n_254),
.C(n_230),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_577),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_491),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_543),
.B(n_220),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_519),
.B(n_292),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_491),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_562),
.B(n_436),
.Y(n_737)
);

AO22x2_ASAP7_75t_L g738 ( 
.A1(n_572),
.A2(n_307),
.B1(n_247),
.B2(n_281),
.Y(n_738)
);

INVxp67_ASAP7_75t_L g739 ( 
.A(n_510),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_510),
.B(n_237),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_494),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_562),
.B(n_436),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_546),
.Y(n_743)
);

INVx8_ASAP7_75t_L g744 ( 
.A(n_579),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_566),
.B(n_436),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_566),
.B(n_448),
.Y(n_746)
);

BUFx5_ASAP7_75t_L g747 ( 
.A(n_557),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_588),
.B(n_425),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_597),
.B(n_298),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_571),
.B(n_448),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_571),
.B(n_448),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_516),
.A2(n_302),
.B1(n_247),
.B2(n_281),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_558),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_494),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_573),
.A2(n_246),
.B1(n_294),
.B2(n_295),
.Y(n_755)
);

INVx8_ASAP7_75t_L g756 ( 
.A(n_569),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_576),
.B(n_448),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_576),
.B(n_455),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_578),
.B(n_455),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_550),
.B(n_286),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_572),
.B(n_425),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_L g762 ( 
.A1(n_531),
.A2(n_294),
.B1(n_295),
.B2(n_303),
.Y(n_762)
);

AOI221xp5_ASAP7_75t_L g763 ( 
.A1(n_498),
.A2(n_249),
.B1(n_239),
.B2(n_319),
.C(n_318),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_612),
.B(n_244),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_615),
.B(n_418),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_615),
.B(n_418),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_507),
.Y(n_767)
);

A2O1A1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_516),
.A2(n_307),
.B(n_303),
.C(n_411),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_615),
.B(n_418),
.Y(n_769)
);

OR2x6_ASAP7_75t_SL g770 ( 
.A(n_495),
.B(n_253),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_499),
.Y(n_771)
);

INVx8_ASAP7_75t_L g772 ( 
.A(n_569),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_498),
.B(n_260),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_550),
.B(n_286),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_584),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_499),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_616),
.B(n_263),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_593),
.B(n_455),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_593),
.B(n_455),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_516),
.Y(n_780)
);

INVxp67_ASAP7_75t_L g781 ( 
.A(n_610),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_603),
.Y(n_782)
);

INVx8_ASAP7_75t_L g783 ( 
.A(n_569),
.Y(n_783)
);

NAND2xp33_ASAP7_75t_L g784 ( 
.A(n_587),
.B(n_577),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_603),
.B(n_457),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_604),
.B(n_457),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_615),
.B(n_418),
.Y(n_787)
);

BUFx2_ASAP7_75t_L g788 ( 
.A(n_739),
.Y(n_788)
);

BUFx8_ASAP7_75t_SL g789 ( 
.A(n_702),
.Y(n_789)
);

O2A1O1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_690),
.A2(n_618),
.B(n_604),
.C(n_606),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_687),
.A2(n_587),
.B1(n_569),
.B2(n_574),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_687),
.B(n_606),
.Y(n_792)
);

NAND2x1p5_ASAP7_75t_L g793 ( 
.A(n_669),
.B(n_607),
.Y(n_793)
);

AND2x4_ASAP7_75t_L g794 ( 
.A(n_653),
.B(n_547),
.Y(n_794)
);

O2A1O1Ixp5_ASAP7_75t_L g795 ( 
.A1(n_673),
.A2(n_618),
.B(n_565),
.C(n_602),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_644),
.A2(n_587),
.B1(n_574),
.B2(n_607),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_690),
.B(n_577),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_624),
.A2(n_557),
.B1(n_582),
.B2(n_574),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_669),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_701),
.Y(n_800)
);

OAI21xp5_ASAP7_75t_L g801 ( 
.A1(n_625),
.A2(n_589),
.B(n_582),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_644),
.A2(n_587),
.B1(n_574),
.B2(n_550),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_784),
.A2(n_615),
.B(n_580),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_630),
.B(n_587),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_630),
.B(n_587),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_701),
.Y(n_806)
);

O2A1O1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_622),
.A2(n_610),
.B(n_561),
.C(n_542),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_661),
.A2(n_514),
.B(n_538),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_636),
.A2(n_514),
.B(n_538),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_628),
.B(n_547),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_775),
.Y(n_811)
);

AOI21x1_ASAP7_75t_L g812 ( 
.A1(n_724),
.A2(n_749),
.B(n_727),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_782),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_700),
.A2(n_514),
.B(n_538),
.Y(n_814)
);

AOI21x1_ASAP7_75t_L g815 ( 
.A1(n_724),
.A2(n_502),
.B(n_512),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_654),
.B(n_573),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_619),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_703),
.A2(n_617),
.B(n_608),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_681),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_658),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_781),
.A2(n_614),
.B(n_570),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_626),
.A2(n_617),
.B(n_508),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_L g823 ( 
.A1(n_627),
.A2(n_504),
.B1(n_555),
.B2(n_549),
.Y(n_823)
);

NOR2xp67_ASAP7_75t_L g824 ( 
.A(n_731),
.B(n_656),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_631),
.A2(n_617),
.B(n_575),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_688),
.B(n_573),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_633),
.A2(n_575),
.B(n_528),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_669),
.A2(n_575),
.B(n_528),
.Y(n_828)
);

A2O1A1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_715),
.A2(n_535),
.B(n_504),
.C(n_555),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_638),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_620),
.Y(n_831)
);

NOR2x1_ASAP7_75t_L g832 ( 
.A(n_643),
.B(n_610),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_683),
.B(n_490),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_632),
.B(n_266),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_702),
.B(n_508),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_683),
.A2(n_477),
.B(n_534),
.C(n_548),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_642),
.B(n_508),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_669),
.A2(n_528),
.B(n_575),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_623),
.B(n_684),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_699),
.A2(n_528),
.B(n_575),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_627),
.A2(n_548),
.B1(n_477),
.B2(n_534),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_L g842 ( 
.A1(n_781),
.A2(n_500),
.B(n_505),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_650),
.A2(n_508),
.B(n_528),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_697),
.B(n_425),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_623),
.B(n_490),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_650),
.A2(n_508),
.B(n_477),
.Y(n_846)
);

AOI21x1_ASAP7_75t_L g847 ( 
.A1(n_727),
.A2(n_613),
.B(n_502),
.Y(n_847)
);

O2A1O1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_709),
.A2(n_613),
.B(n_601),
.C(n_594),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_684),
.B(n_490),
.Y(n_849)
);

OR2x6_ASAP7_75t_SL g850 ( 
.A(n_716),
.B(n_267),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_705),
.B(n_490),
.Y(n_851)
);

BUFx4f_ASAP7_75t_L g852 ( 
.A(n_756),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_682),
.A2(n_548),
.B(n_567),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_SL g854 ( 
.A(n_637),
.B(n_286),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_665),
.A2(n_534),
.B(n_567),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_705),
.A2(n_505),
.B1(n_490),
.B2(n_500),
.Y(n_856)
);

BUFx8_ASAP7_75t_SL g857 ( 
.A(n_664),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_635),
.Y(n_858)
);

NAND2xp33_ASAP7_75t_SL g859 ( 
.A(n_722),
.B(n_270),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_739),
.B(n_567),
.Y(n_860)
);

NAND2xp33_ASAP7_75t_L g861 ( 
.A(n_660),
.B(n_500),
.Y(n_861)
);

O2A1O1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_761),
.A2(n_563),
.B(n_601),
.C(n_594),
.Y(n_862)
);

O2A1O1Ixp5_ASAP7_75t_L g863 ( 
.A1(n_621),
.A2(n_563),
.B(n_512),
.C(n_544),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_671),
.A2(n_600),
.B(n_599),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_718),
.B(n_500),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_672),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_718),
.B(n_500),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_647),
.B(n_274),
.Y(n_868)
);

BUFx12f_ASAP7_75t_L g869 ( 
.A(n_767),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_740),
.B(n_275),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_740),
.B(n_276),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_641),
.B(n_500),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_657),
.A2(n_600),
.B(n_599),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_780),
.A2(n_609),
.B1(n_581),
.B2(n_583),
.Y(n_874)
);

NOR3xp33_ASAP7_75t_L g875 ( 
.A(n_670),
.B(n_279),
.C(n_280),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_639),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_674),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_707),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_659),
.A2(n_600),
.B(n_599),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_642),
.B(n_286),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_641),
.B(n_505),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_717),
.B(n_505),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_642),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_642),
.Y(n_884)
);

OAI21xp5_ASAP7_75t_L g885 ( 
.A1(n_645),
.A2(n_505),
.B(n_552),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_743),
.B(n_505),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_655),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_725),
.A2(n_287),
.B1(n_590),
.B2(n_583),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_646),
.A2(n_544),
.B(n_552),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_662),
.A2(n_749),
.B(n_693),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_753),
.B(n_581),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_660),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_660),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_723),
.B(n_581),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_691),
.A2(n_600),
.B(n_599),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_679),
.A2(n_600),
.B(n_599),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_667),
.B(n_284),
.Y(n_897)
);

INVxp67_ASAP7_75t_L g898 ( 
.A(n_748),
.Y(n_898)
);

A2O1A1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_667),
.A2(n_590),
.B(n_406),
.C(n_411),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_655),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_679),
.A2(n_732),
.B(n_721),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_649),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_634),
.B(n_652),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_676),
.Y(n_904)
);

INVxp67_ASAP7_75t_L g905 ( 
.A(n_647),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_721),
.A2(n_457),
.B(n_465),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_675),
.A2(n_406),
.B(n_411),
.C(n_461),
.Y(n_907)
);

A2O1A1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_675),
.A2(n_406),
.B(n_411),
.C(n_461),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_732),
.A2(n_457),
.B(n_465),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_651),
.A2(n_465),
.B(n_461),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_629),
.A2(n_458),
.B(n_404),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_695),
.B(n_458),
.Y(n_912)
);

NOR3xp33_ASAP7_75t_L g913 ( 
.A(n_670),
.B(n_297),
.C(n_313),
.Y(n_913)
);

A2O1A1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_678),
.A2(n_406),
.B(n_411),
.C(n_458),
.Y(n_914)
);

INVx6_ASAP7_75t_L g915 ( 
.A(n_655),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_629),
.A2(n_414),
.B(n_406),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_655),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_629),
.A2(n_414),
.B(n_406),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_704),
.A2(n_411),
.B(n_396),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_678),
.A2(n_408),
.B(n_410),
.C(n_396),
.Y(n_920)
);

O2A1O1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_728),
.A2(n_403),
.B(n_412),
.C(n_410),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_648),
.B(n_308),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_695),
.B(n_408),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_648),
.A2(n_408),
.B(n_410),
.C(n_396),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_764),
.B(n_777),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_773),
.B(n_311),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_664),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_L g928 ( 
.A1(n_725),
.A2(n_609),
.B1(n_310),
.B2(n_401),
.Y(n_928)
);

OAI321xp33_ASAP7_75t_L g929 ( 
.A1(n_763),
.A2(n_401),
.A3(n_403),
.B1(n_405),
.B2(n_412),
.C(n_423),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_629),
.B(n_287),
.Y(n_930)
);

O2A1O1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_692),
.A2(n_755),
.B(n_768),
.C(n_762),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_787),
.A2(n_414),
.B(n_401),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_787),
.A2(n_765),
.B(n_766),
.Y(n_933)
);

OAI21xp33_ASAP7_75t_L g934 ( 
.A1(n_663),
.A2(n_412),
.B(n_405),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_666),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_765),
.A2(n_414),
.B(n_403),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_680),
.Y(n_937)
);

BUFx12f_ASAP7_75t_L g938 ( 
.A(n_734),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_764),
.B(n_405),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_766),
.A2(n_423),
.B(n_407),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_706),
.A2(n_423),
.B(n_609),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_685),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_769),
.A2(n_423),
.B(n_407),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_686),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_710),
.A2(n_609),
.B(n_301),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_769),
.A2(n_407),
.B(n_301),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_777),
.B(n_422),
.Y(n_947)
);

O2A1O1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_755),
.A2(n_287),
.B(n_21),
.C(n_22),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_752),
.A2(n_422),
.B(n_421),
.C(n_418),
.Y(n_949)
);

NOR2x1_ASAP7_75t_L g950 ( 
.A(n_714),
.B(n_422),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_698),
.B(n_287),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_734),
.B(n_422),
.Y(n_952)
);

NAND2xp33_ASAP7_75t_L g953 ( 
.A(n_676),
.B(n_422),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_696),
.B(n_421),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_696),
.B(n_422),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_696),
.B(n_422),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_640),
.B(n_20),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_711),
.A2(n_407),
.B(n_421),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_689),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_696),
.B(n_422),
.Y(n_960)
);

INVxp67_ASAP7_75t_SL g961 ( 
.A(n_696),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_696),
.B(n_422),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_713),
.A2(n_407),
.B(n_421),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_738),
.B(n_722),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_720),
.A2(n_407),
.B(n_421),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_738),
.B(n_421),
.Y(n_966)
);

INVx4_ASAP7_75t_L g967 ( 
.A(n_676),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_747),
.B(n_421),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_712),
.Y(n_969)
);

NOR3xp33_ASAP7_75t_L g970 ( 
.A(n_677),
.B(n_20),
.C(n_23),
.Y(n_970)
);

A2O1A1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_760),
.A2(n_421),
.B(n_418),
.C(n_28),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_747),
.B(n_421),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_747),
.B(n_418),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_747),
.B(n_159),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_726),
.A2(n_158),
.B(n_151),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_747),
.B(n_25),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_892),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_892),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_839),
.B(n_747),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_915),
.Y(n_980)
);

O2A1O1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_925),
.A2(n_719),
.B(n_774),
.C(n_735),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_792),
.B(n_737),
.Y(n_982)
);

AND2x2_ASAP7_75t_SL g983 ( 
.A(n_897),
.B(n_770),
.Y(n_983)
);

BUFx3_ASAP7_75t_L g984 ( 
.A(n_869),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_SL g985 ( 
.A(n_789),
.B(n_756),
.Y(n_985)
);

HB1xp67_ASAP7_75t_L g986 ( 
.A(n_819),
.Y(n_986)
);

INVxp67_ASAP7_75t_L g987 ( 
.A(n_788),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_922),
.A2(n_870),
.B(n_871),
.C(n_957),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_898),
.B(n_742),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_794),
.B(n_730),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_898),
.B(n_905),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_905),
.B(n_783),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_857),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_809),
.A2(n_712),
.B(n_744),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_797),
.B(n_786),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_L g996 ( 
.A1(n_820),
.A2(n_738),
.B1(n_783),
.B2(n_756),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_870),
.A2(n_871),
.B(n_922),
.C(n_957),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_961),
.A2(n_712),
.B(n_744),
.Y(n_998)
);

NOR4xp25_ASAP7_75t_SL g999 ( 
.A(n_951),
.B(n_668),
.C(n_772),
.D(n_783),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_892),
.Y(n_1000)
);

A2O1A1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_931),
.A2(n_772),
.B(n_744),
.C(n_778),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_811),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_939),
.B(n_785),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_807),
.A2(n_772),
.B(n_750),
.C(n_779),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_810),
.B(n_745),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_866),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_794),
.B(n_746),
.Y(n_1007)
);

INVxp67_ASAP7_75t_L g1008 ( 
.A(n_819),
.Y(n_1008)
);

BUFx2_ASAP7_75t_L g1009 ( 
.A(n_938),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_868),
.B(n_751),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_813),
.B(n_668),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_877),
.B(n_668),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_875),
.A2(n_757),
.B(n_758),
.C(n_759),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_800),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_875),
.A2(n_776),
.B(n_771),
.C(n_754),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_913),
.B(n_741),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_961),
.A2(n_805),
.B(n_804),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_SL g1018 ( 
.A(n_852),
.B(n_668),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_878),
.B(n_668),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_816),
.A2(n_733),
.B1(n_729),
.B2(n_708),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_912),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_923),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_894),
.B(n_826),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_945),
.A2(n_736),
.B(n_694),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_860),
.B(n_146),
.Y(n_1025)
);

INVx2_ASAP7_75t_SL g1026 ( 
.A(n_830),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_800),
.B(n_27),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_R g1028 ( 
.A(n_859),
.B(n_141),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_892),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_830),
.B(n_29),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_926),
.A2(n_29),
.B(n_31),
.C(n_32),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_893),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_860),
.B(n_136),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_913),
.A2(n_134),
.B1(n_132),
.B2(n_130),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_953),
.A2(n_119),
.B(n_118),
.Y(n_1035)
);

INVx3_ASAP7_75t_L g1036 ( 
.A(n_883),
.Y(n_1036)
);

BUFx3_ASAP7_75t_L g1037 ( 
.A(n_927),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_806),
.B(n_926),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_806),
.B(n_33),
.Y(n_1039)
);

OR2x6_ASAP7_75t_L g1040 ( 
.A(n_927),
.B(n_117),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_801),
.A2(n_116),
.B(n_115),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_791),
.A2(n_35),
.B1(n_37),
.B2(n_41),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_831),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_803),
.A2(n_113),
.B(n_82),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_858),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_937),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_790),
.B(n_73),
.Y(n_1047)
);

BUFx2_ASAP7_75t_R g1048 ( 
.A(n_850),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_876),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_955),
.A2(n_70),
.B(n_44),
.Y(n_1050)
);

NAND3xp33_ASAP7_75t_SL g1051 ( 
.A(n_854),
.B(n_58),
.C(n_45),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_956),
.A2(n_962),
.B(n_960),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_834),
.B(n_35),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_968),
.A2(n_45),
.B(n_46),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_884),
.B(n_46),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_884),
.B(n_47),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_973),
.A2(n_58),
.B(n_49),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_821),
.B(n_48),
.Y(n_1058)
);

INVxp67_ASAP7_75t_SL g1059 ( 
.A(n_799),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_967),
.B(n_893),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_SL g1061 ( 
.A1(n_902),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_1061)
);

NAND3xp33_ASAP7_75t_SL g1062 ( 
.A(n_970),
.B(n_57),
.C(n_54),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_844),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_893),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_935),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_942),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_964),
.B(n_53),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_944),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_903),
.B(n_55),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_959),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_852),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_844),
.B(n_55),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_890),
.A2(n_56),
.B(n_57),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_824),
.A2(n_796),
.B(n_948),
.C(n_802),
.Y(n_1074)
);

OAI22xp33_ASAP7_75t_L g1075 ( 
.A1(n_823),
.A2(n_817),
.B1(n_929),
.B2(n_833),
.Y(n_1075)
);

BUFx4f_ASAP7_75t_L g1076 ( 
.A(n_893),
.Y(n_1076)
);

OAI21xp33_ASAP7_75t_L g1077 ( 
.A1(n_934),
.A2(n_888),
.B(n_880),
.Y(n_1077)
);

O2A1O1Ixp5_ASAP7_75t_L g1078 ( 
.A1(n_845),
.A2(n_867),
.B(n_865),
.C(n_849),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_799),
.B(n_872),
.Y(n_1079)
);

O2A1O1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_829),
.A2(n_970),
.B(n_971),
.C(n_924),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_R g1081 ( 
.A(n_904),
.B(n_969),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_888),
.A2(n_793),
.B1(n_798),
.B2(n_976),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_799),
.B(n_793),
.Y(n_1083)
);

NOR2xp67_ASAP7_75t_L g1084 ( 
.A(n_967),
.B(n_930),
.Y(n_1084)
);

AOI33xp33_ASAP7_75t_L g1085 ( 
.A1(n_966),
.A2(n_917),
.A3(n_921),
.B1(n_862),
.B2(n_848),
.B3(n_856),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_799),
.B(n_904),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_808),
.A2(n_851),
.B(n_825),
.Y(n_1087)
);

O2A1O1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_920),
.A2(n_899),
.B(n_907),
.C(n_908),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_883),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_SL g1090 ( 
.A1(n_910),
.A2(n_963),
.B(n_842),
.C(n_919),
.Y(n_1090)
);

O2A1O1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_914),
.A2(n_836),
.B(n_949),
.C(n_881),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_822),
.A2(n_818),
.B(n_947),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_887),
.B(n_900),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_832),
.A2(n_933),
.B(n_795),
.C(n_886),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_887),
.B(n_900),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_904),
.B(n_969),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_882),
.A2(n_841),
.B1(n_891),
.B2(n_952),
.Y(n_1097)
);

INVx4_ASAP7_75t_L g1098 ( 
.A(n_904),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_969),
.B(n_835),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_928),
.A2(n_974),
.B1(n_885),
.B2(n_837),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_969),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_874),
.A2(n_950),
.B1(n_861),
.B2(n_972),
.Y(n_1102)
);

OAI22x1_ASAP7_75t_L g1103 ( 
.A1(n_812),
.A2(n_815),
.B1(n_847),
.B2(n_954),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_828),
.A2(n_838),
.B(n_843),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_901),
.B(n_853),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_889),
.B(n_932),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_840),
.B(n_827),
.Y(n_1107)
);

OR2x6_ASAP7_75t_L g1108 ( 
.A(n_975),
.B(n_855),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_936),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_863),
.Y(n_1110)
);

NOR3xp33_ASAP7_75t_SL g1111 ( 
.A(n_946),
.B(n_943),
.C(n_940),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_941),
.B(n_795),
.Y(n_1112)
);

NOR3xp33_ASAP7_75t_L g1113 ( 
.A(n_863),
.B(n_896),
.C(n_846),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_864),
.B(n_873),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_895),
.B(n_879),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_814),
.B(n_906),
.Y(n_1116)
);

AOI33xp33_ASAP7_75t_L g1117 ( 
.A1(n_909),
.A2(n_911),
.A3(n_958),
.B1(n_965),
.B2(n_916),
.B3(n_918),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_905),
.B(n_839),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_839),
.A2(n_925),
.B(n_897),
.C(n_922),
.Y(n_1119)
);

INVx4_ASAP7_75t_L g1120 ( 
.A(n_892),
.Y(n_1120)
);

AND2x2_ASAP7_75t_SL g1121 ( 
.A(n_839),
.B(n_547),
.Y(n_1121)
);

OR2x2_ASAP7_75t_SL g1122 ( 
.A(n_839),
.B(n_389),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_819),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_809),
.A2(n_476),
.B(n_784),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_988),
.A2(n_1119),
.B1(n_997),
.B2(n_1118),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1104),
.A2(n_1087),
.B(n_1124),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1017),
.A2(n_1092),
.B(n_979),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_979),
.A2(n_1107),
.B(n_994),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1003),
.A2(n_1115),
.B(n_1090),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1006),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1002),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_987),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1043),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1024),
.A2(n_1052),
.B(n_1105),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1046),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1116),
.A2(n_998),
.B(n_1088),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1022),
.B(n_1038),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_991),
.B(n_989),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1078),
.A2(n_1091),
.B(n_1074),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_SL g1140 ( 
.A(n_1048),
.B(n_983),
.Y(n_1140)
);

INVx3_ASAP7_75t_SL g1141 ( 
.A(n_993),
.Y(n_1141)
);

OAI22x1_ASAP7_75t_L g1142 ( 
.A1(n_1067),
.A2(n_1053),
.B1(n_1039),
.B2(n_1027),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_986),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1003),
.A2(n_982),
.B(n_1001),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_990),
.B(n_1060),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_991),
.B(n_989),
.Y(n_1146)
);

INVx1_ASAP7_75t_SL g1147 ( 
.A(n_1123),
.Y(n_1147)
);

O2A1O1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_1031),
.A2(n_1062),
.B(n_1042),
.C(n_1051),
.Y(n_1148)
);

OR2x6_ASAP7_75t_L g1149 ( 
.A(n_1040),
.B(n_1060),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_984),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1021),
.B(n_1023),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_982),
.A2(n_1094),
.B(n_995),
.Y(n_1152)
);

AOI221xp5_ASAP7_75t_L g1153 ( 
.A1(n_1042),
.A2(n_1058),
.B1(n_1077),
.B2(n_1061),
.C(n_981),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1058),
.A2(n_1080),
.B(n_1041),
.C(n_1069),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1079),
.A2(n_1020),
.B(n_1097),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_1008),
.B(n_1026),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1023),
.B(n_1005),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_SL g1158 ( 
.A(n_985),
.B(n_1018),
.Y(n_1158)
);

AO31x2_ASAP7_75t_L g1159 ( 
.A1(n_1103),
.A2(n_1082),
.A3(n_1004),
.B(n_1097),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_1014),
.Y(n_1160)
);

AO21x2_ASAP7_75t_L g1161 ( 
.A1(n_1112),
.A2(n_1113),
.B(n_1082),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1010),
.B(n_1121),
.Y(n_1162)
);

OAI21xp33_ASAP7_75t_L g1163 ( 
.A1(n_1072),
.A2(n_1030),
.B(n_1056),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_1096),
.Y(n_1164)
);

INVx1_ASAP7_75t_SL g1165 ( 
.A(n_1055),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_977),
.Y(n_1166)
);

OAI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1075),
.A2(n_1106),
.B(n_1013),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_SL g1168 ( 
.A1(n_1025),
.A2(n_1033),
.B(n_1019),
.C(n_1012),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1070),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1066),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1068),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1063),
.B(n_1007),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1045),
.Y(n_1173)
);

AO31x2_ASAP7_75t_L g1174 ( 
.A1(n_1073),
.A2(n_1025),
.A3(n_1033),
.B(n_996),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1100),
.A2(n_1102),
.B1(n_1083),
.B2(n_1011),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1109),
.A2(n_1015),
.B(n_995),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_996),
.A2(n_1047),
.A3(n_1050),
.B(n_1054),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1016),
.A2(n_1047),
.B(n_1114),
.Y(n_1178)
);

OR2x2_ASAP7_75t_L g1179 ( 
.A(n_1122),
.B(n_1049),
.Y(n_1179)
);

AO31x2_ASAP7_75t_L g1180 ( 
.A1(n_1057),
.A2(n_1044),
.A3(n_1056),
.B(n_1055),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1065),
.Y(n_1181)
);

OA21x2_ASAP7_75t_L g1182 ( 
.A1(n_1111),
.A2(n_1114),
.B(n_1035),
.Y(n_1182)
);

CKINVDCx20_ASAP7_75t_R g1183 ( 
.A(n_1009),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_992),
.B(n_1089),
.Y(n_1184)
);

CKINVDCx11_ASAP7_75t_R g1185 ( 
.A(n_1037),
.Y(n_1185)
);

AO31x2_ASAP7_75t_L g1186 ( 
.A1(n_1093),
.A2(n_1095),
.A3(n_1085),
.B(n_1108),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1108),
.A2(n_999),
.B(n_1099),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1108),
.A2(n_1086),
.B(n_1059),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1040),
.B(n_980),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1034),
.A2(n_1084),
.B(n_1117),
.C(n_1076),
.Y(n_1190)
);

OR2x2_ASAP7_75t_L g1191 ( 
.A(n_1036),
.B(n_1040),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_SL g1192 ( 
.A1(n_1098),
.A2(n_1120),
.B(n_978),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1036),
.A2(n_1120),
.B1(n_1098),
.B2(n_1000),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1081),
.A2(n_977),
.B(n_978),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_977),
.B(n_978),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1000),
.A2(n_1029),
.B1(n_1032),
.B2(n_1064),
.Y(n_1196)
);

OR2x2_ASAP7_75t_L g1197 ( 
.A(n_1064),
.B(n_1101),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1028),
.A2(n_988),
.B(n_997),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1101),
.B(n_1118),
.Y(n_1199)
);

AOI221xp5_ASAP7_75t_L g1200 ( 
.A1(n_997),
.A2(n_988),
.B1(n_871),
.B2(n_870),
.C(n_444),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1104),
.A2(n_1087),
.B(n_847),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1124),
.A2(n_476),
.B(n_784),
.Y(n_1202)
);

CKINVDCx11_ASAP7_75t_R g1203 ( 
.A(n_1009),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1124),
.A2(n_476),
.B(n_784),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_SL g1205 ( 
.A1(n_988),
.A2(n_1119),
.B(n_839),
.C(n_997),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1118),
.B(n_905),
.Y(n_1206)
);

NAND3xp33_ASAP7_75t_L g1207 ( 
.A(n_997),
.B(n_988),
.C(n_1119),
.Y(n_1207)
);

HB1xp67_ASAP7_75t_L g1208 ( 
.A(n_986),
.Y(n_1208)
);

O2A1O1Ixp5_ASAP7_75t_L g1209 ( 
.A1(n_988),
.A2(n_839),
.B(n_1119),
.C(n_925),
.Y(n_1209)
);

OAI221xp5_ASAP7_75t_L g1210 ( 
.A1(n_988),
.A2(n_997),
.B1(n_1119),
.B2(n_870),
.C(n_871),
.Y(n_1210)
);

AO32x2_ASAP7_75t_L g1211 ( 
.A1(n_1042),
.A2(n_996),
.A3(n_1082),
.B1(n_1097),
.B2(n_1020),
.Y(n_1211)
);

AOI221xp5_ASAP7_75t_SL g1212 ( 
.A1(n_997),
.A2(n_988),
.B1(n_1119),
.B2(n_1042),
.C(n_898),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1124),
.A2(n_476),
.B(n_784),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1104),
.A2(n_1087),
.B(n_847),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_977),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1124),
.A2(n_476),
.B(n_784),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_986),
.Y(n_1217)
);

NAND2xp33_ASAP7_75t_L g1218 ( 
.A(n_988),
.B(n_1119),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_988),
.A2(n_997),
.B(n_1119),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1124),
.A2(n_476),
.B(n_784),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_SL g1221 ( 
.A1(n_988),
.A2(n_997),
.B(n_1119),
.Y(n_1221)
);

AO31x2_ASAP7_75t_L g1222 ( 
.A1(n_988),
.A2(n_1094),
.A3(n_1103),
.B(n_1082),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_988),
.A2(n_1119),
.B1(n_997),
.B2(n_839),
.Y(n_1223)
);

NAND3xp33_ASAP7_75t_L g1224 ( 
.A(n_997),
.B(n_988),
.C(n_1119),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1104),
.A2(n_1087),
.B(n_847),
.Y(n_1225)
);

AO32x2_ASAP7_75t_L g1226 ( 
.A1(n_1042),
.A2(n_996),
.A3(n_1082),
.B1(n_1097),
.B2(n_1020),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_986),
.Y(n_1227)
);

O2A1O1Ixp33_ASAP7_75t_SL g1228 ( 
.A1(n_988),
.A2(n_1119),
.B(n_839),
.C(n_997),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1118),
.B(n_905),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_988),
.A2(n_1094),
.A3(n_1103),
.B(n_1082),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1006),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1006),
.Y(n_1232)
);

BUFx8_ASAP7_75t_SL g1233 ( 
.A(n_993),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1104),
.A2(n_1087),
.B(n_847),
.Y(n_1234)
);

AOI221x1_ASAP7_75t_L g1235 ( 
.A1(n_988),
.A2(n_1119),
.B1(n_839),
.B2(n_1042),
.C(n_1073),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_988),
.A2(n_476),
.B1(n_1119),
.B2(n_501),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1124),
.A2(n_476),
.B(n_784),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1118),
.B(n_905),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1104),
.A2(n_1087),
.B(n_847),
.Y(n_1239)
);

INVx4_ASAP7_75t_L g1240 ( 
.A(n_1076),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_988),
.A2(n_1094),
.A3(n_1103),
.B(n_1082),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1104),
.A2(n_1087),
.B(n_847),
.Y(n_1242)
);

AO21x1_ASAP7_75t_L g1243 ( 
.A1(n_997),
.A2(n_839),
.B(n_1058),
.Y(n_1243)
);

O2A1O1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_988),
.A2(n_997),
.B(n_1119),
.C(n_839),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1124),
.A2(n_476),
.B(n_784),
.Y(n_1245)
);

A2O1A1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_997),
.A2(n_988),
.B(n_1119),
.C(n_839),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1104),
.A2(n_1087),
.B(n_847),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1006),
.Y(n_1248)
);

NAND2xp33_ASAP7_75t_L g1249 ( 
.A(n_988),
.B(n_1119),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1118),
.B(n_515),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_997),
.A2(n_988),
.B(n_1119),
.C(n_839),
.Y(n_1251)
);

AO32x1_ASAP7_75t_L g1252 ( 
.A1(n_1042),
.A2(n_1082),
.A3(n_996),
.B1(n_1112),
.B2(n_1110),
.Y(n_1252)
);

INVx1_ASAP7_75t_SL g1253 ( 
.A(n_986),
.Y(n_1253)
);

BUFx4_ASAP7_75t_SL g1254 ( 
.A(n_984),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_977),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_986),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1006),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1006),
.Y(n_1258)
);

O2A1O1Ixp33_ASAP7_75t_SL g1259 ( 
.A1(n_988),
.A2(n_1119),
.B(n_839),
.C(n_997),
.Y(n_1259)
);

AOI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1124),
.A2(n_812),
.B(n_1103),
.Y(n_1260)
);

BUFx2_ASAP7_75t_SL g1261 ( 
.A(n_1071),
.Y(n_1261)
);

CKINVDCx8_ASAP7_75t_R g1262 ( 
.A(n_993),
.Y(n_1262)
);

O2A1O1Ixp5_ASAP7_75t_L g1263 ( 
.A1(n_988),
.A2(n_839),
.B(n_1119),
.C(n_925),
.Y(n_1263)
);

BUFx12f_ASAP7_75t_L g1264 ( 
.A(n_993),
.Y(n_1264)
);

A2O1A1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_997),
.A2(n_988),
.B(n_1119),
.C(n_839),
.Y(n_1265)
);

BUFx8_ASAP7_75t_L g1266 ( 
.A(n_1264),
.Y(n_1266)
);

BUFx4f_ASAP7_75t_SL g1267 ( 
.A(n_1183),
.Y(n_1267)
);

INVx2_ASAP7_75t_SL g1268 ( 
.A(n_1254),
.Y(n_1268)
);

BUFx2_ASAP7_75t_L g1269 ( 
.A(n_1160),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1200),
.A2(n_1210),
.B1(n_1207),
.B2(n_1224),
.Y(n_1270)
);

INVx6_ASAP7_75t_L g1271 ( 
.A(n_1240),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_SL g1272 ( 
.A1(n_1140),
.A2(n_1198),
.B1(n_1207),
.B2(n_1224),
.Y(n_1272)
);

BUFx2_ASAP7_75t_L g1273 ( 
.A(n_1143),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1218),
.A2(n_1249),
.B(n_1221),
.Y(n_1274)
);

BUFx12f_ASAP7_75t_L g1275 ( 
.A(n_1185),
.Y(n_1275)
);

BUFx12f_ASAP7_75t_L g1276 ( 
.A(n_1203),
.Y(n_1276)
);

CKINVDCx6p67_ASAP7_75t_R g1277 ( 
.A(n_1141),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1132),
.Y(n_1278)
);

INVx2_ASAP7_75t_SL g1279 ( 
.A(n_1208),
.Y(n_1279)
);

BUFx2_ASAP7_75t_SL g1280 ( 
.A(n_1240),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_1217),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1206),
.A2(n_1238),
.B1(n_1229),
.B2(n_1137),
.Y(n_1282)
);

CKINVDCx11_ASAP7_75t_R g1283 ( 
.A(n_1262),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1152),
.A2(n_1223),
.B(n_1205),
.Y(n_1284)
);

CKINVDCx11_ASAP7_75t_R g1285 ( 
.A(n_1147),
.Y(n_1285)
);

CKINVDCx6p67_ASAP7_75t_R g1286 ( 
.A(n_1261),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1153),
.A2(n_1125),
.B1(n_1219),
.B2(n_1198),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_SL g1288 ( 
.A1(n_1140),
.A2(n_1125),
.B1(n_1219),
.B2(n_1236),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1130),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_1194),
.Y(n_1290)
);

CKINVDCx6p67_ASAP7_75t_R g1291 ( 
.A(n_1166),
.Y(n_1291)
);

NAND2x1p5_ASAP7_75t_L g1292 ( 
.A(n_1165),
.B(n_1172),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1131),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1227),
.Y(n_1294)
);

BUFx12f_ASAP7_75t_L g1295 ( 
.A(n_1150),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1250),
.B(n_1165),
.Y(n_1296)
);

BUFx12f_ASAP7_75t_L g1297 ( 
.A(n_1179),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1243),
.A2(n_1236),
.B1(n_1142),
.B2(n_1167),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_1233),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1167),
.A2(n_1163),
.B1(n_1139),
.B2(n_1157),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1246),
.A2(n_1265),
.B1(n_1251),
.B2(n_1162),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1231),
.Y(n_1302)
);

OAI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1235),
.A2(n_1158),
.B1(n_1146),
.B2(n_1138),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1147),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1232),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1163),
.A2(n_1139),
.B1(n_1151),
.B2(n_1161),
.Y(n_1306)
);

BUFx4f_ASAP7_75t_SL g1307 ( 
.A(n_1166),
.Y(n_1307)
);

CKINVDCx20_ASAP7_75t_R g1308 ( 
.A(n_1189),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_SL g1309 ( 
.A1(n_1158),
.A2(n_1149),
.B1(n_1178),
.B2(n_1175),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1253),
.Y(n_1310)
);

INVx1_ASAP7_75t_SL g1311 ( 
.A(n_1253),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_SL g1312 ( 
.A1(n_1149),
.A2(n_1178),
.B1(n_1145),
.B2(n_1199),
.Y(n_1312)
);

AOI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1212),
.A2(n_1145),
.B1(n_1228),
.B2(n_1259),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1248),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1209),
.A2(n_1263),
.B(n_1244),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1161),
.A2(n_1129),
.B1(n_1144),
.B2(n_1171),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1256),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1257),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_SL g1319 ( 
.A1(n_1149),
.A2(n_1256),
.B1(n_1184),
.B2(n_1148),
.Y(n_1319)
);

INVx8_ASAP7_75t_L g1320 ( 
.A(n_1166),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_SL g1321 ( 
.A1(n_1212),
.A2(n_1182),
.B1(n_1258),
.B2(n_1135),
.Y(n_1321)
);

CKINVDCx6p67_ASAP7_75t_R g1322 ( 
.A(n_1215),
.Y(n_1322)
);

OAI22x1_ASAP7_75t_L g1323 ( 
.A1(n_1169),
.A2(n_1191),
.B1(n_1196),
.B2(n_1170),
.Y(n_1323)
);

CKINVDCx11_ASAP7_75t_R g1324 ( 
.A(n_1215),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1173),
.A2(n_1181),
.B1(n_1155),
.B2(n_1182),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1187),
.A2(n_1176),
.B1(n_1164),
.B2(n_1156),
.Y(n_1326)
);

AOI21xp33_ASAP7_75t_L g1327 ( 
.A1(n_1154),
.A2(n_1190),
.B(n_1136),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1202),
.A2(n_1220),
.B1(n_1216),
.B2(n_1213),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1188),
.A2(n_1245),
.B1(n_1237),
.B2(n_1204),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1197),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1196),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1193),
.A2(n_1195),
.B1(n_1192),
.B2(n_1128),
.Y(n_1332)
);

INVx6_ASAP7_75t_L g1333 ( 
.A(n_1255),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1186),
.Y(n_1334)
);

OAI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1211),
.A2(n_1226),
.B1(n_1127),
.B2(n_1252),
.Y(n_1335)
);

OAI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1211),
.A2(n_1226),
.B1(n_1252),
.B2(n_1260),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1211),
.A2(n_1226),
.B1(n_1134),
.B2(n_1126),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1247),
.A2(n_1242),
.B1(n_1239),
.B2(n_1225),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1180),
.Y(n_1339)
);

OAI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1174),
.A2(n_1241),
.B1(n_1230),
.B2(n_1222),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1201),
.A2(n_1214),
.B1(n_1234),
.B2(n_1174),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1174),
.A2(n_1177),
.B1(n_1230),
.B2(n_1241),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_1177),
.Y(n_1343)
);

OAI21xp5_ASAP7_75t_SL g1344 ( 
.A1(n_1177),
.A2(n_1159),
.B(n_1168),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1159),
.B(n_1250),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1159),
.A2(n_1200),
.B1(n_1210),
.B2(n_1207),
.Y(n_1346)
);

BUFx3_ASAP7_75t_L g1347 ( 
.A(n_1160),
.Y(n_1347)
);

INVx1_ASAP7_75t_SL g1348 ( 
.A(n_1132),
.Y(n_1348)
);

CKINVDCx11_ASAP7_75t_R g1349 ( 
.A(n_1262),
.Y(n_1349)
);

AOI22x1_ASAP7_75t_SL g1350 ( 
.A1(n_1183),
.A2(n_495),
.B1(n_504),
.B2(n_471),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1250),
.B(n_1118),
.Y(n_1351)
);

CKINVDCx11_ASAP7_75t_R g1352 ( 
.A(n_1262),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1233),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1200),
.A2(n_1210),
.B1(n_1224),
.B2(n_1207),
.Y(n_1354)
);

BUFx12f_ASAP7_75t_L g1355 ( 
.A(n_1185),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_SL g1356 ( 
.A1(n_1140),
.A2(n_983),
.B1(n_1210),
.B2(n_870),
.Y(n_1356)
);

OAI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1210),
.A2(n_988),
.B1(n_997),
.B2(n_1119),
.Y(n_1357)
);

BUFx12f_ASAP7_75t_L g1358 ( 
.A(n_1185),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1160),
.Y(n_1359)
);

BUFx4f_ASAP7_75t_SL g1360 ( 
.A(n_1264),
.Y(n_1360)
);

CKINVDCx11_ASAP7_75t_R g1361 ( 
.A(n_1262),
.Y(n_1361)
);

BUFx12f_ASAP7_75t_L g1362 ( 
.A(n_1185),
.Y(n_1362)
);

BUFx8_ASAP7_75t_SL g1363 ( 
.A(n_1233),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1160),
.Y(n_1364)
);

CKINVDCx14_ASAP7_75t_R g1365 ( 
.A(n_1203),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1200),
.A2(n_1210),
.B1(n_1224),
.B2(n_1207),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1250),
.B(n_1118),
.Y(n_1367)
);

INVx6_ASAP7_75t_L g1368 ( 
.A(n_1240),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1200),
.A2(n_1210),
.B1(n_1224),
.B2(n_1207),
.Y(n_1369)
);

CKINVDCx11_ASAP7_75t_R g1370 ( 
.A(n_1262),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1133),
.Y(n_1371)
);

CKINVDCx6p67_ASAP7_75t_R g1372 ( 
.A(n_1141),
.Y(n_1372)
);

CKINVDCx11_ASAP7_75t_R g1373 ( 
.A(n_1262),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1210),
.B(n_997),
.Y(n_1374)
);

INVx4_ASAP7_75t_L g1375 ( 
.A(n_1240),
.Y(n_1375)
);

INVx5_ASAP7_75t_L g1376 ( 
.A(n_1240),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1200),
.A2(n_1210),
.B1(n_1224),
.B2(n_1207),
.Y(n_1377)
);

NOR2x1_ASAP7_75t_L g1378 ( 
.A(n_1240),
.B(n_1137),
.Y(n_1378)
);

INVx3_ASAP7_75t_L g1379 ( 
.A(n_1240),
.Y(n_1379)
);

CKINVDCx11_ASAP7_75t_R g1380 ( 
.A(n_1262),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1334),
.Y(n_1381)
);

AO21x2_ASAP7_75t_L g1382 ( 
.A1(n_1327),
.A2(n_1315),
.B(n_1357),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1374),
.A2(n_1356),
.B1(n_1287),
.B2(n_1354),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1284),
.A2(n_1341),
.B(n_1329),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1374),
.B(n_1300),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1339),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_L g1387 ( 
.A(n_1301),
.B(n_1272),
.Y(n_1387)
);

INVx3_ASAP7_75t_L g1388 ( 
.A(n_1290),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1341),
.A2(n_1329),
.B(n_1338),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1343),
.Y(n_1390)
);

INVx2_ASAP7_75t_SL g1391 ( 
.A(n_1290),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1282),
.B(n_1351),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1323),
.Y(n_1393)
);

BUFx3_ASAP7_75t_L g1394 ( 
.A(n_1292),
.Y(n_1394)
);

NAND2x1p5_ASAP7_75t_L g1395 ( 
.A(n_1274),
.B(n_1313),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1342),
.B(n_1337),
.Y(n_1396)
);

BUFx12f_ASAP7_75t_L g1397 ( 
.A(n_1283),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_1342),
.B(n_1337),
.Y(n_1398)
);

BUFx3_ASAP7_75t_L g1399 ( 
.A(n_1292),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_L g1400 ( 
.A(n_1345),
.Y(n_1400)
);

INVx3_ASAP7_75t_L g1401 ( 
.A(n_1305),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1340),
.B(n_1344),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1314),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1346),
.B(n_1287),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1338),
.A2(n_1316),
.B(n_1325),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1314),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1316),
.A2(n_1325),
.B(n_1332),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1326),
.A2(n_1298),
.B(n_1346),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1310),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1298),
.B(n_1318),
.Y(n_1410)
);

OAI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1367),
.A2(n_1303),
.B1(n_1304),
.B2(n_1311),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1331),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1289),
.Y(n_1413)
);

AND4x1_ASAP7_75t_L g1414 ( 
.A(n_1270),
.B(n_1369),
.C(n_1377),
.D(n_1366),
.Y(n_1414)
);

OA21x2_ASAP7_75t_L g1415 ( 
.A1(n_1306),
.A2(n_1300),
.B(n_1377),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1340),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1326),
.B(n_1306),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1335),
.B(n_1336),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1336),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1293),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1270),
.B(n_1354),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1302),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1376),
.Y(n_1423)
);

BUFx2_ASAP7_75t_L g1424 ( 
.A(n_1317),
.Y(n_1424)
);

INVx2_ASAP7_75t_SL g1425 ( 
.A(n_1376),
.Y(n_1425)
);

INVx1_ASAP7_75t_SL g1426 ( 
.A(n_1294),
.Y(n_1426)
);

AOI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1288),
.A2(n_1303),
.B1(n_1319),
.B2(n_1309),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1321),
.Y(n_1428)
);

AOI21xp33_ASAP7_75t_L g1429 ( 
.A1(n_1378),
.A2(n_1312),
.B(n_1328),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1296),
.B(n_1371),
.Y(n_1430)
);

INVxp33_ASAP7_75t_L g1431 ( 
.A(n_1285),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_SL g1432 ( 
.A(n_1297),
.B(n_1281),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1330),
.Y(n_1433)
);

CKINVDCx11_ASAP7_75t_R g1434 ( 
.A(n_1349),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1347),
.B(n_1359),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1347),
.B(n_1359),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1269),
.Y(n_1437)
);

INVx2_ASAP7_75t_SL g1438 ( 
.A(n_1271),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1379),
.A2(n_1322),
.B(n_1291),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1279),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1273),
.B(n_1364),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1275),
.A2(n_1355),
.B1(n_1362),
.B2(n_1358),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1278),
.B(n_1308),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1280),
.A2(n_1307),
.B(n_1320),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1348),
.Y(n_1445)
);

INVx5_ASAP7_75t_L g1446 ( 
.A(n_1271),
.Y(n_1446)
);

INVx3_ASAP7_75t_L g1447 ( 
.A(n_1375),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1271),
.B(n_1368),
.Y(n_1448)
);

NAND2xp33_ASAP7_75t_R g1449 ( 
.A(n_1387),
.B(n_1353),
.Y(n_1449)
);

BUFx4f_ASAP7_75t_SL g1450 ( 
.A(n_1397),
.Y(n_1450)
);

INVx11_ASAP7_75t_L g1451 ( 
.A(n_1397),
.Y(n_1451)
);

INVx4_ASAP7_75t_SL g1452 ( 
.A(n_1397),
.Y(n_1452)
);

OA21x2_ASAP7_75t_L g1453 ( 
.A1(n_1405),
.A2(n_1333),
.B(n_1307),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1433),
.B(n_1324),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1392),
.B(n_1267),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1433),
.B(n_1286),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1389),
.A2(n_1368),
.B(n_1320),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1420),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1392),
.B(n_1368),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1435),
.B(n_1277),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1435),
.B(n_1372),
.Y(n_1461)
);

CKINVDCx8_ASAP7_75t_R g1462 ( 
.A(n_1437),
.Y(n_1462)
);

O2A1O1Ixp33_ASAP7_75t_SL g1463 ( 
.A1(n_1387),
.A2(n_1299),
.B(n_1268),
.C(n_1365),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1394),
.B(n_1360),
.Y(n_1464)
);

AOI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1383),
.A2(n_1358),
.B1(n_1275),
.B2(n_1355),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1385),
.B(n_1412),
.Y(n_1466)
);

OA21x2_ASAP7_75t_L g1467 ( 
.A1(n_1405),
.A2(n_1389),
.B(n_1384),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1400),
.B(n_1267),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1400),
.B(n_1362),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1385),
.B(n_1295),
.Y(n_1470)
);

A2O1A1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1427),
.A2(n_1350),
.B(n_1360),
.C(n_1380),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1400),
.B(n_1295),
.Y(n_1472)
);

CKINVDCx20_ASAP7_75t_R g1473 ( 
.A(n_1434),
.Y(n_1473)
);

CKINVDCx6p67_ASAP7_75t_R g1474 ( 
.A(n_1446),
.Y(n_1474)
);

A2O1A1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1427),
.A2(n_1352),
.B(n_1361),
.C(n_1370),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1394),
.B(n_1266),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1422),
.Y(n_1477)
);

AOI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1383),
.A2(n_1276),
.B1(n_1373),
.B2(n_1266),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1436),
.B(n_1276),
.Y(n_1479)
);

NOR2xp33_ASAP7_75t_L g1480 ( 
.A(n_1431),
.B(n_1363),
.Y(n_1480)
);

OAI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1414),
.A2(n_1411),
.B(n_1408),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1400),
.B(n_1441),
.Y(n_1482)
);

AND2x2_ASAP7_75t_SL g1483 ( 
.A(n_1414),
.B(n_1404),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1422),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1430),
.B(n_1400),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1443),
.B(n_1441),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1412),
.B(n_1410),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1399),
.B(n_1409),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1443),
.B(n_1393),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1413),
.Y(n_1490)
);

NAND4xp25_ASAP7_75t_L g1491 ( 
.A(n_1421),
.B(n_1442),
.C(n_1404),
.D(n_1441),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1410),
.B(n_1403),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1413),
.Y(n_1493)
);

AND2x6_ASAP7_75t_L g1494 ( 
.A(n_1410),
.B(n_1417),
.Y(n_1494)
);

INVx1_ASAP7_75t_SL g1495 ( 
.A(n_1426),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1410),
.B(n_1403),
.Y(n_1496)
);

OAI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1411),
.A2(n_1408),
.B(n_1421),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1401),
.B(n_1424),
.Y(n_1498)
);

AND2x6_ASAP7_75t_L g1499 ( 
.A(n_1410),
.B(n_1417),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1381),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1421),
.A2(n_1404),
.B1(n_1395),
.B2(n_1402),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_L g1502 ( 
.A(n_1443),
.B(n_1445),
.Y(n_1502)
);

AO32x2_ASAP7_75t_L g1503 ( 
.A1(n_1391),
.A2(n_1418),
.A3(n_1423),
.B1(n_1425),
.B2(n_1438),
.Y(n_1503)
);

INVx4_ASAP7_75t_L g1504 ( 
.A(n_1446),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1403),
.B(n_1406),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1395),
.A2(n_1402),
.B1(n_1415),
.B2(n_1426),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1393),
.B(n_1437),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_1442),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1458),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1485),
.B(n_1419),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1495),
.B(n_1445),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1490),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1482),
.B(n_1416),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1487),
.B(n_1416),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1486),
.B(n_1382),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1477),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1484),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1487),
.B(n_1418),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1500),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1493),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1492),
.B(n_1496),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1483),
.A2(n_1395),
.B1(n_1417),
.B2(n_1415),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1489),
.B(n_1390),
.Y(n_1523)
);

NAND2x1_ASAP7_75t_L g1524 ( 
.A(n_1504),
.B(n_1388),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1473),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1500),
.Y(n_1526)
);

AND2x4_ASAP7_75t_SL g1527 ( 
.A(n_1474),
.B(n_1388),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1507),
.B(n_1503),
.Y(n_1528)
);

INVxp67_ASAP7_75t_L g1529 ( 
.A(n_1502),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1503),
.B(n_1390),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1492),
.B(n_1396),
.Y(n_1531)
);

AOI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1465),
.A2(n_1478),
.B1(n_1481),
.B2(n_1491),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1496),
.B(n_1396),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1505),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_1455),
.B(n_1432),
.Y(n_1535)
);

NOR2xp67_ASAP7_75t_L g1536 ( 
.A(n_1470),
.B(n_1469),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1505),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1503),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1466),
.Y(n_1539)
);

OR2x6_ASAP7_75t_L g1540 ( 
.A(n_1457),
.B(n_1407),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1506),
.B(n_1396),
.Y(n_1541)
);

BUFx2_ASAP7_75t_L g1542 ( 
.A(n_1488),
.Y(n_1542)
);

INVx5_ASAP7_75t_L g1543 ( 
.A(n_1540),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1528),
.B(n_1542),
.Y(n_1544)
);

INVxp67_ASAP7_75t_L g1545 ( 
.A(n_1511),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1519),
.Y(n_1546)
);

INVx5_ASAP7_75t_SL g1547 ( 
.A(n_1540),
.Y(n_1547)
);

OAI33xp33_ASAP7_75t_L g1548 ( 
.A1(n_1515),
.A2(n_1506),
.A3(n_1501),
.B1(n_1491),
.B2(n_1440),
.B3(n_1459),
.Y(n_1548)
);

INVxp67_ASAP7_75t_L g1549 ( 
.A(n_1539),
.Y(n_1549)
);

INVx5_ASAP7_75t_L g1550 ( 
.A(n_1540),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1529),
.B(n_1498),
.Y(n_1551)
);

NOR2xp33_ASAP7_75t_L g1552 ( 
.A(n_1535),
.B(n_1508),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1528),
.B(n_1453),
.Y(n_1553)
);

AND2x4_ASAP7_75t_L g1554 ( 
.A(n_1530),
.B(n_1488),
.Y(n_1554)
);

INVxp67_ASAP7_75t_SL g1555 ( 
.A(n_1514),
.Y(n_1555)
);

OAI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1532),
.A2(n_1481),
.B1(n_1497),
.B2(n_1478),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_SL g1557 ( 
.A1(n_1522),
.A2(n_1497),
.B1(n_1499),
.B2(n_1494),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1512),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1542),
.B(n_1510),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_SL g1560 ( 
.A1(n_1525),
.A2(n_1465),
.B1(n_1462),
.B2(n_1450),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1530),
.Y(n_1561)
);

BUFx3_ASAP7_75t_L g1562 ( 
.A(n_1524),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1525),
.Y(n_1563)
);

OAI221xp5_ASAP7_75t_L g1564 ( 
.A1(n_1541),
.A2(n_1475),
.B1(n_1471),
.B2(n_1459),
.C(n_1536),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1518),
.B(n_1467),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1526),
.Y(n_1566)
);

OAI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1541),
.A2(n_1415),
.B1(n_1428),
.B2(n_1429),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1523),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1520),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1518),
.B(n_1467),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1531),
.B(n_1398),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1527),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1520),
.Y(n_1573)
);

INVx5_ASAP7_75t_L g1574 ( 
.A(n_1540),
.Y(n_1574)
);

AO21x2_ASAP7_75t_L g1575 ( 
.A1(n_1538),
.A2(n_1381),
.B(n_1386),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1509),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1521),
.B(n_1498),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1538),
.Y(n_1578)
);

AOI21xp33_ASAP7_75t_L g1579 ( 
.A1(n_1514),
.A2(n_1382),
.B(n_1449),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1516),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1555),
.B(n_1534),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1561),
.B(n_1553),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1578),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1544),
.B(n_1521),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1556),
.B(n_1472),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1578),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1565),
.B(n_1570),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1565),
.B(n_1570),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1575),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1575),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1549),
.B(n_1537),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1575),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1569),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1569),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1546),
.B(n_1531),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1558),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1571),
.B(n_1533),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1554),
.B(n_1533),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1573),
.Y(n_1599)
);

INVx1_ASAP7_75t_SL g1600 ( 
.A(n_1571),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1554),
.B(n_1513),
.Y(n_1601)
);

BUFx2_ASAP7_75t_L g1602 ( 
.A(n_1562),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1573),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1558),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1546),
.B(n_1517),
.Y(n_1605)
);

BUFx3_ASAP7_75t_L g1606 ( 
.A(n_1562),
.Y(n_1606)
);

AND2x2_ASAP7_75t_SL g1607 ( 
.A(n_1559),
.B(n_1417),
.Y(n_1607)
);

INVx4_ASAP7_75t_L g1608 ( 
.A(n_1563),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1559),
.B(n_1543),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1605),
.Y(n_1610)
);

OAI221xp5_ASAP7_75t_L g1611 ( 
.A1(n_1585),
.A2(n_1557),
.B1(n_1564),
.B2(n_1560),
.C(n_1579),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1608),
.B(n_1563),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1605),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1593),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1585),
.A2(n_1560),
.B1(n_1567),
.B2(n_1548),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1608),
.B(n_1451),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1593),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1597),
.B(n_1566),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1593),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1597),
.B(n_1566),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1594),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1600),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1597),
.B(n_1568),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1609),
.B(n_1562),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1600),
.B(n_1580),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1594),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1594),
.Y(n_1627)
);

OAI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1607),
.A2(n_1552),
.B(n_1545),
.Y(n_1628)
);

INVxp67_ASAP7_75t_SL g1629 ( 
.A(n_1581),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1599),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1592),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1592),
.Y(n_1632)
);

NAND2x1_ASAP7_75t_L g1633 ( 
.A(n_1602),
.B(n_1576),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1592),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1595),
.B(n_1581),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1592),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1609),
.B(n_1607),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1599),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1606),
.B(n_1543),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1609),
.B(n_1547),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1589),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1589),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1591),
.B(n_1577),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1599),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1607),
.B(n_1547),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1602),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1607),
.B(n_1547),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1603),
.Y(n_1648)
);

NOR2x1_ASAP7_75t_L g1649 ( 
.A(n_1606),
.B(n_1572),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1603),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1601),
.B(n_1547),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1591),
.B(n_1595),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1614),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1615),
.B(n_1629),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1635),
.B(n_1587),
.Y(n_1655)
);

INVxp67_ASAP7_75t_L g1656 ( 
.A(n_1646),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_1637),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1635),
.B(n_1587),
.Y(n_1658)
);

INVx3_ASAP7_75t_L g1659 ( 
.A(n_1633),
.Y(n_1659)
);

BUFx2_ASAP7_75t_L g1660 ( 
.A(n_1649),
.Y(n_1660)
);

CKINVDCx16_ASAP7_75t_R g1661 ( 
.A(n_1612),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1649),
.B(n_1606),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1614),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1637),
.B(n_1606),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1645),
.B(n_1602),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1622),
.B(n_1587),
.Y(n_1666)
);

INVxp67_ASAP7_75t_L g1667 ( 
.A(n_1611),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1628),
.A2(n_1382),
.B1(n_1608),
.B2(n_1547),
.Y(n_1668)
);

NAND2xp33_ASAP7_75t_L g1669 ( 
.A(n_1615),
.B(n_1479),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1645),
.B(n_1647),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1647),
.B(n_1598),
.Y(n_1671)
);

NOR2x1_ASAP7_75t_L g1672 ( 
.A(n_1633),
.B(n_1608),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1617),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1618),
.B(n_1588),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1618),
.B(n_1588),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1617),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1643),
.B(n_1584),
.Y(n_1677)
);

CKINVDCx16_ASAP7_75t_R g1678 ( 
.A(n_1616),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1619),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1619),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1624),
.B(n_1598),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1624),
.B(n_1598),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1652),
.B(n_1584),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1621),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1621),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1620),
.B(n_1588),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1626),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1640),
.B(n_1651),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1667),
.B(n_1610),
.Y(n_1689)
);

OA21x2_ASAP7_75t_L g1690 ( 
.A1(n_1654),
.A2(n_1632),
.B(n_1631),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1659),
.Y(n_1691)
);

INVxp33_ASAP7_75t_L g1692 ( 
.A(n_1672),
.Y(n_1692)
);

OAI211xp5_ASAP7_75t_SL g1693 ( 
.A1(n_1669),
.A2(n_1613),
.B(n_1610),
.C(n_1463),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1688),
.B(n_1640),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1657),
.B(n_1669),
.Y(n_1695)
);

AOI32xp33_ASAP7_75t_L g1696 ( 
.A1(n_1668),
.A2(n_1639),
.A3(n_1651),
.B1(n_1608),
.B2(n_1613),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1656),
.B(n_1601),
.Y(n_1697)
);

OAI21xp33_ASAP7_75t_L g1698 ( 
.A1(n_1688),
.A2(n_1639),
.B(n_1623),
.Y(n_1698)
);

NAND2x1_ASAP7_75t_SL g1699 ( 
.A(n_1662),
.B(n_1659),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1653),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1653),
.Y(n_1701)
);

NAND3xp33_ASAP7_75t_L g1702 ( 
.A(n_1660),
.B(n_1639),
.C(n_1627),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1664),
.B(n_1601),
.Y(n_1703)
);

OAI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1661),
.A2(n_1574),
.B1(n_1550),
.B2(n_1543),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1663),
.Y(n_1705)
);

OA22x2_ASAP7_75t_L g1706 ( 
.A1(n_1660),
.A2(n_1639),
.B1(n_1648),
.B2(n_1644),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1673),
.Y(n_1707)
);

AOI221xp5_ASAP7_75t_SL g1708 ( 
.A1(n_1664),
.A2(n_1665),
.B1(n_1670),
.B2(n_1671),
.C(n_1682),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1678),
.B(n_1480),
.Y(n_1709)
);

NAND2x1p5_ASAP7_75t_L g1710 ( 
.A(n_1662),
.B(n_1446),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1687),
.Y(n_1711)
);

OAI21xp5_ASAP7_75t_L g1712 ( 
.A1(n_1662),
.A2(n_1625),
.B(n_1626),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_1666),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1676),
.Y(n_1714)
);

INVxp67_ASAP7_75t_L g1715 ( 
.A(n_1713),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1713),
.Y(n_1716)
);

AOI222xp33_ASAP7_75t_L g1717 ( 
.A1(n_1695),
.A2(n_1670),
.B1(n_1665),
.B2(n_1671),
.C1(n_1683),
.C2(n_1682),
.Y(n_1717)
);

INVxp67_ASAP7_75t_L g1718 ( 
.A(n_1709),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1699),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1694),
.B(n_1681),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1708),
.B(n_1681),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1700),
.Y(n_1722)
);

AOI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1693),
.A2(n_1666),
.B1(n_1677),
.B2(n_1659),
.Y(n_1723)
);

AOI221xp5_ASAP7_75t_L g1724 ( 
.A1(n_1692),
.A2(n_1679),
.B1(n_1685),
.B2(n_1684),
.C(n_1680),
.Y(n_1724)
);

OAI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1692),
.A2(n_1550),
.B1(n_1543),
.B2(n_1574),
.Y(n_1725)
);

INVxp67_ASAP7_75t_SL g1726 ( 
.A(n_1709),
.Y(n_1726)
);

AOI31xp33_ASAP7_75t_L g1727 ( 
.A1(n_1694),
.A2(n_1658),
.A3(n_1655),
.B(n_1476),
.Y(n_1727)
);

INVxp67_ASAP7_75t_L g1728 ( 
.A(n_1691),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1701),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1697),
.B(n_1655),
.Y(n_1730)
);

O2A1O1Ixp33_ASAP7_75t_L g1731 ( 
.A1(n_1689),
.A2(n_1658),
.B(n_1675),
.C(n_1674),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1705),
.Y(n_1732)
);

AOI22xp33_ASAP7_75t_L g1733 ( 
.A1(n_1698),
.A2(n_1574),
.B1(n_1550),
.B2(n_1543),
.Y(n_1733)
);

OAI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1718),
.A2(n_1702),
.B(n_1706),
.Y(n_1734)
);

O2A1O1Ixp5_ASAP7_75t_L g1735 ( 
.A1(n_1726),
.A2(n_1712),
.B(n_1704),
.C(n_1691),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1718),
.B(n_1703),
.Y(n_1736)
);

AOI21xp33_ASAP7_75t_L g1737 ( 
.A1(n_1731),
.A2(n_1719),
.B(n_1727),
.Y(n_1737)
);

AOI211xp5_ASAP7_75t_SL g1738 ( 
.A1(n_1715),
.A2(n_1714),
.B(n_1711),
.C(n_1707),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1716),
.Y(n_1739)
);

AOI221xp5_ASAP7_75t_L g1740 ( 
.A1(n_1724),
.A2(n_1696),
.B1(n_1706),
.B2(n_1710),
.C(n_1674),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1715),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1728),
.Y(n_1742)
);

INVxp67_ASAP7_75t_SL g1743 ( 
.A(n_1728),
.Y(n_1743)
);

AOI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1721),
.A2(n_1690),
.B(n_1710),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1717),
.A2(n_1690),
.B1(n_1382),
.B2(n_1543),
.Y(n_1745)
);

OAI211xp5_ASAP7_75t_SL g1746 ( 
.A1(n_1740),
.A2(n_1723),
.B(n_1732),
.C(n_1733),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1736),
.B(n_1720),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1743),
.Y(n_1748)
);

AOI31xp33_ASAP7_75t_L g1749 ( 
.A1(n_1737),
.A2(n_1734),
.A3(n_1741),
.B(n_1742),
.Y(n_1749)
);

AOI211xp5_ASAP7_75t_L g1750 ( 
.A1(n_1744),
.A2(n_1725),
.B(n_1730),
.C(n_1729),
.Y(n_1750)
);

NAND3xp33_ASAP7_75t_L g1751 ( 
.A(n_1735),
.B(n_1690),
.C(n_1722),
.Y(n_1751)
);

NOR4xp25_ASAP7_75t_L g1752 ( 
.A(n_1739),
.B(n_1745),
.C(n_1738),
.D(n_1686),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1745),
.B(n_1675),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1736),
.B(n_1452),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1743),
.Y(n_1755)
);

AOI211xp5_ASAP7_75t_L g1756 ( 
.A1(n_1752),
.A2(n_1686),
.B(n_1476),
.C(n_1464),
.Y(n_1756)
);

NAND4xp25_ASAP7_75t_L g1757 ( 
.A(n_1746),
.B(n_1464),
.C(n_1454),
.D(n_1460),
.Y(n_1757)
);

NAND4xp25_ASAP7_75t_L g1758 ( 
.A(n_1750),
.B(n_1461),
.C(n_1452),
.D(n_1468),
.Y(n_1758)
);

NOR4xp75_ASAP7_75t_L g1759 ( 
.A(n_1753),
.B(n_1452),
.C(n_1448),
.D(n_1551),
.Y(n_1759)
);

OAI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1752),
.A2(n_1625),
.B(n_1627),
.Y(n_1760)
);

OAI221xp5_ASAP7_75t_L g1761 ( 
.A1(n_1756),
.A2(n_1749),
.B1(n_1751),
.B2(n_1748),
.C(n_1755),
.Y(n_1761)
);

AOI211xp5_ASAP7_75t_L g1762 ( 
.A1(n_1758),
.A2(n_1747),
.B(n_1754),
.C(n_1641),
.Y(n_1762)
);

OAI211xp5_ASAP7_75t_SL g1763 ( 
.A1(n_1760),
.A2(n_1631),
.B(n_1632),
.C(n_1634),
.Y(n_1763)
);

OAI21xp5_ASAP7_75t_SL g1764 ( 
.A1(n_1757),
.A2(n_1440),
.B(n_1456),
.Y(n_1764)
);

AOI211xp5_ASAP7_75t_L g1765 ( 
.A1(n_1759),
.A2(n_1641),
.B(n_1642),
.C(n_1644),
.Y(n_1765)
);

AOI211xp5_ASAP7_75t_L g1766 ( 
.A1(n_1758),
.A2(n_1642),
.B(n_1648),
.C(n_1650),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1761),
.B(n_1620),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1762),
.Y(n_1768)
);

AOI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1764),
.A2(n_1650),
.B1(n_1638),
.B2(n_1630),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1766),
.B(n_1623),
.Y(n_1770)
);

BUFx2_ASAP7_75t_L g1771 ( 
.A(n_1763),
.Y(n_1771)
);

A2O1A1Ixp33_ASAP7_75t_SL g1772 ( 
.A1(n_1768),
.A2(n_1765),
.B(n_1634),
.C(n_1636),
.Y(n_1772)
);

NOR2x1_ASAP7_75t_L g1773 ( 
.A(n_1771),
.B(n_1638),
.Y(n_1773)
);

NOR2x1_ASAP7_75t_L g1774 ( 
.A(n_1767),
.B(n_1630),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1773),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_SL g1776 ( 
.A1(n_1775),
.A2(n_1770),
.B1(n_1772),
.B2(n_1774),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1776),
.Y(n_1777)
);

OR3x1_ASAP7_75t_L g1778 ( 
.A(n_1776),
.B(n_1769),
.C(n_1590),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1778),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1777),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1780),
.A2(n_1636),
.B1(n_1550),
.B2(n_1574),
.Y(n_1781)
);

AOI22xp5_ASAP7_75t_SL g1782 ( 
.A1(n_1779),
.A2(n_1572),
.B1(n_1438),
.B2(n_1447),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1782),
.Y(n_1783)
);

OAI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1783),
.A2(n_1781),
.B(n_1582),
.Y(n_1784)
);

OAI22xp33_ASAP7_75t_L g1785 ( 
.A1(n_1784),
.A2(n_1596),
.B1(n_1604),
.B2(n_1586),
.Y(n_1785)
);

OAI221xp5_ASAP7_75t_R g1786 ( 
.A1(n_1785),
.A2(n_1574),
.B1(n_1550),
.B2(n_1583),
.C(n_1586),
.Y(n_1786)
);

AOI211xp5_ASAP7_75t_L g1787 ( 
.A1(n_1786),
.A2(n_1444),
.B(n_1439),
.C(n_1448),
.Y(n_1787)
);


endmodule