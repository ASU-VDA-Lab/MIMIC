module fake_jpeg_26099_n_173 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_173);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_25),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVxp33_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_11),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_56),
.Y(n_87)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g81 ( 
.A(n_72),
.Y(n_81)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_0),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_54),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_76),
.B(n_70),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_47),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_77),
.B(n_69),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_78),
.B(n_84),
.Y(n_100)
);

AND2x4_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_57),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_79),
.Y(n_93)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_80),
.Y(n_94)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_83),
.Y(n_104)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_59),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_85),
.B(n_90),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_97),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_84),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_96),
.Y(n_109)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_90),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_101),
.B(n_79),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_73),
.B1(n_49),
.B2(n_59),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_102),
.A2(n_106),
.B1(n_80),
.B2(n_68),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_79),
.A2(n_58),
.B1(n_53),
.B2(n_61),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_110),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_86),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_48),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_114),
.B(n_91),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_75),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_92),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_117),
.B1(n_98),
.B2(n_95),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_106),
.A2(n_58),
.B1(n_50),
.B2(n_65),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_99),
.B1(n_94),
.B2(n_97),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_119),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_125),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_110),
.A2(n_100),
.B1(n_95),
.B2(n_104),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_121),
.A2(n_128),
.B1(n_129),
.B2(n_0),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_122),
.A2(n_124),
.B1(n_113),
.B2(n_54),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_114),
.A2(n_63),
.B(n_64),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_123),
.A2(n_112),
.B(n_1),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_94),
.B1(n_55),
.B2(n_66),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_127),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_51),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_115),
.A2(n_60),
.B1(n_62),
.B2(n_65),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_115),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_136),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_129),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_132),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_20),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_133),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_138),
.B1(n_139),
.B2(n_142),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_56),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_67),
.C(n_16),
.Y(n_137)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_125),
.A2(n_67),
.B1(n_15),
.B2(n_18),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_14),
.Y(n_140)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_127),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_141),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_144),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_122),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_145),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_148),
.A2(n_152),
.B1(n_8),
.B2(n_9),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_135),
.A2(n_138),
.B1(n_142),
.B2(n_143),
.Y(n_150)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_143),
.A2(n_31),
.B1(n_45),
.B2(n_43),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_153),
.Y(n_157)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_157),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_158),
.A2(n_160),
.B1(n_151),
.B2(n_146),
.Y(n_161)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_154),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_161),
.A2(n_159),
.B(n_156),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_150),
.C(n_159),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_147),
.C(n_152),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_165),
.A2(n_162),
.B1(n_155),
.B2(n_32),
.Y(n_166)
);

OAI21x1_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_26),
.B(n_46),
.Y(n_167)
);

AOI221xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_21),
.B1(n_39),
.B2(n_36),
.C(n_34),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_33),
.C(n_30),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_169),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_149),
.C(n_12),
.Y(n_171)
);

BUFx24_ASAP7_75t_SL g172 ( 
.A(n_171),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_149),
.Y(n_173)
);


endmodule