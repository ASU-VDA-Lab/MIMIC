module fake_jpeg_3129_n_418 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_418);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_418;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_4),
.B(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_15),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_60),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_45),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVxp67_ASAP7_75t_SL g54 ( 
.A(n_36),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_19),
.B(n_1),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_55),
.B(n_65),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_19),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_56),
.A2(n_55),
.B1(n_24),
.B2(n_35),
.Y(n_79)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_62),
.B(n_64),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_63),
.Y(n_109)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_66),
.B(n_67),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_23),
.B(n_1),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx5_ASAP7_75t_SL g100 ( 
.A(n_68),
.Y(n_100)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_69),
.A2(n_65),
.B(n_48),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_28),
.B(n_14),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_70),
.B(n_72),
.Y(n_95)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_71),
.A2(n_21),
.B1(n_22),
.B2(n_33),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_28),
.B(n_14),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_23),
.B(n_38),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_38),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_29),
.B(n_12),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_74),
.B(n_27),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_38),
.B1(n_35),
.B2(n_24),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_76),
.A2(n_45),
.B1(n_68),
.B2(n_63),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_78),
.B(n_89),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_79),
.A2(n_85),
.B1(n_102),
.B2(n_108),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_37),
.B1(n_31),
.B2(n_21),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_82),
.A2(n_106),
.B1(n_57),
.B2(n_47),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_73),
.A2(n_24),
.B1(n_35),
.B2(n_29),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_42),
.B(n_37),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_69),
.A2(n_22),
.B1(n_16),
.B2(n_30),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_96),
.A2(n_61),
.B1(n_46),
.B2(n_21),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_37),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_98),
.B(n_102),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_40),
.B(n_21),
.C(n_30),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_105),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_59),
.B(n_27),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_62),
.B(n_20),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_116),
.Y(n_126)
);

INVx4_ASAP7_75t_SL g134 ( 
.A(n_113),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_41),
.A2(n_22),
.B1(n_20),
.B2(n_16),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_52),
.B(n_21),
.C(n_33),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_117),
.Y(n_194)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_118),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

AO22x1_ASAP7_75t_L g120 ( 
.A1(n_76),
.A2(n_91),
.B1(n_103),
.B2(n_82),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_120),
.A2(n_116),
.B(n_80),
.Y(n_168)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_98),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_127),
.Y(n_164)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_84),
.B(n_53),
.Y(n_127)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_128),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_129),
.A2(n_50),
.B1(n_39),
.B2(n_43),
.Y(n_181)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_132),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_109),
.B1(n_130),
.B2(n_144),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_93),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_156),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

INVx13_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_138),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_112),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_143),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_141),
.A2(n_150),
.B1(n_100),
.B2(n_21),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_142),
.B(n_154),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_81),
.B(n_51),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_103),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_144),
.B(n_146),
.Y(n_191)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_103),
.Y(n_146)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_147),
.Y(n_195)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_107),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_149),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_78),
.A2(n_66),
.B1(n_71),
.B2(n_53),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_82),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_151),
.Y(n_185)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

OR2x2_ASAP7_75t_SL g153 ( 
.A(n_99),
.B(n_51),
.Y(n_153)
);

NAND3xp33_ASAP7_75t_SL g197 ( 
.A(n_153),
.B(n_134),
.C(n_146),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_86),
.B(n_49),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_75),
.Y(n_155)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_80),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_158),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_82),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_159),
.A2(n_171),
.B1(n_178),
.B2(n_183),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_124),
.B(n_114),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_179),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_197),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_151),
.A2(n_75),
.B1(n_88),
.B2(n_90),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_126),
.A2(n_88),
.B(n_93),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_175),
.A2(n_181),
.B(n_190),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_123),
.A2(n_77),
.B1(n_92),
.B2(n_90),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_124),
.B(n_133),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_142),
.A2(n_92),
.B1(n_77),
.B2(n_100),
.Y(n_183)
);

XNOR2x1_ASAP7_75t_L g186 ( 
.A(n_120),
.B(n_94),
.Y(n_186)
);

NOR2x1_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_129),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_121),
.B(n_94),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_188),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_1),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_190),
.A2(n_135),
.B1(n_136),
.B2(n_139),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_120),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_192),
.A2(n_132),
.B1(n_117),
.B2(n_122),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_161),
.A2(n_139),
.B(n_134),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_198),
.A2(n_210),
.B(n_216),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_125),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_199),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_201),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_157),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_203),
.B(n_211),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_118),
.C(n_150),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_204),
.B(n_235),
.C(n_182),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_177),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_205),
.B(n_215),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_206),
.A2(n_225),
.B1(n_230),
.B2(n_2),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_208),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_155),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_209),
.B(n_219),
.Y(n_257)
);

OA21x2_ASAP7_75t_L g210 ( 
.A1(n_161),
.A2(n_129),
.B(n_145),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_119),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_213),
.A2(n_228),
.B1(n_192),
.B2(n_173),
.Y(n_236)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_162),
.Y(n_214)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_177),
.Y(n_215)
);

BUFx8_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

BUFx5_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_163),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_218),
.B(n_220),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_131),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_179),
.B(n_138),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_168),
.B(n_129),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_221),
.A2(n_222),
.B(n_176),
.Y(n_243)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_162),
.Y(n_223)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_223),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_152),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_224),
.B(n_227),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_196),
.A2(n_148),
.B1(n_128),
.B2(n_147),
.Y(n_225)
);

BUFx12_ASAP7_75t_L g226 ( 
.A(n_184),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_226),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_163),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_196),
.A2(n_137),
.B1(n_3),
.B2(n_5),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_160),
.Y(n_229)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_167),
.A2(n_183),
.B1(n_159),
.B2(n_188),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_178),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_169),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_175),
.B(n_137),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_232),
.Y(n_270)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_160),
.Y(n_233)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_180),
.Y(n_234)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_167),
.B(n_137),
.C(n_5),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_236),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_221),
.A2(n_191),
.B1(n_171),
.B2(n_186),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_237),
.A2(n_242),
.B(n_243),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_221),
.A2(n_189),
.B1(n_195),
.B2(n_194),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_268),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_212),
.A2(n_172),
.B1(n_176),
.B2(n_193),
.Y(n_242)
);

OA21x2_ASAP7_75t_L g245 ( 
.A1(n_198),
.A2(n_193),
.B(n_172),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_245),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_200),
.B(n_182),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_247),
.B(n_204),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_212),
.Y(n_278)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_258),
.Y(n_282)
);

AOI32xp33_ASAP7_75t_L g259 ( 
.A1(n_205),
.A2(n_195),
.A3(n_169),
.B1(n_166),
.B2(n_194),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_264),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_210),
.A2(n_189),
.B1(n_166),
.B2(n_170),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_261),
.A2(n_206),
.B1(n_202),
.B2(n_231),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_216),
.A2(n_170),
.B(n_5),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_262),
.A2(n_217),
.B(n_213),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_263),
.A2(n_269),
.B1(n_217),
.B2(n_208),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_209),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_214),
.Y(n_266)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_266),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_200),
.B(n_6),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_201),
.C(n_235),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_219),
.B(n_6),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_230),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_272),
.A2(n_287),
.B1(n_270),
.B2(n_245),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_218),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_276),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_227),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_248),
.C(n_254),
.Y(n_303)
);

OAI21xp33_ASAP7_75t_L g279 ( 
.A1(n_240),
.A2(n_212),
.B(n_207),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_279),
.B(n_280),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_281),
.B(n_247),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_246),
.B(n_223),
.Y(n_283)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_283),
.Y(n_313)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_239),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_284),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_240),
.B(n_229),
.Y(n_285)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_285),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_237),
.A2(n_202),
.B1(n_222),
.B2(n_210),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_253),
.B(n_207),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_288),
.B(n_290),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_241),
.A2(n_215),
.B(n_225),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_289),
.A2(n_291),
.B(n_245),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_256),
.B(n_228),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_241),
.A2(n_243),
.B(n_270),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_258),
.Y(n_292)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_292),
.Y(n_322)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_239),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_294),
.A2(n_295),
.B1(n_297),
.B2(n_298),
.Y(n_309)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_250),
.Y(n_295)
);

NAND2x1_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_238),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_265),
.B(n_233),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_257),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_299),
.A2(n_236),
.B1(n_261),
.B2(n_242),
.Y(n_307)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_250),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_300),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_302),
.A2(n_324),
.B1(n_325),
.B2(n_296),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_303),
.B(n_317),
.C(n_291),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_304),
.B(n_312),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_285),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_306),
.B(n_288),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_314),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_293),
.A2(n_264),
.B1(n_262),
.B2(n_254),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_308),
.A2(n_316),
.B1(n_319),
.B2(n_321),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_310),
.A2(n_314),
.B(n_325),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_278),
.B(n_267),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_281),
.B(n_268),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_315),
.B(n_274),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_293),
.A2(n_298),
.B1(n_275),
.B2(n_271),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_280),
.B(n_266),
.C(n_251),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_275),
.A2(n_251),
.B1(n_252),
.B2(n_255),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_275),
.A2(n_252),
.B1(n_255),
.B2(n_260),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_287),
.A2(n_249),
.B1(n_260),
.B2(n_234),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_271),
.A2(n_249),
.B1(n_217),
.B2(n_244),
.Y(n_325)
);

OA22x2_ASAP7_75t_L g326 ( 
.A1(n_282),
.A2(n_244),
.B1(n_226),
.B2(n_8),
.Y(n_326)
);

OA21x2_ASAP7_75t_L g340 ( 
.A1(n_326),
.A2(n_272),
.B(n_295),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_327),
.B(n_343),
.Y(n_356)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_318),
.Y(n_329)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_329),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_277),
.C(n_289),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_330),
.B(n_335),
.C(n_342),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_L g331 ( 
.A1(n_313),
.A2(n_273),
.B1(n_283),
.B2(n_297),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_331),
.A2(n_340),
.B1(n_346),
.B2(n_323),
.Y(n_357)
);

NAND3xp33_ASAP7_75t_L g358 ( 
.A(n_332),
.B(n_339),
.C(n_311),
.Y(n_358)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_305),
.Y(n_334)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_334),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_317),
.B(n_277),
.C(n_276),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_337),
.Y(n_360)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_309),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_338),
.B(n_341),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_320),
.B(n_290),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_322),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_312),
.B(n_292),
.C(n_282),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_301),
.B(n_274),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_344),
.B(n_304),
.Y(n_349)
);

FAx1_ASAP7_75t_SL g345 ( 
.A(n_310),
.B(n_300),
.CI(n_294),
.CON(n_345),
.SN(n_345)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_345),
.B(n_347),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_316),
.A2(n_286),
.B1(n_284),
.B2(n_226),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_311),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_348),
.A2(n_302),
.B(n_324),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_349),
.B(n_333),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_327),
.B(n_286),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_351),
.B(n_353),
.Y(n_367)
);

BUFx12_ASAP7_75t_L g352 ( 
.A(n_345),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_352),
.Y(n_368)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_336),
.Y(n_353)
);

XNOR2x1_ASAP7_75t_L g373 ( 
.A(n_355),
.B(n_336),
.Y(n_373)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_357),
.Y(n_369)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_358),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_333),
.B(n_315),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_361),
.B(n_365),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_346),
.Y(n_363)
);

AO22x1_ASAP7_75t_L g379 ( 
.A1(n_363),
.A2(n_328),
.B1(n_307),
.B2(n_345),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_343),
.B(n_308),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_366),
.B(n_354),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_356),
.B(n_335),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_370),
.B(n_378),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_356),
.B(n_330),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_372),
.B(n_374),
.Y(n_380)
);

MAJx2_ASAP7_75t_L g387 ( 
.A(n_373),
.B(n_340),
.C(n_352),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_364),
.B(n_342),
.C(n_344),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_364),
.B(n_328),
.C(n_321),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_376),
.B(n_377),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_361),
.B(n_328),
.C(n_319),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_349),
.B(n_360),
.C(n_365),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_379),
.A2(n_368),
.B1(n_363),
.B2(n_360),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_382),
.Y(n_396)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_383),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_375),
.B(n_362),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_384),
.B(n_385),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_370),
.B(n_359),
.C(n_340),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_367),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_386),
.B(n_391),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_387),
.B(n_379),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_376),
.A2(n_352),
.B(n_350),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_388),
.A2(n_389),
.B(n_377),
.Y(n_395)
);

NAND2x1p5_ASAP7_75t_L g389 ( 
.A(n_373),
.B(n_347),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_371),
.B(n_326),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_380),
.A2(n_381),
.B(n_369),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_393),
.A2(n_395),
.B(n_401),
.Y(n_405)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_397),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_390),
.B(n_374),
.C(n_366),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_398),
.B(n_385),
.Y(n_407)
);

OAI22xp33_ASAP7_75t_L g399 ( 
.A1(n_387),
.A2(n_326),
.B1(n_7),
.B2(n_9),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_399),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_391),
.A2(n_326),
.B(n_7),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_394),
.B(n_400),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_402),
.A2(n_6),
.B(n_10),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_392),
.B(n_382),
.Y(n_403)
);

INVxp33_ASAP7_75t_L g409 ( 
.A(n_403),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_407),
.B(n_408),
.Y(n_411)
);

MAJx2_ASAP7_75t_L g408 ( 
.A(n_396),
.B(n_389),
.C(n_9),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_405),
.A2(n_396),
.B(n_399),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_410),
.A2(n_404),
.B(n_402),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_412),
.A2(n_406),
.B1(n_10),
.B2(n_11),
.Y(n_414)
);

NOR3xp33_ASAP7_75t_L g415 ( 
.A(n_413),
.B(n_414),
.C(n_411),
.Y(n_415)
);

OA21x2_ASAP7_75t_L g416 ( 
.A1(n_415),
.A2(n_409),
.B(n_10),
.Y(n_416)
);

AOI21x1_ASAP7_75t_L g417 ( 
.A1(n_416),
.A2(n_11),
.B(n_273),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_417),
.B(n_11),
.Y(n_418)
);


endmodule