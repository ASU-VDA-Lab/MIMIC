module fake_aes_1226_n_1325 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_272, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_270, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_1325);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_272;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
output n_1325;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1079;
wire n_315;
wire n_409;
wire n_295;
wire n_1321;
wire n_677;
wire n_1242;
wire n_283;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_281;
wire n_487;
wire n_451;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_280;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_275;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_287;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_286;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_282;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_285;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_288;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_276;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_405;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g275 ( .A(n_126), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_9), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_140), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_19), .Y(n_278) );
BUFx3_ASAP7_75t_L g279 ( .A(n_175), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_128), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_189), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_162), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_34), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_78), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_231), .Y(n_285) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_21), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g287 ( .A(n_72), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_15), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_206), .Y(n_289) );
INVxp67_ASAP7_75t_SL g290 ( .A(n_44), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_122), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_236), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_75), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_91), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_55), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_184), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_84), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_130), .Y(n_298) );
INVxp67_ASAP7_75t_SL g299 ( .A(n_104), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_67), .Y(n_300) );
CKINVDCx20_ASAP7_75t_R g301 ( .A(n_183), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_235), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_202), .Y(n_303) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_35), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_147), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_174), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_81), .Y(n_307) );
CKINVDCx20_ASAP7_75t_R g308 ( .A(n_237), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_27), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_109), .Y(n_310) );
CKINVDCx16_ASAP7_75t_R g311 ( .A(n_196), .Y(n_311) );
INVxp33_ASAP7_75t_SL g312 ( .A(n_120), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_254), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_43), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_114), .Y(n_315) );
CKINVDCx20_ASAP7_75t_R g316 ( .A(n_227), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_192), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_219), .Y(n_318) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_65), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_40), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_226), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_273), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_150), .Y(n_323) );
NOR2xp67_ASAP7_75t_L g324 ( .A(n_33), .B(n_137), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_46), .Y(n_325) );
INVxp67_ASAP7_75t_L g326 ( .A(n_180), .Y(n_326) );
INVxp67_ASAP7_75t_SL g327 ( .A(n_95), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_1), .Y(n_328) );
INVxp33_ASAP7_75t_SL g329 ( .A(n_272), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_68), .Y(n_330) );
CKINVDCx20_ASAP7_75t_R g331 ( .A(n_63), .Y(n_331) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_212), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_124), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_25), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_145), .Y(n_335) );
CKINVDCx14_ASAP7_75t_R g336 ( .A(n_56), .Y(n_336) );
INVxp33_ASAP7_75t_SL g337 ( .A(n_188), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_48), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_61), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_34), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_53), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_198), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_129), .Y(n_343) );
INVxp67_ASAP7_75t_SL g344 ( .A(n_4), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_83), .Y(n_345) );
INVxp33_ASAP7_75t_L g346 ( .A(n_131), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_148), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_70), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_271), .Y(n_349) );
INVxp67_ASAP7_75t_L g350 ( .A(n_40), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_65), .Y(n_351) );
BUFx3_ASAP7_75t_L g352 ( .A(n_89), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_252), .Y(n_353) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_105), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_135), .Y(n_355) );
BUFx3_ASAP7_75t_L g356 ( .A(n_117), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_247), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_144), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_166), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_45), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_30), .Y(n_361) );
CKINVDCx16_ASAP7_75t_R g362 ( .A(n_18), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_76), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_268), .Y(n_364) );
INVx1_ASAP7_75t_SL g365 ( .A(n_172), .Y(n_365) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_197), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_8), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_178), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_204), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_77), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_88), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_82), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_136), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_35), .Y(n_374) );
INVx3_ASAP7_75t_L g375 ( .A(n_79), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_171), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_241), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_238), .Y(n_378) );
INVxp33_ASAP7_75t_L g379 ( .A(n_127), .Y(n_379) );
CKINVDCx20_ASAP7_75t_R g380 ( .A(n_10), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_228), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_23), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_222), .Y(n_383) );
INVx1_ASAP7_75t_SL g384 ( .A(n_11), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_107), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_99), .Y(n_386) );
BUFx5_ASAP7_75t_L g387 ( .A(n_133), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_4), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_232), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_94), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_260), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_90), .Y(n_392) );
CKINVDCx20_ASAP7_75t_R g393 ( .A(n_165), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_208), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_52), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_80), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_6), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_20), .Y(n_398) );
INVxp33_ASAP7_75t_L g399 ( .A(n_158), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_199), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_60), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_125), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_154), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_57), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_161), .Y(n_405) );
CKINVDCx16_ASAP7_75t_R g406 ( .A(n_121), .Y(n_406) );
INVxp33_ASAP7_75t_SL g407 ( .A(n_46), .Y(n_407) );
CKINVDCx20_ASAP7_75t_R g408 ( .A(n_92), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_101), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_214), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_38), .Y(n_411) );
INVxp33_ASAP7_75t_SL g412 ( .A(n_53), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_152), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_300), .Y(n_414) );
INVx3_ASAP7_75t_L g415 ( .A(n_375), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_346), .B(n_0), .Y(n_416) );
AND2x4_ASAP7_75t_SL g417 ( .A(n_287), .B(n_71), .Y(n_417) );
INVxp67_ASAP7_75t_L g418 ( .A(n_353), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_300), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_325), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_375), .B(n_387), .Y(n_421) );
NOR2x1_ASAP7_75t_L g422 ( .A(n_375), .B(n_0), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_346), .B(n_1), .Y(n_423) );
BUFx2_ASAP7_75t_L g424 ( .A(n_336), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_325), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_387), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_351), .Y(n_427) );
HAxp5_ASAP7_75t_SL g428 ( .A(n_278), .B(n_2), .CON(n_428), .SN(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_379), .B(n_2), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_351), .Y(n_430) );
CKINVDCx5p33_ASAP7_75t_R g431 ( .A(n_311), .Y(n_431) );
BUFx2_ASAP7_75t_L g432 ( .A(n_336), .Y(n_432) );
OAI21x1_ASAP7_75t_L g433 ( .A1(n_292), .A2(n_74), .B(n_73), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_362), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_387), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_286), .Y(n_436) );
INVx6_ASAP7_75t_L g437 ( .A(n_387), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_387), .Y(n_438) );
INVx6_ASAP7_75t_L g439 ( .A(n_387), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_407), .A2(n_3), .B1(n_5), .B2(n_6), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_407), .A2(n_3), .B1(n_5), .B2(n_7), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_404), .Y(n_442) );
AND2x4_ASAP7_75t_L g443 ( .A(n_404), .B(n_7), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_379), .B(n_8), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_283), .B(n_9), .Y(n_445) );
NOR2xp33_ASAP7_75t_SL g446 ( .A(n_406), .B(n_274), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_331), .Y(n_447) );
BUFx2_ASAP7_75t_L g448 ( .A(n_424), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_424), .B(n_399), .Y(n_449) );
INVx4_ASAP7_75t_L g450 ( .A(n_437), .Y(n_450) );
INVx4_ASAP7_75t_SL g451 ( .A(n_437), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_426), .Y(n_452) );
INVx3_ASAP7_75t_L g453 ( .A(n_415), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_431), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_432), .B(n_399), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_426), .Y(n_456) );
INVx4_ASAP7_75t_L g457 ( .A(n_437), .Y(n_457) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_440), .A2(n_380), .B1(n_331), .B2(n_412), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_426), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_432), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_418), .B(n_326), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_435), .Y(n_462) );
NAND2xp33_ASAP7_75t_L g463 ( .A(n_423), .B(n_387), .Y(n_463) );
INVx4_ASAP7_75t_L g464 ( .A(n_437), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_418), .B(n_304), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_423), .B(n_294), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_435), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_435), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_415), .B(n_292), .Y(n_469) );
CKINVDCx16_ASAP7_75t_R g470 ( .A(n_434), .Y(n_470) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_433), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_438), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_415), .B(n_276), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_415), .B(n_307), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_438), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_438), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_437), .Y(n_477) );
INVx1_ASAP7_75t_SL g478 ( .A(n_417), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_439), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_436), .B(n_312), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_439), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_423), .B(n_307), .Y(n_482) );
INVx1_ASAP7_75t_SL g483 ( .A(n_417), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_439), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_436), .B(n_319), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_429), .B(n_310), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_429), .B(n_276), .Y(n_487) );
NAND2xp33_ASAP7_75t_R g488 ( .A(n_429), .B(n_412), .Y(n_488) );
BUFx10_ASAP7_75t_L g489 ( .A(n_439), .Y(n_489) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_433), .Y(n_490) );
AND2x2_ASAP7_75t_SL g491 ( .A(n_417), .B(n_310), .Y(n_491) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_433), .Y(n_492) );
INVx3_ASAP7_75t_L g493 ( .A(n_443), .Y(n_493) );
AND2x4_ASAP7_75t_L g494 ( .A(n_422), .B(n_288), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_453), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_453), .Y(n_496) );
BUFx3_ASAP7_75t_L g497 ( .A(n_489), .Y(n_497) );
BUFx2_ASAP7_75t_L g498 ( .A(n_448), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_453), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_453), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_493), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_480), .A2(n_444), .B1(n_416), .B2(n_446), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_493), .Y(n_503) );
INVx4_ASAP7_75t_L g504 ( .A(n_489), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_468), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_493), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_494), .A2(n_443), .B1(n_439), .B2(n_416), .Y(n_507) );
INVx3_ASAP7_75t_SL g508 ( .A(n_491), .Y(n_508) );
INVx1_ASAP7_75t_SL g509 ( .A(n_460), .Y(n_509) );
INVx3_ASAP7_75t_L g510 ( .A(n_493), .Y(n_510) );
BUFx3_ASAP7_75t_L g511 ( .A(n_489), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_485), .B(n_444), .Y(n_512) );
AND2x4_ASAP7_75t_L g513 ( .A(n_494), .B(n_443), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_482), .B(n_443), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_482), .B(n_422), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_486), .B(n_294), .Y(n_516) );
NAND2x1p5_ASAP7_75t_L g517 ( .A(n_491), .B(n_440), .Y(n_517) );
OR2x2_ASAP7_75t_SL g518 ( .A(n_470), .B(n_428), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_469), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_468), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_468), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_448), .Y(n_522) );
OAI22xp5_ASAP7_75t_SL g523 ( .A1(n_458), .A2(n_447), .B1(n_380), .B2(n_441), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_494), .B(n_446), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_460), .B(n_295), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_472), .Y(n_526) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_489), .Y(n_527) );
INVx3_ASAP7_75t_L g528 ( .A(n_494), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_472), .Y(n_529) );
INVxp67_ASAP7_75t_SL g530 ( .A(n_486), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_463), .A2(n_490), .B1(n_492), .B2(n_471), .Y(n_531) );
NAND2x1p5_ASAP7_75t_L g532 ( .A(n_491), .B(n_441), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_469), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_471), .B(n_275), .Y(n_534) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_487), .Y(n_535) );
BUFx2_ASAP7_75t_L g536 ( .A(n_487), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_449), .B(n_297), .Y(n_537) );
NOR2xp33_ASAP7_75t_SL g538 ( .A(n_478), .B(n_287), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_488), .A2(n_308), .B1(n_316), .B2(n_301), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_449), .B(n_297), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_474), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_470), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_471), .B(n_277), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_455), .B(n_295), .Y(n_544) );
NAND2x1p5_ASAP7_75t_L g545 ( .A(n_478), .B(n_309), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_472), .Y(n_546) );
INVxp67_ASAP7_75t_L g547 ( .A(n_485), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_476), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_455), .B(n_317), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_461), .B(n_317), .Y(n_550) );
AND2x4_ASAP7_75t_L g551 ( .A(n_473), .B(n_445), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_471), .B(n_280), .Y(n_552) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_465), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_465), .B(n_343), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_466), .B(n_343), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_474), .B(n_349), .Y(n_556) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_471), .Y(n_557) );
OR2x2_ASAP7_75t_SL g558 ( .A(n_458), .B(n_428), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_452), .Y(n_559) );
BUFx2_ASAP7_75t_L g560 ( .A(n_483), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_452), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_456), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_483), .B(n_349), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_454), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_456), .B(n_355), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_459), .Y(n_566) );
NAND3xp33_ASAP7_75t_SL g567 ( .A(n_459), .B(n_308), .C(n_301), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_462), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_471), .B(n_281), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_462), .B(n_355), .Y(n_570) );
AOI22xp5_ASAP7_75t_L g571 ( .A1(n_467), .A2(n_332), .B1(n_393), .B2(n_316), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_490), .B(n_284), .Y(n_572) );
INVx3_ASAP7_75t_L g573 ( .A(n_490), .Y(n_573) );
INVx2_ASAP7_75t_SL g574 ( .A(n_492), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_467), .B(n_445), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_475), .B(n_366), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_490), .B(n_285), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_475), .B(n_366), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_450), .B(n_376), .Y(n_579) );
BUFx12f_ASAP7_75t_L g580 ( .A(n_490), .Y(n_580) );
INVxp67_ASAP7_75t_SL g581 ( .A(n_450), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_490), .A2(n_419), .B1(n_420), .B2(n_414), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_450), .B(n_376), .Y(n_583) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_492), .Y(n_584) );
INVxp67_ASAP7_75t_L g585 ( .A(n_476), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_492), .A2(n_419), .B1(n_420), .B2(n_414), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_450), .B(n_377), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_509), .A2(n_332), .B1(n_408), .B2(n_393), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_510), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_510), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_530), .Y(n_591) );
O2A1O1Ixp33_ASAP7_75t_L g592 ( .A1(n_547), .A2(n_350), .B(n_421), .C(n_344), .Y(n_592) );
BUFx6f_ASAP7_75t_L g593 ( .A(n_527), .Y(n_593) );
AND2x4_ASAP7_75t_L g594 ( .A(n_528), .B(n_513), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_505), .Y(n_595) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_527), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_553), .B(n_312), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_512), .B(n_329), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_575), .A2(n_408), .B1(n_337), .B2(n_329), .Y(n_599) );
CKINVDCx5p33_ASAP7_75t_R g600 ( .A(n_564), .Y(n_600) );
INVx2_ASAP7_75t_SL g601 ( .A(n_560), .Y(n_601) );
AND2x4_ASAP7_75t_L g602 ( .A(n_528), .B(n_290), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_545), .B(n_457), .Y(n_603) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_527), .Y(n_604) );
BUFx4f_ASAP7_75t_L g605 ( .A(n_508), .Y(n_605) );
OAI22xp5_ASAP7_75t_SL g606 ( .A1(n_518), .A2(n_428), .B1(n_361), .B2(n_337), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_507), .A2(n_492), .B1(n_361), .B2(n_378), .Y(n_607) );
BUFx4f_ASAP7_75t_L g608 ( .A(n_508), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_535), .B(n_457), .Y(n_609) );
CKINVDCx6p67_ASAP7_75t_R g610 ( .A(n_564), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_544), .B(n_457), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_519), .Y(n_612) );
AOI22xp33_ASAP7_75t_SL g613 ( .A1(n_538), .A2(n_330), .B1(n_382), .B2(n_340), .Y(n_613) );
A2O1A1Ixp33_ASAP7_75t_L g614 ( .A1(n_533), .A2(n_476), .B(n_492), .C(n_320), .Y(n_614) );
BUFx2_ASAP7_75t_L g615 ( .A(n_522), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_536), .B(n_457), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_541), .Y(n_617) );
AOI21xp5_ASAP7_75t_L g618 ( .A1(n_534), .A2(n_464), .B(n_477), .Y(n_618) );
O2A1O1Ixp33_ASAP7_75t_L g619 ( .A1(n_524), .A2(n_328), .B(n_334), .C(n_314), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_551), .B(n_464), .Y(n_620) );
A2O1A1Ixp33_ASAP7_75t_L g621 ( .A1(n_515), .A2(n_338), .B(n_341), .C(n_339), .Y(n_621) );
AOI21xp5_ASAP7_75t_L g622 ( .A1(n_534), .A2(n_552), .B(n_543), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_505), .Y(n_623) );
CKINVDCx8_ASAP7_75t_R g624 ( .A(n_542), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_554), .B(n_384), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_516), .B(n_378), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_520), .Y(n_627) );
BUFx2_ASAP7_75t_L g628 ( .A(n_522), .Y(n_628) );
O2A1O1Ixp33_ASAP7_75t_SL g629 ( .A1(n_543), .A2(n_484), .B(n_477), .C(n_291), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_504), .B(n_451), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_537), .B(n_484), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_520), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_501), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g634 ( .A1(n_552), .A2(n_481), .B(n_479), .Y(n_634) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_527), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_503), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_507), .A2(n_360), .B1(n_367), .B2(n_348), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_521), .Y(n_638) );
BUFx6f_ASAP7_75t_L g639 ( .A(n_497), .Y(n_639) );
INVxp67_ASAP7_75t_SL g640 ( .A(n_571), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_513), .A2(n_388), .B1(n_395), .B2(n_374), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_521), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_506), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_502), .A2(n_398), .B1(n_401), .B2(n_397), .Y(n_644) );
INVx4_ASAP7_75t_L g645 ( .A(n_504), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g646 ( .A(n_504), .B(n_451), .Y(n_646) );
INVx1_ASAP7_75t_SL g647 ( .A(n_498), .Y(n_647) );
BUFx3_ASAP7_75t_L g648 ( .A(n_542), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_513), .Y(n_649) );
OR2x6_ASAP7_75t_L g650 ( .A(n_517), .B(n_411), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_517), .A2(n_327), .B1(n_299), .B2(n_425), .Y(n_651) );
O2A1O1Ixp33_ASAP7_75t_L g652 ( .A1(n_514), .A2(n_540), .B(n_549), .C(n_567), .Y(n_652) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_525), .Y(n_653) );
A2O1A1Ixp33_ASAP7_75t_L g654 ( .A1(n_559), .A2(n_324), .B(n_427), .C(n_425), .Y(n_654) );
BUFx6f_ASAP7_75t_L g655 ( .A(n_497), .Y(n_655) );
INVx1_ASAP7_75t_SL g656 ( .A(n_539), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_561), .Y(n_657) );
INVx3_ASAP7_75t_L g658 ( .A(n_580), .Y(n_658) );
AND2x6_ASAP7_75t_L g659 ( .A(n_511), .B(n_279), .Y(n_659) );
INVx3_ASAP7_75t_L g660 ( .A(n_580), .Y(n_660) );
BUFx6f_ASAP7_75t_L g661 ( .A(n_511), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_562), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_569), .A2(n_481), .B(n_479), .Y(n_663) );
AOI222xp33_ASAP7_75t_L g664 ( .A1(n_523), .A2(n_427), .B1(n_430), .B2(n_442), .C1(n_293), .C2(n_289), .Y(n_664) );
AO32x1_ASAP7_75t_L g665 ( .A1(n_574), .A2(n_318), .A3(n_296), .B1(n_321), .B2(n_322), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_566), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_532), .A2(n_303), .B1(n_305), .B2(n_298), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_556), .B(n_430), .Y(n_668) );
OAI22xp5_ASAP7_75t_SL g669 ( .A1(n_558), .A2(n_442), .B1(n_282), .B2(n_391), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_563), .B(n_451), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_550), .B(n_479), .Y(n_671) );
INVx1_ASAP7_75t_SL g672 ( .A(n_565), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_526), .Y(n_673) );
A2O1A1Ixp33_ASAP7_75t_L g674 ( .A1(n_568), .A2(n_306), .B(n_323), .C(n_313), .Y(n_674) );
A2O1A1Ixp33_ASAP7_75t_SL g675 ( .A1(n_531), .A2(n_481), .B(n_315), .C(n_335), .Y(n_675) );
O2A1O1Ixp33_ASAP7_75t_L g676 ( .A1(n_570), .A2(n_347), .B(n_357), .C(n_345), .Y(n_676) );
BUFx6f_ASAP7_75t_L g677 ( .A(n_557), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_555), .B(n_365), .Y(n_678) );
BUFx2_ASAP7_75t_L g679 ( .A(n_585), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_526), .Y(n_680) );
BUFx6f_ASAP7_75t_L g681 ( .A(n_557), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_531), .A2(n_364), .B1(n_368), .B2(n_358), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_529), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_569), .A2(n_372), .B(n_371), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_576), .B(n_10), .Y(n_685) );
AND2x4_ASAP7_75t_L g686 ( .A(n_495), .B(n_451), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_572), .A2(n_381), .B(n_373), .Y(n_687) );
BUFx2_ASAP7_75t_L g688 ( .A(n_578), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_582), .A2(n_389), .B1(n_392), .B2(n_385), .Y(n_689) );
O2A1O1Ixp33_ASAP7_75t_L g690 ( .A1(n_587), .A2(n_396), .B(n_402), .C(n_394), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_529), .B(n_451), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_577), .A2(n_410), .B(n_405), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_496), .Y(n_693) );
O2A1O1Ixp33_ASAP7_75t_L g694 ( .A1(n_579), .A2(n_413), .B(n_403), .C(n_390), .Y(n_694) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_583), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_499), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_500), .A2(n_409), .B1(n_386), .B2(n_400), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_582), .A2(n_363), .B1(n_390), .B2(n_383), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_546), .B(n_11), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_581), .B(n_12), .Y(n_700) );
INVx2_ASAP7_75t_SL g701 ( .A(n_546), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_548), .B(n_279), .Y(n_702) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_548), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_586), .A2(n_403), .B1(n_383), .B2(n_370), .Y(n_704) );
AND2x4_ASAP7_75t_L g705 ( .A(n_586), .B(n_352), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_573), .Y(n_706) );
NAND3xp33_ASAP7_75t_L g707 ( .A(n_577), .B(n_333), .C(n_315), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_573), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_557), .Y(n_709) );
BUFx6f_ASAP7_75t_L g710 ( .A(n_557), .Y(n_710) );
AO21x1_ASAP7_75t_L g711 ( .A1(n_584), .A2(n_335), .B(n_333), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_584), .Y(n_712) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_584), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_584), .A2(n_369), .B(n_359), .Y(n_714) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_547), .B(n_12), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_547), .B(n_13), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_595), .Y(n_717) );
INVx2_ASAP7_75t_SL g718 ( .A(n_601), .Y(n_718) );
OAI21x1_ASAP7_75t_L g719 ( .A1(n_709), .A2(n_369), .B(n_359), .Y(n_719) );
INVx2_ASAP7_75t_L g720 ( .A(n_623), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_612), .Y(n_721) );
OA21x2_ASAP7_75t_L g722 ( .A1(n_711), .A2(n_370), .B(n_342), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_617), .B(n_13), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_679), .Y(n_724) );
AND2x4_ASAP7_75t_L g725 ( .A(n_645), .B(n_356), .Y(n_725) );
BUFx8_ASAP7_75t_L g726 ( .A(n_615), .Y(n_726) );
BUFx3_ASAP7_75t_L g727 ( .A(n_639), .Y(n_727) );
AO31x2_ASAP7_75t_L g728 ( .A1(n_614), .A2(n_354), .A3(n_342), .B(n_302), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_591), .Y(n_729) );
OAI21x1_ASAP7_75t_L g730 ( .A1(n_712), .A2(n_342), .B(n_302), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_606), .A2(n_354), .B1(n_342), .B2(n_302), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_672), .B(n_14), .Y(n_732) );
BUFx2_ASAP7_75t_R g733 ( .A(n_600), .Y(n_733) );
INVx6_ASAP7_75t_L g734 ( .A(n_645), .Y(n_734) );
OAI21x1_ASAP7_75t_L g735 ( .A1(n_634), .A2(n_354), .B(n_302), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_664), .A2(n_354), .B1(n_17), .B2(n_18), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_644), .B(n_16), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_650), .A2(n_17), .B1(n_19), .B2(n_20), .Y(n_738) );
BUFx2_ASAP7_75t_L g739 ( .A(n_628), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_653), .B(n_21), .Y(n_740) );
INVx3_ASAP7_75t_L g741 ( .A(n_658), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_657), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_662), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_650), .A2(n_22), .B1(n_23), .B2(n_24), .Y(n_744) );
NAND2x1p5_ASAP7_75t_L g745 ( .A(n_658), .B(n_22), .Y(n_745) );
BUFx3_ASAP7_75t_L g746 ( .A(n_639), .Y(n_746) );
NAND2x1p5_ASAP7_75t_L g747 ( .A(n_660), .B(n_24), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_666), .Y(n_748) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_588), .A2(n_25), .B1(n_26), .B2(n_27), .Y(n_749) );
INVx3_ASAP7_75t_L g750 ( .A(n_660), .Y(n_750) );
INVx3_ASAP7_75t_L g751 ( .A(n_639), .Y(n_751) );
INVxp33_ASAP7_75t_L g752 ( .A(n_599), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_602), .Y(n_753) );
BUFx4f_ASAP7_75t_L g754 ( .A(n_610), .Y(n_754) );
INVx2_ASAP7_75t_L g755 ( .A(n_627), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_602), .Y(n_756) );
OAI21x1_ASAP7_75t_L g757 ( .A1(n_663), .A2(n_86), .B(n_85), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_668), .Y(n_758) );
AOI22xp33_ASAP7_75t_SL g759 ( .A1(n_640), .A2(n_26), .B1(n_28), .B2(n_29), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_685), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g761 ( .A(n_656), .B(n_28), .Y(n_761) );
INVx6_ASAP7_75t_L g762 ( .A(n_655), .Y(n_762) );
BUFx3_ASAP7_75t_L g763 ( .A(n_655), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_669), .A2(n_29), .B1(n_30), .B2(n_31), .Y(n_764) );
INVx2_ASAP7_75t_L g765 ( .A(n_632), .Y(n_765) );
AO31x2_ASAP7_75t_L g766 ( .A1(n_654), .A2(n_31), .A3(n_32), .B(n_33), .Y(n_766) );
OR2x2_ASAP7_75t_L g767 ( .A(n_647), .B(n_32), .Y(n_767) );
BUFx3_ASAP7_75t_L g768 ( .A(n_655), .Y(n_768) );
BUFx6f_ASAP7_75t_L g769 ( .A(n_677), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_703), .A2(n_36), .B1(n_37), .B2(n_38), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_633), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_594), .B(n_36), .Y(n_772) );
OAI21x1_ASAP7_75t_SL g773 ( .A1(n_652), .A2(n_37), .B(n_39), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_636), .Y(n_774) );
BUFx10_ASAP7_75t_L g775 ( .A(n_659), .Y(n_775) );
OAI21x1_ASAP7_75t_L g776 ( .A1(n_714), .A2(n_93), .B(n_87), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_594), .B(n_39), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_638), .Y(n_778) );
OAI211xp5_ASAP7_75t_SL g779 ( .A1(n_621), .A2(n_41), .B(n_42), .C(n_43), .Y(n_779) );
NAND3xp33_ASAP7_75t_L g780 ( .A(n_625), .B(n_41), .C(n_42), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_642), .Y(n_781) );
NOR3xp33_ASAP7_75t_L g782 ( .A(n_651), .B(n_44), .C(n_45), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_637), .A2(n_47), .B1(n_48), .B2(n_49), .Y(n_783) );
OAI21x1_ASAP7_75t_L g784 ( .A1(n_622), .A2(n_97), .B(n_96), .Y(n_784) );
O2A1O1Ixp33_ASAP7_75t_SL g785 ( .A1(n_675), .A2(n_176), .B(n_269), .C(n_267), .Y(n_785) );
OA21x2_ASAP7_75t_L g786 ( .A1(n_707), .A2(n_100), .B(n_98), .Y(n_786) );
AOI22xp33_ASAP7_75t_SL g787 ( .A1(n_715), .A2(n_47), .B1(n_49), .B2(n_50), .Y(n_787) );
AND2x2_ASAP7_75t_L g788 ( .A(n_598), .B(n_50), .Y(n_788) );
OA21x2_ASAP7_75t_L g789 ( .A1(n_702), .A2(n_179), .B(n_266), .Y(n_789) );
OA21x2_ASAP7_75t_L g790 ( .A1(n_684), .A2(n_177), .B(n_265), .Y(n_790) );
OA21x2_ASAP7_75t_L g791 ( .A1(n_687), .A2(n_173), .B(n_264), .Y(n_791) );
BUFx8_ASAP7_75t_L g792 ( .A(n_648), .Y(n_792) );
OAI21x1_ASAP7_75t_L g793 ( .A1(n_706), .A2(n_170), .B(n_263), .Y(n_793) );
INVx2_ASAP7_75t_L g794 ( .A(n_673), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_688), .B(n_51), .Y(n_795) );
OAI21x1_ASAP7_75t_L g796 ( .A1(n_708), .A2(n_169), .B(n_262), .Y(n_796) );
AOI21xp5_ASAP7_75t_L g797 ( .A1(n_691), .A2(n_168), .B(n_261), .Y(n_797) );
INVx2_ASAP7_75t_SL g798 ( .A(n_605), .Y(n_798) );
OAI21x1_ASAP7_75t_L g799 ( .A1(n_618), .A2(n_167), .B(n_259), .Y(n_799) );
OAI22x1_ASAP7_75t_L g800 ( .A1(n_667), .A2(n_51), .B1(n_52), .B2(n_54), .Y(n_800) );
O2A1O1Ixp33_ASAP7_75t_SL g801 ( .A1(n_713), .A2(n_181), .B(n_258), .C(n_257), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_643), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_649), .Y(n_803) );
AND2x4_ASAP7_75t_L g804 ( .A(n_661), .B(n_54), .Y(n_804) );
INVx1_ASAP7_75t_SL g805 ( .A(n_695), .Y(n_805) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_597), .B(n_55), .Y(n_806) );
OAI22xp33_ASAP7_75t_L g807 ( .A1(n_605), .A2(n_56), .B1(n_57), .B2(n_58), .Y(n_807) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_626), .B(n_58), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_680), .Y(n_809) );
INVx4_ASAP7_75t_L g810 ( .A(n_608), .Y(n_810) );
OAI21x1_ASAP7_75t_L g811 ( .A1(n_670), .A2(n_182), .B(n_256), .Y(n_811) );
AND2x2_ASAP7_75t_L g812 ( .A(n_613), .B(n_59), .Y(n_812) );
AOI221xp5_ASAP7_75t_L g813 ( .A1(n_641), .A2(n_59), .B1(n_60), .B2(n_61), .C(n_62), .Y(n_813) );
OAI21x1_ASAP7_75t_L g814 ( .A1(n_630), .A2(n_185), .B(n_255), .Y(n_814) );
OAI21x1_ASAP7_75t_L g815 ( .A1(n_646), .A2(n_164), .B(n_253), .Y(n_815) );
OAI21x1_ASAP7_75t_L g816 ( .A1(n_682), .A2(n_163), .B(n_251), .Y(n_816) );
INVx4_ASAP7_75t_L g817 ( .A(n_608), .Y(n_817) );
OAI21xp5_ASAP7_75t_L g818 ( .A1(n_620), .A2(n_160), .B(n_250), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_678), .B(n_62), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_699), .Y(n_820) );
NAND2xp5_ASAP7_75t_SL g821 ( .A(n_593), .B(n_102), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_607), .A2(n_63), .B1(n_64), .B2(n_66), .Y(n_822) );
A2O1A1Ixp33_ASAP7_75t_L g823 ( .A1(n_619), .A2(n_64), .B(n_66), .C(n_67), .Y(n_823) );
BUFx3_ASAP7_75t_L g824 ( .A(n_661), .Y(n_824) );
AO31x2_ASAP7_75t_L g825 ( .A1(n_698), .A2(n_68), .A3(n_69), .B(n_70), .Y(n_825) );
AOI222xp33_ASAP7_75t_L g826 ( .A1(n_716), .A2(n_69), .B1(n_103), .B2(n_106), .C1(n_108), .C2(n_110), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_700), .A2(n_111), .B1(n_112), .B2(n_113), .Y(n_827) );
BUFx2_ASAP7_75t_L g828 ( .A(n_659), .Y(n_828) );
BUFx12f_ASAP7_75t_L g829 ( .A(n_659), .Y(n_829) );
O2A1O1Ixp33_ASAP7_75t_SL g830 ( .A1(n_674), .A2(n_115), .B(n_116), .C(n_118), .Y(n_830) );
AO21x2_ASAP7_75t_L g831 ( .A1(n_692), .A2(n_119), .B(n_123), .Y(n_831) );
INVx2_ASAP7_75t_L g832 ( .A(n_683), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_693), .Y(n_833) );
OAI21x1_ASAP7_75t_L g834 ( .A1(n_696), .A2(n_132), .B(n_134), .Y(n_834) );
HB1xp67_ASAP7_75t_L g835 ( .A(n_661), .Y(n_835) );
BUFx2_ASAP7_75t_L g836 ( .A(n_659), .Y(n_836) );
INVx3_ASAP7_75t_L g837 ( .A(n_593), .Y(n_837) );
AO221x2_ASAP7_75t_L g838 ( .A1(n_704), .A2(n_138), .B1(n_139), .B2(n_141), .C(n_142), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_611), .A2(n_143), .B1(n_146), .B2(n_149), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_701), .Y(n_840) );
OAI21xp5_ASAP7_75t_L g841 ( .A1(n_671), .A2(n_151), .B(n_153), .Y(n_841) );
AOI21x1_ASAP7_75t_L g842 ( .A1(n_705), .A2(n_155), .B(n_156), .Y(n_842) );
O2A1O1Ixp33_ASAP7_75t_SL g843 ( .A1(n_603), .A2(n_157), .B(n_159), .C(n_186), .Y(n_843) );
CKINVDCx5p33_ASAP7_75t_R g844 ( .A(n_624), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_589), .Y(n_845) );
AND2x4_ASAP7_75t_L g846 ( .A(n_593), .B(n_187), .Y(n_846) );
OAI22xp5_ASAP7_75t_L g847 ( .A1(n_705), .A2(n_190), .B1(n_191), .B2(n_193), .Y(n_847) );
HB1xp67_ASAP7_75t_L g848 ( .A(n_596), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_590), .Y(n_849) );
OAI21x1_ASAP7_75t_L g850 ( .A1(n_694), .A2(n_194), .B(n_195), .Y(n_850) );
BUFx3_ASAP7_75t_L g851 ( .A(n_596), .Y(n_851) );
INVx2_ASAP7_75t_L g852 ( .A(n_596), .Y(n_852) );
HB1xp67_ASAP7_75t_L g853 ( .A(n_604), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_592), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_758), .B(n_676), .Y(n_855) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_752), .A2(n_690), .B1(n_689), .B2(n_604), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_721), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_729), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_752), .A2(n_631), .B1(n_609), .B2(n_616), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_742), .Y(n_860) );
AND2x2_ASAP7_75t_L g861 ( .A(n_795), .B(n_697), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_743), .Y(n_862) );
BUFx12f_ASAP7_75t_L g863 ( .A(n_726), .Y(n_863) );
NOR2xp33_ASAP7_75t_L g864 ( .A(n_724), .B(n_686), .Y(n_864) );
OAI22xp33_ASAP7_75t_L g865 ( .A1(n_745), .A2(n_604), .B1(n_635), .B2(n_681), .Y(n_865) );
CKINVDCx5p33_ASAP7_75t_R g866 ( .A(n_733), .Y(n_866) );
AND2x2_ASAP7_75t_L g867 ( .A(n_795), .B(n_635), .Y(n_867) );
AOI221xp5_ASAP7_75t_L g868 ( .A1(n_760), .A2(n_629), .B1(n_686), .B2(n_635), .C(n_665), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_748), .B(n_710), .Y(n_869) );
AOI221xp5_ASAP7_75t_L g870 ( .A1(n_806), .A2(n_665), .B1(n_681), .B2(n_677), .C(n_710), .Y(n_870) );
AOI21xp5_ASAP7_75t_L g871 ( .A1(n_785), .A2(n_710), .B(n_681), .Y(n_871) );
OAI221xp5_ASAP7_75t_L g872 ( .A1(n_736), .A2(n_665), .B1(n_201), .B2(n_203), .C(n_205), .Y(n_872) );
OR3x1_ASAP7_75t_L g873 ( .A(n_779), .B(n_200), .C(n_207), .Y(n_873) );
OR2x2_ASAP7_75t_L g874 ( .A(n_805), .B(n_209), .Y(n_874) );
INVx2_ASAP7_75t_L g875 ( .A(n_717), .Y(n_875) );
OAI21x1_ASAP7_75t_L g876 ( .A1(n_735), .A2(n_210), .B(n_211), .Y(n_876) );
A2O1A1Ixp33_ASAP7_75t_L g877 ( .A1(n_819), .A2(n_213), .B(n_215), .C(n_216), .Y(n_877) );
NOR2x1p5_ASAP7_75t_L g878 ( .A(n_810), .B(n_217), .Y(n_878) );
OAI21xp5_ASAP7_75t_L g879 ( .A1(n_808), .A2(n_218), .B(n_220), .Y(n_879) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_736), .A2(n_221), .B1(n_223), .B2(n_224), .Y(n_880) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_738), .A2(n_225), .B1(n_229), .B2(n_230), .Y(n_881) );
AOI222xp33_ASAP7_75t_L g882 ( .A1(n_754), .A2(n_233), .B1(n_234), .B2(n_239), .C1(n_240), .C2(n_242), .Y(n_882) );
AOI221xp5_ASAP7_75t_L g883 ( .A1(n_806), .A2(n_243), .B1(n_244), .B2(n_245), .C(n_246), .Y(n_883) );
CKINVDCx5p33_ASAP7_75t_R g884 ( .A(n_754), .Y(n_884) );
OAI22xp5_ASAP7_75t_L g885 ( .A1(n_738), .A2(n_248), .B1(n_249), .B2(n_270), .Y(n_885) );
CKINVDCx5p33_ASAP7_75t_R g886 ( .A(n_844), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_771), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_774), .Y(n_888) );
INVx3_ASAP7_75t_L g889 ( .A(n_734), .Y(n_889) );
CKINVDCx5p33_ASAP7_75t_R g890 ( .A(n_792), .Y(n_890) );
AOI22xp33_ASAP7_75t_SL g891 ( .A1(n_838), .A2(n_745), .B1(n_747), .B2(n_819), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_782), .A2(n_854), .B1(n_761), .B2(n_779), .Y(n_892) );
OA21x2_ASAP7_75t_L g893 ( .A1(n_719), .A2(n_793), .B(n_834), .Y(n_893) );
HB1xp67_ASAP7_75t_L g894 ( .A(n_717), .Y(n_894) );
OAI22xp33_ASAP7_75t_L g895 ( .A1(n_747), .A2(n_807), .B1(n_800), .B2(n_749), .Y(n_895) );
BUFx3_ASAP7_75t_L g896 ( .A(n_792), .Y(n_896) );
NOR2xp33_ASAP7_75t_SL g897 ( .A(n_810), .B(n_817), .Y(n_897) );
OAI22xp5_ASAP7_75t_SL g898 ( .A1(n_759), .A2(n_764), .B1(n_744), .B2(n_787), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_802), .Y(n_899) );
AOI321xp33_ASAP7_75t_L g900 ( .A1(n_764), .A2(n_782), .A3(n_744), .B1(n_731), .B2(n_807), .C(n_783), .Y(n_900) );
INVx2_ASAP7_75t_SL g901 ( .A(n_726), .Y(n_901) );
CKINVDCx11_ASAP7_75t_R g902 ( .A(n_739), .Y(n_902) );
O2A1O1Ixp33_ASAP7_75t_L g903 ( .A1(n_737), .A2(n_823), .B(n_761), .C(n_773), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_808), .A2(n_731), .B1(n_788), .B2(n_759), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_753), .B(n_756), .Y(n_905) );
BUFx6f_ASAP7_75t_L g906 ( .A(n_769), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_820), .A2(n_813), .B1(n_780), .B2(n_787), .Y(n_907) );
INVx2_ASAP7_75t_SL g908 ( .A(n_817), .Y(n_908) );
AOI21x1_ASAP7_75t_L g909 ( .A1(n_722), .A2(n_842), .B(n_821), .Y(n_909) );
OAI21xp5_ASAP7_75t_L g910 ( .A1(n_723), .A2(n_772), .B(n_777), .Y(n_910) );
OAI22xp33_ASAP7_75t_L g911 ( .A1(n_770), .A2(n_767), .B1(n_829), .B2(n_828), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_833), .B(n_803), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_838), .A2(n_783), .B1(n_812), .B2(n_822), .Y(n_913) );
NAND3xp33_ASAP7_75t_SL g914 ( .A(n_826), .B(n_822), .C(n_823), .Y(n_914) );
AOI21xp5_ASAP7_75t_L g915 ( .A1(n_720), .A2(n_809), .B(n_778), .Y(n_915) );
AOI332xp33_ASAP7_75t_L g916 ( .A1(n_740), .A2(n_732), .A3(n_725), .B1(n_750), .B2(n_741), .B3(n_804), .C1(n_845), .C2(n_849), .Y(n_916) );
A2O1A1Ixp33_ASAP7_75t_L g917 ( .A1(n_818), .A2(n_778), .B(n_809), .C(n_841), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_825), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_718), .B(n_741), .Y(n_919) );
AOI21xp5_ASAP7_75t_L g920 ( .A1(n_830), .A2(n_769), .B(n_801), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_825), .Y(n_921) );
AOI222xp33_ASAP7_75t_L g922 ( .A1(n_798), .A2(n_804), .B1(n_725), .B2(n_750), .C1(n_847), .C2(n_836), .Y(n_922) );
INVx2_ASAP7_75t_L g923 ( .A(n_755), .Y(n_923) );
INVx2_ASAP7_75t_L g924 ( .A(n_765), .Y(n_924) );
INVx2_ASAP7_75t_L g925 ( .A(n_781), .Y(n_925) );
AOI22xp5_ASAP7_75t_L g926 ( .A1(n_734), .A2(n_840), .B1(n_838), .B2(n_832), .Y(n_926) );
AND2x2_ASAP7_75t_L g927 ( .A(n_794), .B(n_734), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_825), .Y(n_928) );
AND2x2_ASAP7_75t_L g929 ( .A(n_825), .B(n_766), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_827), .A2(n_839), .B1(n_831), .B2(n_835), .Y(n_930) );
AOI221xp5_ASAP7_75t_L g931 ( .A1(n_843), .A2(n_801), .B1(n_797), .B2(n_835), .C(n_846), .Y(n_931) );
AOI21xp33_ASAP7_75t_L g932 ( .A1(n_848), .A2(n_853), .B(n_751), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_766), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_831), .A2(n_746), .B1(n_727), .B2(n_768), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_727), .A2(n_763), .B1(n_768), .B2(n_746), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_763), .A2(n_824), .B1(n_846), .B2(n_762), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_766), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_824), .B(n_751), .Y(n_938) );
OAI22xp5_ASAP7_75t_L g939 ( .A1(n_762), .A2(n_853), .B1(n_848), .B2(n_851), .Y(n_939) );
INVx2_ASAP7_75t_L g940 ( .A(n_728), .Y(n_940) );
OA21x2_ASAP7_75t_L g941 ( .A1(n_730), .A2(n_796), .B(n_850), .Y(n_941) );
OAI22xp33_ASAP7_75t_SL g942 ( .A1(n_762), .A2(n_821), .B1(n_837), .B2(n_851), .Y(n_942) );
HB1xp67_ASAP7_75t_L g943 ( .A(n_837), .Y(n_943) );
AOI21xp5_ASAP7_75t_L g944 ( .A1(n_769), .A2(n_789), .B(n_722), .Y(n_944) );
INVx2_ASAP7_75t_L g945 ( .A(n_728), .Y(n_945) );
INVx2_ASAP7_75t_SL g946 ( .A(n_775), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_775), .A2(n_722), .B1(n_791), .B2(n_790), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g948 ( .A(n_766), .B(n_852), .Y(n_948) );
AND2x2_ASAP7_75t_L g949 ( .A(n_728), .B(n_816), .Y(n_949) );
AOI21xp5_ASAP7_75t_L g950 ( .A1(n_789), .A2(n_790), .B(n_791), .Y(n_950) );
AO21x2_ASAP7_75t_L g951 ( .A1(n_811), .A2(n_757), .B(n_784), .Y(n_951) );
CKINVDCx20_ASAP7_75t_R g952 ( .A(n_786), .Y(n_952) );
AOI222xp33_ASAP7_75t_L g953 ( .A1(n_799), .A2(n_523), .B1(n_606), .B2(n_458), .C1(n_640), .C2(n_656), .Y(n_953) );
OAI21x1_ASAP7_75t_L g954 ( .A1(n_814), .A2(n_815), .B(n_776), .Y(n_954) );
AND2x4_ASAP7_75t_L g955 ( .A(n_786), .B(n_810), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_786), .A2(n_752), .B1(n_523), .B2(n_782), .Y(n_956) );
AOI22xp33_ASAP7_75t_SL g957 ( .A1(n_838), .A2(n_523), .B1(n_538), .B2(n_522), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_752), .A2(n_523), .B1(n_782), .B2(n_736), .Y(n_958) );
AND2x2_ASAP7_75t_L g959 ( .A(n_795), .B(n_547), .Y(n_959) );
OAI21x1_ASAP7_75t_L g960 ( .A1(n_735), .A2(n_730), .B(n_719), .Y(n_960) );
INVx2_ASAP7_75t_L g961 ( .A(n_729), .Y(n_961) );
INVx2_ASAP7_75t_L g962 ( .A(n_729), .Y(n_962) );
INVx2_ASAP7_75t_L g963 ( .A(n_729), .Y(n_963) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_758), .B(n_530), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_758), .B(n_530), .Y(n_965) );
HB1xp67_ASAP7_75t_L g966 ( .A(n_717), .Y(n_966) );
AOI33xp33_ASAP7_75t_L g967 ( .A1(n_759), .A2(n_641), .A3(n_440), .B1(n_441), .B2(n_656), .B3(n_787), .Y(n_967) );
AOI221xp5_ASAP7_75t_L g968 ( .A1(n_752), .A2(n_458), .B1(n_523), .B2(n_547), .C(n_598), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_721), .Y(n_969) );
INVx2_ASAP7_75t_L g970 ( .A(n_729), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_752), .A2(n_523), .B1(n_782), .B2(n_736), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_752), .A2(n_523), .B1(n_782), .B2(n_736), .Y(n_972) );
OAI22xp5_ASAP7_75t_L g973 ( .A1(n_752), .A2(n_588), .B1(n_650), .B2(n_571), .Y(n_973) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_752), .A2(n_588), .B1(n_650), .B2(n_571), .Y(n_974) );
INVx2_ASAP7_75t_L g975 ( .A(n_729), .Y(n_975) );
OA21x2_ASAP7_75t_L g976 ( .A1(n_735), .A2(n_719), .B(n_793), .Y(n_976) );
AND2x4_ASAP7_75t_L g977 ( .A(n_810), .B(n_817), .Y(n_977) );
HB1xp67_ASAP7_75t_L g978 ( .A(n_717), .Y(n_978) );
AOI21xp33_ASAP7_75t_SL g979 ( .A1(n_844), .A2(n_470), .B(n_600), .Y(n_979) );
OAI221xp5_ASAP7_75t_L g980 ( .A1(n_958), .A2(n_971), .B1(n_972), .B2(n_968), .C(n_957), .Y(n_980) );
AOI22xp33_ASAP7_75t_SL g981 ( .A1(n_898), .A2(n_974), .B1(n_973), .B2(n_957), .Y(n_981) );
AO31x2_ASAP7_75t_L g982 ( .A1(n_933), .A2(n_937), .A3(n_918), .B(n_928), .Y(n_982) );
INVx2_ASAP7_75t_L g983 ( .A(n_894), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_894), .B(n_966), .Y(n_984) );
BUFx6f_ASAP7_75t_L g985 ( .A(n_906), .Y(n_985) );
AND2x2_ASAP7_75t_L g986 ( .A(n_966), .B(n_978), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_978), .Y(n_987) );
AOI221xp5_ASAP7_75t_L g988 ( .A1(n_958), .A2(n_972), .B1(n_971), .B2(n_895), .C(n_959), .Y(n_988) );
INVxp67_ASAP7_75t_SL g989 ( .A(n_875), .Y(n_989) );
AND2x2_ASAP7_75t_L g990 ( .A(n_923), .B(n_924), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_857), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_860), .Y(n_992) );
OR2x2_ASAP7_75t_L g993 ( .A(n_921), .B(n_858), .Y(n_993) );
NOR2x1_ASAP7_75t_L g994 ( .A(n_878), .B(n_896), .Y(n_994) );
BUFx2_ASAP7_75t_L g995 ( .A(n_906), .Y(n_995) );
INVx2_ASAP7_75t_L g996 ( .A(n_940), .Y(n_996) );
AND2x2_ASAP7_75t_L g997 ( .A(n_925), .B(n_961), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_862), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_887), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_888), .Y(n_1000) );
INVxp67_ASAP7_75t_L g1001 ( .A(n_964), .Y(n_1001) );
INVx2_ASAP7_75t_L g1002 ( .A(n_945), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_962), .B(n_963), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_899), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_970), .B(n_975), .Y(n_1005) );
OR2x2_ASAP7_75t_L g1006 ( .A(n_912), .B(n_969), .Y(n_1006) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_967), .B(n_953), .Y(n_1007) );
HB1xp67_ASAP7_75t_L g1008 ( .A(n_927), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_929), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_948), .Y(n_1010) );
INVx1_ASAP7_75t_L g1011 ( .A(n_869), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_914), .A2(n_913), .B1(n_895), .B2(n_891), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_891), .B(n_892), .Y(n_1013) );
CKINVDCx5p33_ASAP7_75t_R g1014 ( .A(n_863), .Y(n_1014) );
AND2x2_ASAP7_75t_L g1015 ( .A(n_892), .B(n_956), .Y(n_1015) );
NAND3xp33_ASAP7_75t_L g1016 ( .A(n_956), .B(n_900), .C(n_882), .Y(n_1016) );
INVxp33_ASAP7_75t_L g1017 ( .A(n_902), .Y(n_1017) );
NAND2xp5_ASAP7_75t_L g1018 ( .A(n_861), .B(n_965), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_867), .B(n_913), .Y(n_1019) );
OR2x6_ASAP7_75t_L g1020 ( .A(n_955), .B(n_903), .Y(n_1020) );
INVx2_ASAP7_75t_L g1021 ( .A(n_906), .Y(n_1021) );
OA21x2_ASAP7_75t_L g1022 ( .A1(n_950), .A2(n_944), .B(n_947), .Y(n_1022) );
OR2x2_ASAP7_75t_L g1023 ( .A(n_905), .B(n_855), .Y(n_1023) );
HB1xp67_ASAP7_75t_L g1024 ( .A(n_864), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_919), .Y(n_1025) );
INVx2_ASAP7_75t_L g1026 ( .A(n_906), .Y(n_1026) );
INVx2_ASAP7_75t_L g1027 ( .A(n_976), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_907), .B(n_904), .Y(n_1028) );
OR2x6_ASAP7_75t_L g1029 ( .A(n_955), .B(n_946), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_864), .Y(n_1030) );
INVxp67_ASAP7_75t_SL g1031 ( .A(n_865), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_907), .B(n_904), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_915), .B(n_926), .Y(n_1033) );
OR2x2_ASAP7_75t_L g1034 ( .A(n_943), .B(n_911), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g1035 ( .A(n_911), .B(n_977), .Y(n_1035) );
INVx2_ASAP7_75t_SL g1036 ( .A(n_977), .Y(n_1036) );
OAI22xp33_ASAP7_75t_L g1037 ( .A1(n_897), .A2(n_872), .B1(n_866), .B2(n_901), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_943), .Y(n_1038) );
INVx2_ASAP7_75t_L g1039 ( .A(n_876), .Y(n_1039) );
NOR2x1p5_ASAP7_75t_L g1040 ( .A(n_890), .B(n_884), .Y(n_1040) );
INVx2_ASAP7_75t_L g1041 ( .A(n_960), .Y(n_1041) );
HB1xp67_ASAP7_75t_L g1042 ( .A(n_889), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_874), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_908), .Y(n_1044) );
OR2x2_ASAP7_75t_L g1045 ( .A(n_938), .B(n_910), .Y(n_1045) );
BUFx3_ASAP7_75t_L g1046 ( .A(n_889), .Y(n_1046) );
INVx5_ASAP7_75t_SL g1047 ( .A(n_865), .Y(n_1047) );
OR2x2_ASAP7_75t_L g1048 ( .A(n_939), .B(n_936), .Y(n_1048) );
OAI22xp5_ASAP7_75t_L g1049 ( .A1(n_859), .A2(n_936), .B1(n_873), .B2(n_856), .Y(n_1049) );
INVx2_ASAP7_75t_L g1050 ( .A(n_949), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g1051 ( .A(n_859), .B(n_922), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_880), .Y(n_1052) );
BUFx2_ASAP7_75t_L g1053 ( .A(n_952), .Y(n_1053) );
INVx1_ASAP7_75t_SL g1054 ( .A(n_886), .Y(n_1054) );
HB1xp67_ASAP7_75t_L g1055 ( .A(n_932), .Y(n_1055) );
INVxp67_ASAP7_75t_SL g1056 ( .A(n_935), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g1057 ( .A(n_979), .B(n_935), .Y(n_1057) );
INVx1_ASAP7_75t_L g1058 ( .A(n_881), .Y(n_1058) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_868), .B(n_930), .Y(n_1059) );
BUFx6f_ASAP7_75t_L g1060 ( .A(n_954), .Y(n_1060) );
BUFx3_ASAP7_75t_L g1061 ( .A(n_893), .Y(n_1061) );
INVx2_ASAP7_75t_L g1062 ( .A(n_893), .Y(n_1062) );
HB1xp67_ASAP7_75t_L g1063 ( .A(n_879), .Y(n_1063) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_934), .B(n_930), .Y(n_1064) );
BUFx6f_ASAP7_75t_L g1065 ( .A(n_941), .Y(n_1065) );
INVx2_ASAP7_75t_SL g1066 ( .A(n_885), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_877), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_883), .A2(n_870), .B1(n_916), .B2(n_931), .Y(n_1068) );
INVxp67_ASAP7_75t_SL g1069 ( .A(n_942), .Y(n_1069) );
OR2x2_ASAP7_75t_L g1070 ( .A(n_934), .B(n_917), .Y(n_1070) );
BUFx2_ASAP7_75t_L g1071 ( .A(n_941), .Y(n_1071) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_947), .B(n_951), .Y(n_1072) );
INVx2_ASAP7_75t_SL g1073 ( .A(n_941), .Y(n_1073) );
INVx2_ASAP7_75t_L g1074 ( .A(n_909), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1009), .B(n_920), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1076 ( .A(n_1007), .B(n_871), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_1028), .B(n_1032), .Y(n_1077) );
INVx1_ASAP7_75t_L g1078 ( .A(n_993), .Y(n_1078) );
NAND2xp5_ASAP7_75t_L g1079 ( .A(n_1028), .B(n_1032), .Y(n_1079) );
AND2x4_ASAP7_75t_L g1080 ( .A(n_1009), .B(n_1050), .Y(n_1080) );
INVx2_ASAP7_75t_L g1081 ( .A(n_1027), .Y(n_1081) );
INVxp67_ASAP7_75t_SL g1082 ( .A(n_984), .Y(n_1082) );
AND2x2_ASAP7_75t_SL g1083 ( .A(n_1053), .B(n_1034), .Y(n_1083) );
OAI211xp5_ASAP7_75t_SL g1084 ( .A1(n_988), .A2(n_980), .B(n_1025), .C(n_1044), .Y(n_1084) );
INVx1_ASAP7_75t_L g1085 ( .A(n_993), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_1003), .B(n_1005), .Y(n_1086) );
INVx1_ASAP7_75t_L g1087 ( .A(n_982), .Y(n_1087) );
HB1xp67_ASAP7_75t_L g1088 ( .A(n_984), .Y(n_1088) );
INVx1_ASAP7_75t_L g1089 ( .A(n_982), .Y(n_1089) );
NAND2xp5_ASAP7_75t_L g1090 ( .A(n_1003), .B(n_1005), .Y(n_1090) );
OR2x2_ASAP7_75t_L g1091 ( .A(n_987), .B(n_983), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_1019), .B(n_986), .Y(n_1092) );
NOR2xp33_ASAP7_75t_L g1093 ( .A(n_1017), .B(n_1054), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1094 ( .A(n_1019), .B(n_986), .Y(n_1094) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_1015), .B(n_983), .Y(n_1095) );
NAND2x1_ASAP7_75t_L g1096 ( .A(n_1020), .B(n_1029), .Y(n_1096) );
OAI221xp5_ASAP7_75t_L g1097 ( .A1(n_981), .A2(n_1016), .B1(n_1012), .B2(n_1018), .C(n_1001), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_1015), .B(n_1013), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g1099 ( .A(n_997), .B(n_1006), .Y(n_1099) );
NOR2xp67_ASAP7_75t_R g1100 ( .A(n_1053), .B(n_994), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1013), .B(n_1050), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g1102 ( .A1(n_1051), .A2(n_1035), .B1(n_1034), .B2(n_1049), .Y(n_1102) );
OAI21xp33_ASAP7_75t_L g1103 ( .A1(n_1068), .A2(n_1069), .B(n_1064), .Y(n_1103) );
OR2x2_ASAP7_75t_L g1104 ( .A(n_987), .B(n_1038), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_1064), .B(n_997), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_1010), .B(n_990), .Y(n_1106) );
AND2x4_ASAP7_75t_L g1107 ( .A(n_1029), .B(n_1020), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1010), .B(n_990), .Y(n_1108) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_1006), .B(n_991), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_982), .B(n_1033), .Y(n_1110) );
INVxp67_ASAP7_75t_SL g1111 ( .A(n_989), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_1066), .A2(n_1024), .B1(n_1052), .B2(n_1048), .Y(n_1112) );
AOI221xp5_ASAP7_75t_L g1113 ( .A1(n_1030), .A2(n_1043), .B1(n_998), .B2(n_992), .C(n_1004), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_982), .Y(n_1114) );
AOI33xp33_ASAP7_75t_L g1115 ( .A1(n_999), .A2(n_1000), .A3(n_1038), .B1(n_1037), .B2(n_1072), .B3(n_1036), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_996), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1117 ( .A(n_1033), .B(n_1072), .Y(n_1117) );
OAI33xp33_ASAP7_75t_L g1118 ( .A1(n_1045), .A2(n_1057), .A3(n_1023), .B1(n_1059), .B2(n_1070), .B3(n_1014), .Y(n_1118) );
INVx2_ASAP7_75t_SL g1119 ( .A(n_1036), .Y(n_1119) );
INVx1_ASAP7_75t_SL g1120 ( .A(n_1014), .Y(n_1120) );
BUFx3_ASAP7_75t_L g1121 ( .A(n_1046), .Y(n_1121) );
HB1xp67_ASAP7_75t_L g1122 ( .A(n_1008), .Y(n_1122) );
OR2x2_ASAP7_75t_L g1123 ( .A(n_1045), .B(n_1023), .Y(n_1123) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1002), .Y(n_1124) );
INVx2_ASAP7_75t_SL g1125 ( .A(n_1029), .Y(n_1125) );
NAND2xp5_ASAP7_75t_L g1126 ( .A(n_1011), .B(n_1042), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_1002), .B(n_1011), .Y(n_1127) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_1020), .B(n_1070), .Y(n_1128) );
INVx4_ASAP7_75t_L g1129 ( .A(n_995), .Y(n_1129) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1071), .Y(n_1130) );
INVxp67_ASAP7_75t_L g1131 ( .A(n_1046), .Y(n_1131) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_1066), .A2(n_1048), .B1(n_1058), .B2(n_1056), .Y(n_1132) );
AND2x4_ASAP7_75t_L g1133 ( .A(n_1029), .B(n_1020), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1062), .Y(n_1134) );
OAI21xp33_ASAP7_75t_L g1135 ( .A1(n_1055), .A2(n_1017), .B(n_1063), .Y(n_1135) );
HB1xp67_ASAP7_75t_L g1136 ( .A(n_995), .Y(n_1136) );
INVxp67_ASAP7_75t_L g1137 ( .A(n_1040), .Y(n_1137) );
INVx4_ASAP7_75t_L g1138 ( .A(n_985), .Y(n_1138) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1073), .Y(n_1139) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_1117), .B(n_1022), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1117), .B(n_1022), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1110), .B(n_1022), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1143 ( .A(n_1110), .B(n_1061), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1105), .B(n_1061), .Y(n_1144) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_1098), .B(n_1031), .Y(n_1145) );
AND2x4_ASAP7_75t_L g1146 ( .A(n_1107), .B(n_1133), .Y(n_1146) );
OR2x2_ASAP7_75t_L g1147 ( .A(n_1088), .B(n_1047), .Y(n_1147) );
OR2x2_ASAP7_75t_L g1148 ( .A(n_1082), .B(n_1047), .Y(n_1148) );
BUFx2_ASAP7_75t_SL g1149 ( .A(n_1111), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1116), .Y(n_1150) );
OR2x2_ASAP7_75t_L g1151 ( .A(n_1092), .B(n_1047), .Y(n_1151) );
AND2x4_ASAP7_75t_L g1152 ( .A(n_1107), .B(n_1065), .Y(n_1152) );
AND3x2_ASAP7_75t_L g1153 ( .A(n_1137), .B(n_1067), .C(n_1047), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_1105), .B(n_1065), .Y(n_1154) );
INVxp67_ASAP7_75t_L g1155 ( .A(n_1122), .Y(n_1155) );
INVx2_ASAP7_75t_L g1156 ( .A(n_1081), .Y(n_1156) );
HB1xp67_ASAP7_75t_L g1157 ( .A(n_1136), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1124), .Y(n_1158) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_1092), .B(n_1065), .Y(n_1159) );
NOR2xp67_ASAP7_75t_L g1160 ( .A(n_1135), .B(n_1074), .Y(n_1160) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1127), .Y(n_1161) );
HB1xp67_ASAP7_75t_L g1162 ( .A(n_1091), .Y(n_1162) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1127), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1164 ( .A(n_1098), .B(n_1021), .Y(n_1164) );
NOR2xp33_ASAP7_75t_SL g1165 ( .A(n_1120), .B(n_1093), .Y(n_1165) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1080), .Y(n_1166) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1080), .Y(n_1167) );
HB1xp67_ASAP7_75t_L g1168 ( .A(n_1091), .Y(n_1168) );
OR2x2_ASAP7_75t_L g1169 ( .A(n_1094), .B(n_1041), .Y(n_1169) );
AND2x2_ASAP7_75t_L g1170 ( .A(n_1101), .B(n_1041), .Y(n_1170) );
BUFx2_ASAP7_75t_L g1171 ( .A(n_1129), .Y(n_1171) );
NOR2x1_ASAP7_75t_L g1172 ( .A(n_1121), .B(n_1021), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1080), .Y(n_1173) );
OR2x2_ASAP7_75t_L g1174 ( .A(n_1123), .B(n_1026), .Y(n_1174) );
NOR3xp33_ASAP7_75t_L g1175 ( .A(n_1097), .B(n_1026), .C(n_1039), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1134), .Y(n_1176) );
NOR2x1p5_ASAP7_75t_L g1177 ( .A(n_1096), .B(n_1039), .Y(n_1177) );
HB1xp67_ASAP7_75t_L g1178 ( .A(n_1126), .Y(n_1178) );
OAI211xp5_ASAP7_75t_L g1179 ( .A1(n_1103), .A2(n_985), .B(n_1060), .C(n_1102), .Y(n_1179) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1134), .Y(n_1180) );
NAND2xp33_ASAP7_75t_SL g1181 ( .A(n_1096), .B(n_985), .Y(n_1181) );
AOI21xp33_ASAP7_75t_SL g1182 ( .A1(n_1083), .A2(n_1060), .B(n_1133), .Y(n_1182) );
NOR3xp33_ASAP7_75t_L g1183 ( .A(n_1118), .B(n_1060), .C(n_1084), .Y(n_1183) );
OR2x2_ASAP7_75t_L g1184 ( .A(n_1123), .B(n_1095), .Y(n_1184) );
HB1xp67_ASAP7_75t_L g1185 ( .A(n_1121), .Y(n_1185) );
OR2x2_ASAP7_75t_L g1186 ( .A(n_1104), .B(n_1078), .Y(n_1186) );
INVx3_ASAP7_75t_L g1187 ( .A(n_1138), .Y(n_1187) );
NAND3xp33_ASAP7_75t_L g1188 ( .A(n_1076), .B(n_1113), .C(n_1115), .Y(n_1188) );
INVxp67_ASAP7_75t_L g1189 ( .A(n_1100), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1128), .B(n_1075), .Y(n_1190) );
CKINVDCx20_ASAP7_75t_R g1191 ( .A(n_1086), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1140), .B(n_1128), .Y(n_1192) );
NAND2xp5_ASAP7_75t_L g1193 ( .A(n_1178), .B(n_1077), .Y(n_1193) );
INVx2_ASAP7_75t_L g1194 ( .A(n_1156), .Y(n_1194) );
OR2x2_ASAP7_75t_L g1195 ( .A(n_1184), .B(n_1104), .Y(n_1195) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1176), .Y(n_1196) );
NAND2xp5_ASAP7_75t_L g1197 ( .A(n_1162), .B(n_1079), .Y(n_1197) );
NAND2x1p5_ASAP7_75t_L g1198 ( .A(n_1171), .B(n_1133), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1199 ( .A(n_1140), .B(n_1075), .Y(n_1199) );
AND3x2_ASAP7_75t_L g1200 ( .A(n_1189), .B(n_1107), .C(n_1131), .Y(n_1200) );
NAND2xp5_ASAP7_75t_L g1201 ( .A(n_1168), .B(n_1112), .Y(n_1201) );
NAND2xp5_ASAP7_75t_L g1202 ( .A(n_1161), .B(n_1163), .Y(n_1202) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1176), .Y(n_1203) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1180), .Y(n_1204) );
INVx2_ASAP7_75t_SL g1205 ( .A(n_1171), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1180), .Y(n_1206) );
INVx1_ASAP7_75t_SL g1207 ( .A(n_1191), .Y(n_1207) );
OR2x2_ASAP7_75t_L g1208 ( .A(n_1184), .B(n_1078), .Y(n_1208) );
CKINVDCx16_ASAP7_75t_R g1209 ( .A(n_1149), .Y(n_1209) );
INVxp67_ASAP7_75t_L g1210 ( .A(n_1149), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1141), .B(n_1130), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1212 ( .A(n_1161), .B(n_1132), .Y(n_1212) );
NOR2xp33_ASAP7_75t_L g1213 ( .A(n_1165), .B(n_1109), .Y(n_1213) );
NAND2xp5_ASAP7_75t_L g1214 ( .A(n_1163), .B(n_1108), .Y(n_1214) );
OAI22xp5_ASAP7_75t_SL g1215 ( .A1(n_1146), .A2(n_1083), .B1(n_1125), .B2(n_1099), .Y(n_1215) );
NAND2xp5_ASAP7_75t_L g1216 ( .A(n_1186), .B(n_1108), .Y(n_1216) );
AND2x4_ASAP7_75t_L g1217 ( .A(n_1146), .B(n_1139), .Y(n_1217) );
INVx1_ASAP7_75t_SL g1218 ( .A(n_1185), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1219 ( .A(n_1186), .B(n_1106), .Y(n_1219) );
OR2x2_ASAP7_75t_L g1220 ( .A(n_1169), .B(n_1164), .Y(n_1220) );
HB1xp67_ASAP7_75t_L g1221 ( .A(n_1157), .Y(n_1221) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1150), .Y(n_1222) );
NAND2xp5_ASAP7_75t_L g1223 ( .A(n_1145), .B(n_1106), .Y(n_1223) );
NAND2xp5_ASAP7_75t_L g1224 ( .A(n_1155), .B(n_1085), .Y(n_1224) );
INVx2_ASAP7_75t_L g1225 ( .A(n_1156), .Y(n_1225) );
AND2x2_ASAP7_75t_L g1226 ( .A(n_1141), .B(n_1130), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1142), .B(n_1114), .Y(n_1227) );
HB1xp67_ASAP7_75t_L g1228 ( .A(n_1174), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1229 ( .A(n_1190), .B(n_1085), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1230 ( .A(n_1142), .B(n_1114), .Y(n_1230) );
NAND2xp5_ASAP7_75t_L g1231 ( .A(n_1190), .B(n_1090), .Y(n_1231) );
INVx3_ASAP7_75t_L g1232 ( .A(n_1187), .Y(n_1232) );
INVx1_ASAP7_75t_SL g1233 ( .A(n_1187), .Y(n_1233) );
AOI222xp33_ASAP7_75t_L g1234 ( .A1(n_1215), .A2(n_1188), .B1(n_1083), .B2(n_1143), .C1(n_1144), .C2(n_1179), .Y(n_1234) );
OR2x2_ASAP7_75t_L g1235 ( .A(n_1220), .B(n_1169), .Y(n_1235) );
INVx1_ASAP7_75t_SL g1236 ( .A(n_1207), .Y(n_1236) );
AOI21xp5_ASAP7_75t_L g1237 ( .A1(n_1215), .A2(n_1181), .B(n_1182), .Y(n_1237) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1196), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1196), .Y(n_1239) );
AOI22xp33_ASAP7_75t_L g1240 ( .A1(n_1213), .A2(n_1183), .B1(n_1175), .B2(n_1146), .Y(n_1240) );
NOR2xp33_ASAP7_75t_L g1241 ( .A(n_1221), .B(n_1167), .Y(n_1241) );
NAND2xp5_ASAP7_75t_L g1242 ( .A(n_1227), .B(n_1174), .Y(n_1242) );
NAND2xp5_ASAP7_75t_L g1243 ( .A(n_1227), .B(n_1154), .Y(n_1243) );
XNOR2x2_ASAP7_75t_L g1244 ( .A(n_1218), .B(n_1148), .Y(n_1244) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1202), .Y(n_1245) );
OR2x2_ASAP7_75t_L g1246 ( .A(n_1220), .B(n_1154), .Y(n_1246) );
OAI221xp5_ASAP7_75t_SL g1247 ( .A1(n_1210), .A2(n_1151), .B1(n_1147), .B2(n_1148), .C(n_1143), .Y(n_1247) );
NAND3xp33_ASAP7_75t_L g1248 ( .A(n_1209), .B(n_1087), .C(n_1089), .Y(n_1248) );
OAI22xp5_ASAP7_75t_L g1249 ( .A1(n_1209), .A2(n_1151), .B1(n_1147), .B2(n_1119), .Y(n_1249) );
AO21x1_ASAP7_75t_L g1250 ( .A1(n_1224), .A2(n_1129), .B(n_1158), .Y(n_1250) );
INVx2_ASAP7_75t_L g1251 ( .A(n_1194), .Y(n_1251) );
AOI21xp33_ASAP7_75t_L g1252 ( .A1(n_1201), .A2(n_1119), .B(n_1125), .Y(n_1252) );
NAND2xp5_ASAP7_75t_L g1253 ( .A(n_1230), .B(n_1199), .Y(n_1253) );
NAND2xp5_ASAP7_75t_L g1254 ( .A(n_1230), .B(n_1144), .Y(n_1254) );
NAND2xp5_ASAP7_75t_L g1255 ( .A(n_1199), .B(n_1170), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_1192), .B(n_1211), .Y(n_1256) );
OAI21xp5_ASAP7_75t_SL g1257 ( .A1(n_1200), .A2(n_1153), .B(n_1187), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1192), .B(n_1159), .Y(n_1258) );
INVx2_ASAP7_75t_L g1259 ( .A(n_1194), .Y(n_1259) );
OAI21xp5_ASAP7_75t_L g1260 ( .A1(n_1218), .A2(n_1160), .B(n_1172), .Y(n_1260) );
NOR2xp33_ASAP7_75t_L g1261 ( .A(n_1193), .B(n_1166), .Y(n_1261) );
INVxp67_ASAP7_75t_L g1262 ( .A(n_1205), .Y(n_1262) );
INVx2_ASAP7_75t_L g1263 ( .A(n_1225), .Y(n_1263) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1235), .Y(n_1264) );
OAI221xp5_ASAP7_75t_L g1265 ( .A1(n_1240), .A2(n_1212), .B1(n_1198), .B2(n_1197), .C(n_1205), .Y(n_1265) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_1245), .B(n_1226), .Y(n_1266) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1235), .Y(n_1267) );
NAND2xp5_ASAP7_75t_L g1268 ( .A(n_1253), .B(n_1226), .Y(n_1268) );
XOR2x2_ASAP7_75t_L g1269 ( .A(n_1236), .B(n_1198), .Y(n_1269) );
OAI22xp5_ASAP7_75t_L g1270 ( .A1(n_1247), .A2(n_1198), .B1(n_1195), .B2(n_1208), .Y(n_1270) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1246), .Y(n_1271) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1246), .Y(n_1272) );
XNOR2x1_ASAP7_75t_L g1273 ( .A(n_1244), .B(n_1195), .Y(n_1273) );
O2A1O1Ixp5_ASAP7_75t_L g1274 ( .A1(n_1250), .A2(n_1232), .B(n_1217), .C(n_1229), .Y(n_1274) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1238), .Y(n_1275) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1238), .Y(n_1276) );
A2O1A1Ixp33_ASAP7_75t_L g1277 ( .A1(n_1237), .A2(n_1232), .B(n_1217), .C(n_1233), .Y(n_1277) );
OAI21xp5_ASAP7_75t_SL g1278 ( .A1(n_1257), .A2(n_1233), .B(n_1232), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1256), .B(n_1211), .Y(n_1279) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1239), .Y(n_1280) );
OR2x2_ASAP7_75t_L g1281 ( .A(n_1242), .B(n_1228), .Y(n_1281) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1239), .Y(n_1282) );
NAND2xp5_ASAP7_75t_SL g1283 ( .A(n_1250), .B(n_1217), .Y(n_1283) );
AOI22xp5_ASAP7_75t_L g1284 ( .A1(n_1273), .A2(n_1234), .B1(n_1261), .B2(n_1241), .Y(n_1284) );
AOI21xp33_ASAP7_75t_L g1285 ( .A1(n_1265), .A2(n_1248), .B(n_1262), .Y(n_1285) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1273), .B(n_1256), .Y(n_1286) );
INVxp67_ASAP7_75t_L g1287 ( .A(n_1269), .Y(n_1287) );
INVx2_ASAP7_75t_SL g1288 ( .A(n_1281), .Y(n_1288) );
O2A1O1Ixp33_ASAP7_75t_SL g1289 ( .A1(n_1277), .A2(n_1260), .B(n_1249), .C(n_1244), .Y(n_1289) );
OAI32xp33_ASAP7_75t_L g1290 ( .A1(n_1283), .A2(n_1254), .A3(n_1255), .B1(n_1243), .B2(n_1208), .Y(n_1290) );
AOI221xp5_ASAP7_75t_L g1291 ( .A1(n_1270), .A2(n_1252), .B1(n_1231), .B2(n_1216), .C(n_1219), .Y(n_1291) );
OA21x2_ASAP7_75t_SL g1292 ( .A1(n_1283), .A2(n_1217), .B(n_1223), .Y(n_1292) );
NAND2xp5_ASAP7_75t_L g1293 ( .A(n_1264), .B(n_1258), .Y(n_1293) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1275), .Y(n_1294) );
AOI22x1_ASAP7_75t_L g1295 ( .A1(n_1278), .A2(n_1177), .B1(n_1258), .B2(n_1129), .Y(n_1295) );
NAND2xp5_ASAP7_75t_L g1296 ( .A(n_1267), .B(n_1214), .Y(n_1296) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1294), .Y(n_1297) );
AOI221xp5_ASAP7_75t_L g1298 ( .A1(n_1289), .A2(n_1277), .B1(n_1274), .B2(n_1272), .C(n_1271), .Y(n_1298) );
NAND3xp33_ASAP7_75t_L g1299 ( .A(n_1287), .B(n_1274), .C(n_1280), .Y(n_1299) );
OAI21xp5_ASAP7_75t_L g1300 ( .A1(n_1284), .A2(n_1279), .B(n_1266), .Y(n_1300) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1293), .Y(n_1301) );
AO22x1_ASAP7_75t_L g1302 ( .A1(n_1292), .A2(n_1268), .B1(n_1276), .B2(n_1282), .Y(n_1302) );
AND2x4_ASAP7_75t_L g1303 ( .A(n_1288), .B(n_1263), .Y(n_1303) );
HB1xp67_ASAP7_75t_L g1304 ( .A(n_1296), .Y(n_1304) );
AOI221xp5_ASAP7_75t_L g1305 ( .A1(n_1290), .A2(n_1206), .B1(n_1203), .B2(n_1204), .C(n_1222), .Y(n_1305) );
NAND4xp75_ASAP7_75t_L g1306 ( .A(n_1298), .B(n_1291), .C(n_1286), .D(n_1285), .Y(n_1306) );
NOR3xp33_ASAP7_75t_L g1307 ( .A(n_1302), .B(n_1285), .C(n_1263), .Y(n_1307) );
OAI211xp5_ASAP7_75t_SL g1308 ( .A1(n_1300), .A2(n_1295), .B(n_1089), .C(n_1087), .Y(n_1308) );
NOR2xp33_ASAP7_75t_L g1309 ( .A(n_1304), .B(n_1259), .Y(n_1309) );
AND2x4_ASAP7_75t_L g1310 ( .A(n_1303), .B(n_1173), .Y(n_1310) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1297), .Y(n_1311) );
OAI222xp33_ASAP7_75t_L g1312 ( .A1(n_1306), .A2(n_1301), .B1(n_1303), .B2(n_1299), .C1(n_1305), .C2(n_1251), .Y(n_1312) );
OR2x2_ASAP7_75t_L g1313 ( .A(n_1311), .B(n_1259), .Y(n_1313) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1309), .Y(n_1314) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1310), .Y(n_1315) );
HB1xp67_ASAP7_75t_L g1316 ( .A(n_1314), .Y(n_1316) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1313), .Y(n_1317) );
XNOR2xp5_ASAP7_75t_L g1318 ( .A(n_1315), .B(n_1307), .Y(n_1318) );
NAND2xp5_ASAP7_75t_L g1319 ( .A(n_1318), .B(n_1251), .Y(n_1319) );
OAI22xp5_ASAP7_75t_SL g1320 ( .A1(n_1316), .A2(n_1312), .B1(n_1308), .B2(n_1138), .Y(n_1320) );
INVxp67_ASAP7_75t_L g1321 ( .A(n_1319), .Y(n_1321) );
AND3x4_ASAP7_75t_L g1322 ( .A(n_1320), .B(n_1316), .C(n_1317), .Y(n_1322) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1321), .Y(n_1323) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1323), .Y(n_1324) );
AOI22xp33_ASAP7_75t_SL g1325 ( .A1(n_1324), .A2(n_1322), .B1(n_1152), .B2(n_1166), .Y(n_1325) );
endmodule