module real_aes_4846_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_469;
wire n_987;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_974;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_983;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_961;
wire n_271;
wire n_489;
wire n_548;
wire n_678;
wire n_427;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_994;
wire n_528;
wire n_202;
wire n_578;
wire n_495;
wire n_892;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_106;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_984;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_931;
wire n_904;
wire n_174;
wire n_780;
wire n_570;
wire n_675;
wire n_840;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_962;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_656;
wire n_316;
wire n_532;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_996;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_164;
wire n_671;
wire n_973;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_985;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_957;
wire n_995;
wire n_296;
wire n_702;
wire n_954;
wire n_969;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_997;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_649;
wire n_397;
wire n_162;
wire n_293;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_965;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_720;
wire n_265;
wire n_354;
wire n_972;
wire n_968;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_653;
wire n_290;
wire n_365;
wire n_637;
wire n_526;
wire n_155;
wire n_928;
wire n_243;
wire n_899;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_679;
wire n_520;
wire n_922;
wire n_926;
wire n_149;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_134;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_982;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
OAI21xp5_ASAP7_75t_L g105 ( .A1(n_0), .A2(n_106), .B(n_564), .Y(n_105) );
INVx1_ASAP7_75t_L g566 ( .A(n_0), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_1), .B(n_292), .Y(n_622) );
CKINVDCx5p33_ASAP7_75t_R g636 ( .A(n_2), .Y(n_636) );
INVx1_ASAP7_75t_L g255 ( .A(n_3), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_4), .A2(n_94), .B1(n_582), .B2(n_583), .Y(n_581) );
INVx1_ASAP7_75t_L g583 ( .A(n_4), .Y(n_583) );
O2A1O1Ixp33_ASAP7_75t_SL g670 ( .A1(n_5), .A2(n_172), .B(n_671), .C(n_672), .Y(n_670) );
OAI22xp33_ASAP7_75t_L g627 ( .A1(n_6), .A2(n_84), .B1(n_143), .B2(n_164), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_7), .B(n_142), .Y(n_213) );
INVxp67_ASAP7_75t_L g110 ( .A(n_8), .Y(n_110) );
INVx1_ASAP7_75t_L g593 ( .A(n_8), .Y(n_593) );
INVx1_ASAP7_75t_L g969 ( .A(n_8), .Y(n_969) );
BUFx2_ASAP7_75t_L g996 ( .A(n_8), .Y(n_996) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_9), .B(n_215), .Y(n_214) );
AOI22xp33_ASAP7_75t_L g147 ( .A1(n_10), .A2(n_39), .B1(n_141), .B2(n_148), .Y(n_147) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_11), .A2(n_44), .B1(n_185), .B2(n_189), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g270 ( .A1(n_12), .A2(n_66), .B1(n_193), .B2(n_263), .Y(n_270) );
INVx1_ASAP7_75t_L g249 ( .A(n_13), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g654 ( .A(n_14), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_15), .A2(n_74), .B1(n_164), .B2(n_187), .Y(n_689) );
CKINVDCx5p33_ASAP7_75t_R g716 ( .A(n_16), .Y(n_716) );
INVx1_ASAP7_75t_L g253 ( .A(n_17), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_18), .A2(n_64), .B1(n_143), .B2(n_168), .Y(n_688) );
OA21x2_ASAP7_75t_L g131 ( .A1(n_19), .A2(n_73), .B(n_132), .Y(n_131) );
OA21x2_ASAP7_75t_L g175 ( .A1(n_19), .A2(n_73), .B(n_132), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g262 ( .A1(n_20), .A2(n_70), .B1(n_193), .B2(n_263), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_21), .A2(n_104), .B1(n_987), .B2(n_997), .Y(n_103) );
INVx1_ASAP7_75t_L g246 ( .A(n_22), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_23), .Y(n_588) );
CKINVDCx5p33_ASAP7_75t_R g649 ( .A(n_24), .Y(n_649) );
BUFx3_ASAP7_75t_L g576 ( .A(n_25), .Y(n_576) );
O2A1O1Ixp33_ASAP7_75t_L g676 ( .A1(n_26), .A2(n_269), .B(n_677), .C(n_678), .Y(n_676) );
OAI22xp33_ASAP7_75t_SL g625 ( .A1(n_27), .A2(n_48), .B1(n_139), .B2(n_143), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_28), .A2(n_37), .B1(n_139), .B2(n_211), .Y(n_615) );
AO22x1_ASAP7_75t_L g208 ( .A1(n_29), .A2(n_80), .B1(n_170), .B2(n_209), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_30), .Y(n_160) );
AND2x2_ASAP7_75t_L g280 ( .A(n_31), .B(n_189), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_32), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_33), .B(n_170), .Y(n_169) );
O2A1O1Ixp5_ASAP7_75t_L g697 ( .A1(n_34), .A2(n_172), .B(n_698), .C(n_699), .Y(n_697) );
INVx1_ASAP7_75t_L g115 ( .A(n_35), .Y(n_115) );
AOI22x1_ASAP7_75t_L g192 ( .A1(n_36), .A2(n_98), .B1(n_137), .B2(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_38), .B(n_152), .Y(n_151) );
AND2x2_ASAP7_75t_L g994 ( .A(n_40), .B(n_995), .Y(n_994) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_41), .B(n_619), .Y(n_618) );
CKINVDCx5p33_ASAP7_75t_R g700 ( .A(n_42), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_43), .B(n_227), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g674 ( .A(n_45), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_46), .B(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_47), .B(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g132 ( .A(n_49), .Y(n_132) );
AND2x4_ASAP7_75t_L g134 ( .A(n_50), .B(n_135), .Y(n_134) );
AND2x4_ASAP7_75t_L g613 ( .A(n_50), .B(n_135), .Y(n_613) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_51), .Y(n_129) );
INVx2_ASAP7_75t_L g265 ( .A(n_52), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g634 ( .A(n_53), .Y(n_634) );
O2A1O1Ixp33_ASAP7_75t_L g651 ( .A1(n_54), .A2(n_172), .B(n_652), .C(n_653), .Y(n_651) );
CKINVDCx5p33_ASAP7_75t_R g705 ( .A(n_55), .Y(n_705) );
INVx2_ASAP7_75t_L g721 ( .A(n_56), .Y(n_721) );
CKINVDCx5p33_ASAP7_75t_R g633 ( .A(n_57), .Y(n_633) );
INVx1_ASAP7_75t_L g560 ( .A(n_58), .Y(n_560) );
INVx1_ASAP7_75t_L g563 ( .A(n_58), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g136 ( .A1(n_59), .A2(n_76), .B1(n_137), .B2(n_141), .Y(n_136) );
CKINVDCx14_ASAP7_75t_R g218 ( .A(n_60), .Y(n_218) );
AND2x2_ASAP7_75t_L g285 ( .A(n_61), .B(n_170), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_62), .B(n_222), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_63), .A2(n_82), .B1(n_186), .B2(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_65), .B(n_233), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g637 ( .A(n_67), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_68), .B(n_222), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_69), .A2(n_581), .B1(n_584), .B2(n_585), .Y(n_580) );
BUFx4f_ASAP7_75t_SL g586 ( .A(n_69), .Y(n_586) );
NAND2xp33_ASAP7_75t_R g691 ( .A(n_71), .B(n_131), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_71), .A2(n_101), .B1(n_241), .B2(n_619), .Y(n_753) );
NAND2x1p5_ASAP7_75t_L g288 ( .A(n_72), .B(n_179), .Y(n_288) );
CKINVDCx14_ASAP7_75t_R g197 ( .A(n_75), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_77), .B(n_142), .Y(n_228) );
OR2x6_ASAP7_75t_L g112 ( .A(n_78), .B(n_113), .Y(n_112) );
AND3x1_ASAP7_75t_L g993 ( .A(n_78), .B(n_994), .C(n_996), .Y(n_993) );
CKINVDCx5p33_ASAP7_75t_R g720 ( .A(n_79), .Y(n_720) );
CKINVDCx5p33_ASAP7_75t_R g717 ( .A(n_81), .Y(n_717) );
INVx1_ASAP7_75t_L g114 ( .A(n_83), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_83), .B(n_115), .Y(n_992) );
INVx1_ASAP7_75t_L g995 ( .A(n_85), .Y(n_995) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_86), .Y(n_140) );
BUFx5_ASAP7_75t_L g143 ( .A(n_86), .Y(n_143) );
INVx1_ASAP7_75t_L g188 ( .A(n_86), .Y(n_188) );
INVxp33_ASAP7_75t_SL g559 ( .A(n_87), .Y(n_559) );
CKINVDCx5p33_ASAP7_75t_R g561 ( .A(n_87), .Y(n_561) );
INVx2_ASAP7_75t_L g683 ( .A(n_88), .Y(n_683) );
INVx2_ASAP7_75t_L g257 ( .A(n_89), .Y(n_257) );
INVx2_ASAP7_75t_L g656 ( .A(n_90), .Y(n_656) );
CKINVDCx5p33_ASAP7_75t_R g679 ( .A(n_91), .Y(n_679) );
NAND2xp33_ASAP7_75t_L g282 ( .A(n_92), .B(n_138), .Y(n_282) );
INVx2_ASAP7_75t_SL g135 ( .A(n_93), .Y(n_135) );
INVx1_ASAP7_75t_L g582 ( .A(n_94), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_95), .B(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_96), .B(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g703 ( .A(n_97), .Y(n_703) );
INVx2_ASAP7_75t_L g708 ( .A(n_99), .Y(n_708) );
OAI21xp33_ASAP7_75t_SL g647 ( .A1(n_100), .A2(n_143), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_101), .B(n_619), .Y(n_711) );
INVxp67_ASAP7_75t_SL g747 ( .A(n_101), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_102), .B(n_177), .Y(n_176) );
OA21x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_573), .B(n_577), .Y(n_104) );
NAND2x1p5_ASAP7_75t_L g106 ( .A(n_107), .B(n_116), .Y(n_106) );
BUFx12f_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_108), .Y(n_568) );
INVx3_ASAP7_75t_L g572 ( .A(n_108), .Y(n_572) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
OR2x6_ASAP7_75t_L g968 ( .A(n_111), .B(n_969), .Y(n_968) );
INVx8_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OR2x6_ASAP7_75t_L g592 ( .A(n_112), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g599 ( .A(n_112), .B(n_593), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI21xp33_ASAP7_75t_L g564 ( .A1(n_117), .A2(n_565), .B(n_569), .Y(n_564) );
XNOR2x1_ASAP7_75t_L g117 ( .A(n_118), .B(n_557), .Y(n_117) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_118), .A2(n_596), .B1(n_600), .B2(n_966), .Y(n_595) );
AND2x4_ASAP7_75t_L g971 ( .A(n_118), .B(n_972), .Y(n_971) );
AND2x4_ASAP7_75t_L g118 ( .A(n_119), .B(n_450), .Y(n_118) );
NOR3xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_362), .C(n_398), .Y(n_119) );
NAND3xp33_ASAP7_75t_SL g120 ( .A(n_121), .B(n_295), .C(n_340), .Y(n_120) );
AOI22xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_199), .B1(n_271), .B2(n_274), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g553 ( .A(n_123), .Y(n_553) );
OR2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_154), .Y(n_123) );
INVx2_ASAP7_75t_L g315 ( .A(n_124), .Y(n_315) );
INVx2_ASAP7_75t_L g442 ( .A(n_124), .Y(n_442) );
INVx2_ASAP7_75t_SL g124 ( .A(n_125), .Y(n_124) );
AND2x2_ASAP7_75t_L g294 ( .A(n_125), .B(n_155), .Y(n_294) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_144), .Y(n_125) );
NAND2x1p5_ASAP7_75t_L g310 ( .A(n_126), .B(n_144), .Y(n_310) );
OR2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_136), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_130), .Y(n_127) );
OAI22xp5_ASAP7_75t_L g157 ( .A1(n_128), .A2(n_141), .B1(n_158), .B2(n_162), .Y(n_157) );
INVx4_ASAP7_75t_L g161 ( .A(n_128), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_128), .A2(n_226), .B(n_228), .Y(n_225) );
OA22x2_ASAP7_75t_L g614 ( .A1(n_128), .A2(n_146), .B1(n_615), .B2(n_616), .Y(n_614) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g146 ( .A(n_129), .Y(n_146) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_129), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_129), .B(n_246), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_129), .B(n_249), .Y(n_248) );
INVx4_ASAP7_75t_L g252 ( .A(n_129), .Y(n_252) );
INVx3_ASAP7_75t_L g269 ( .A(n_129), .Y(n_269) );
INVxp67_ASAP7_75t_L g283 ( .A(n_129), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_129), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_129), .B(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_130), .B(n_146), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_133), .Y(n_130) );
INVx1_ASAP7_75t_L g153 ( .A(n_131), .Y(n_153) );
INVx2_ASAP7_75t_L g242 ( .A(n_131), .Y(n_242) );
BUFx3_ASAP7_75t_L g612 ( .A(n_131), .Y(n_612) );
INVx1_ASAP7_75t_L g645 ( .A(n_131), .Y(n_645) );
INVx1_ASAP7_75t_L g709 ( .A(n_131), .Y(n_709) );
INVx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_134), .Y(n_173) );
INVx1_ASAP7_75t_L g205 ( .A(n_134), .Y(n_205) );
INVx3_ASAP7_75t_L g236 ( .A(n_134), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_134), .B(n_180), .Y(n_628) );
OAI221xp5_ASAP7_75t_L g631 ( .A1(n_134), .A2(n_172), .B1(n_269), .B2(n_632), .C(n_635), .Y(n_631) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g190 ( .A(n_139), .Y(n_190) );
INVx1_ASAP7_75t_L g227 ( .A(n_139), .Y(n_227) );
INVx2_ASAP7_75t_SL g617 ( .A(n_139), .Y(n_617) );
AOI22xp33_ASAP7_75t_SL g632 ( .A1(n_139), .A2(n_143), .B1(n_633), .B2(n_634), .Y(n_632) );
INVx2_ASAP7_75t_L g673 ( .A(n_139), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_139), .A2(n_143), .B1(n_716), .B2(n_717), .Y(n_715) );
INVx6_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx3_ASAP7_75t_L g150 ( .A(n_140), .Y(n_150) );
INVx2_ASAP7_75t_L g164 ( .A(n_140), .Y(n_164) );
INVx2_ASAP7_75t_L g168 ( .A(n_140), .Y(n_168) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g170 ( .A(n_143), .Y(n_170) );
INVx2_ASAP7_75t_L g194 ( .A(n_143), .Y(n_194) );
INVx2_ASAP7_75t_L g233 ( .A(n_143), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_143), .A2(n_168), .B1(n_636), .B2(n_637), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g648 ( .A(n_143), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_143), .B(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_143), .B(n_705), .Y(n_704) );
OA21x2_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_147), .B(n_151), .Y(n_144) );
INVx1_ASAP7_75t_L g191 ( .A(n_146), .Y(n_191) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g263 ( .A(n_149), .Y(n_263) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g215 ( .A(n_150), .Y(n_215) );
INVx2_ASAP7_75t_L g231 ( .A(n_150), .Y(n_231) );
INVx1_ASAP7_75t_L g652 ( .A(n_150), .Y(n_652) );
INVx1_ASAP7_75t_L g698 ( .A(n_150), .Y(n_698) );
INVx1_ASAP7_75t_L g195 ( .A(n_152), .Y(n_195) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
OR2x2_ASAP7_75t_L g390 ( .A(n_154), .B(n_391), .Y(n_390) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_154), .Y(n_538) );
NAND2x1_ASAP7_75t_L g154 ( .A(n_155), .B(n_181), .Y(n_154) );
AND2x2_ASAP7_75t_L g336 ( .A(n_155), .B(n_310), .Y(n_336) );
AND2x2_ASAP7_75t_L g482 ( .A(n_155), .B(n_318), .Y(n_482) );
OA21x2_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_174), .B(n_176), .Y(n_155) );
OA21x2_ASAP7_75t_L g312 ( .A1(n_156), .A2(n_174), .B(n_176), .Y(n_312) );
OAI21x1_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_165), .B(n_173), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_159), .B(n_161), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
OAI22x1_ASAP7_75t_L g183 ( .A1(n_161), .A2(n_184), .B1(n_191), .B2(n_192), .Y(n_183) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_169), .B(n_171), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_167), .B(n_248), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_167), .A2(n_170), .B1(n_251), .B2(n_254), .Y(n_250) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g677 ( .A(n_168), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_168), .A2(n_211), .B1(n_720), .B2(n_721), .Y(n_719) );
INVxp67_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g207 ( .A(n_172), .Y(n_207) );
INVx2_ASAP7_75t_SL g216 ( .A(n_172), .Y(n_216) );
INVx1_ASAP7_75t_L g234 ( .A(n_172), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_172), .A2(n_252), .B1(n_688), .B2(n_689), .Y(n_687) );
OAI22xp33_ASAP7_75t_L g745 ( .A1(n_172), .A2(n_252), .B1(n_715), .B2(n_719), .Y(n_745) );
AO31x2_ASAP7_75t_L g182 ( .A1(n_173), .A2(n_183), .A3(n_195), .B(n_196), .Y(n_182) );
AO31x2_ASAP7_75t_L g276 ( .A1(n_173), .A2(n_183), .A3(n_195), .B(n_196), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_173), .B(n_611), .Y(n_744) );
INVx3_ASAP7_75t_L g198 ( .A(n_174), .Y(n_198) );
BUFx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx4_ASAP7_75t_L g180 ( .A(n_175), .Y(n_180) );
INVx2_ASAP7_75t_L g223 ( .A(n_175), .Y(n_223) );
OR2x2_ASAP7_75t_L g204 ( .A(n_177), .B(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
OR2x2_ASAP7_75t_L g264 ( .A(n_178), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g292 ( .A(n_180), .Y(n_292) );
INVx2_ASAP7_75t_L g619 ( .A(n_180), .Y(n_619) );
NOR2xp33_ASAP7_75t_SL g682 ( .A(n_180), .B(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g308 ( .A(n_181), .Y(n_308) );
INVx1_ASAP7_75t_L g327 ( .A(n_181), .Y(n_327) );
AND2x2_ASAP7_75t_L g335 ( .A(n_181), .B(n_278), .Y(n_335) );
AND2x2_ASAP7_75t_L g471 ( .A(n_181), .B(n_351), .Y(n_471) );
INVx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g343 ( .A(n_182), .B(n_311), .Y(n_343) );
INVx3_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g671 ( .A(n_186), .Y(n_671) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g211 ( .A(n_188), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_189), .B(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NOR2xp67_ASAP7_75t_SL g196 ( .A(n_197), .B(n_198), .Y(n_196) );
OR2x2_ASAP7_75t_L g217 ( .A(n_198), .B(n_218), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g726 ( .A1(n_198), .A2(n_727), .B(n_728), .Y(n_726) );
INVx2_ASAP7_75t_SL g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g547 ( .A(n_200), .Y(n_547) );
OR2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_237), .Y(n_200) );
OR2x2_ASAP7_75t_L g401 ( .A(n_201), .B(n_321), .Y(n_401) );
OR2x2_ASAP7_75t_SL g511 ( .A(n_201), .B(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g271 ( .A(n_202), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g455 ( .A(n_202), .B(n_414), .Y(n_455) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_219), .Y(n_202) );
INVx2_ASAP7_75t_SL g333 ( .A(n_203), .Y(n_333) );
AND2x2_ASAP7_75t_L g339 ( .A(n_203), .B(n_220), .Y(n_339) );
OAI21x1_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_206), .B(n_217), .Y(n_203) );
OAI21xp5_ASAP7_75t_L g302 ( .A1(n_204), .A2(n_206), .B(n_217), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_205), .B(n_241), .Y(n_240) );
NOR2xp67_ASAP7_75t_L g690 ( .A(n_205), .B(n_222), .Y(n_690) );
AOI21x1_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B(n_212), .Y(n_206) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_211), .B(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_211), .B(n_679), .Y(n_678) );
AOI21x1_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_216), .Y(n_212) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_215), .A2(n_252), .B1(n_702), .B2(n_704), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_216), .B(n_288), .Y(n_289) );
INVx1_ASAP7_75t_L g377 ( .A(n_219), .Y(n_377) );
AND2x2_ASAP7_75t_L g461 ( .A(n_219), .B(n_258), .Y(n_461) );
INVx3_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g299 ( .A(n_220), .Y(n_299) );
AND2x2_ASAP7_75t_L g332 ( .A(n_220), .B(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g220 ( .A(n_221), .B(n_224), .Y(n_220) );
NOR2x1_ASAP7_75t_L g235 ( .A(n_222), .B(n_236), .Y(n_235) );
INVx3_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_223), .B(n_257), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_223), .B(n_656), .Y(n_655) );
BUFx3_ASAP7_75t_L g706 ( .A(n_223), .Y(n_706) );
OAI21x1_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_229), .B(n_235), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_232), .B(n_234), .Y(n_229) );
AOI221xp5_ASAP7_75t_L g713 ( .A1(n_234), .A2(n_650), .B1(n_681), .B2(n_714), .C(n_718), .Y(n_713) );
INVx2_ASAP7_75t_L g261 ( .A(n_236), .Y(n_261) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g338 ( .A(n_238), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_238), .B(n_439), .Y(n_438) );
NAND2x1_ASAP7_75t_SL g476 ( .A(n_238), .B(n_332), .Y(n_476) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_238), .Y(n_487) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_258), .Y(n_238) );
INVx1_ASAP7_75t_L g273 ( .A(n_239), .Y(n_273) );
INVxp67_ASAP7_75t_L g298 ( .A(n_239), .Y(n_298) );
OR2x2_ASAP7_75t_L g323 ( .A(n_239), .B(n_302), .Y(n_323) );
INVx1_ASAP7_75t_L g385 ( .A(n_239), .Y(n_385) );
INVx1_ASAP7_75t_L g397 ( .A(n_239), .Y(n_397) );
AND2x2_ASAP7_75t_L g432 ( .A(n_239), .B(n_333), .Y(n_432) );
AO21x2_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_243), .B(n_256), .Y(n_239) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NAND3xp33_ASAP7_75t_SL g260 ( .A(n_242), .B(n_252), .C(n_261), .Y(n_260) );
NAND3xp33_ASAP7_75t_L g267 ( .A(n_242), .B(n_261), .C(n_268), .Y(n_267) );
NAND3xp33_ASAP7_75t_SL g243 ( .A(n_244), .B(n_247), .C(n_250), .Y(n_243) );
NOR2xp33_ASAP7_75t_SL g251 ( .A(n_252), .B(n_253), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_252), .B(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g650 ( .A(n_252), .Y(n_650) );
AND2x2_ASAP7_75t_L g272 ( .A(n_258), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g303 ( .A(n_258), .Y(n_303) );
INVx1_ASAP7_75t_L g321 ( .A(n_258), .Y(n_321) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_258), .Y(n_366) );
NOR2x1_ASAP7_75t_L g396 ( .A(n_258), .B(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g415 ( .A(n_258), .Y(n_415) );
INVx1_ASAP7_75t_L g418 ( .A(n_258), .Y(n_418) );
OR2x6_ASAP7_75t_L g258 ( .A(n_259), .B(n_266), .Y(n_258) );
OAI21x1_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_262), .B(n_264), .Y(n_259) );
AOI21xp33_ASAP7_75t_SL g290 ( .A1(n_261), .A2(n_291), .B(n_293), .Y(n_290) );
NOR2xp67_ASAP7_75t_L g266 ( .A(n_267), .B(n_270), .Y(n_266) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g626 ( .A1(n_269), .A2(n_627), .B(n_628), .Y(n_626) );
AND2x2_ASAP7_75t_L g414 ( .A(n_273), .B(n_415), .Y(n_414) );
AND2x4_ASAP7_75t_L g274 ( .A(n_275), .B(n_294), .Y(n_274) );
BUFx3_ASAP7_75t_L g345 ( .A(n_275), .Y(n_345) );
INVx3_ASAP7_75t_L g443 ( .A(n_275), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_275), .B(n_349), .Y(n_543) );
AND2x4_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
OR2x2_ASAP7_75t_L g317 ( .A(n_276), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g361 ( .A(n_276), .B(n_318), .Y(n_361) );
INVx1_ASAP7_75t_L g447 ( .A(n_276), .Y(n_447) );
INVx1_ASAP7_75t_L g437 ( .A(n_277), .Y(n_437) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVxp67_ASAP7_75t_L g348 ( .A(n_278), .Y(n_348) );
INVx1_ASAP7_75t_L g429 ( .A(n_278), .Y(n_429) );
AO21x2_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_284), .B(n_290), .Y(n_278) );
AO21x2_ASAP7_75t_L g318 ( .A1(n_279), .A2(n_284), .B(n_290), .Y(n_318) );
OAI21x1_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_281), .B(n_283), .Y(n_279) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OAI21x1_ASAP7_75t_SL g284 ( .A1(n_285), .A2(n_286), .B(n_289), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx1_ASAP7_75t_L g293 ( .A(n_288), .Y(n_293) );
INVx2_ASAP7_75t_L g630 ( .A(n_291), .Y(n_630) );
OR2x2_ASAP7_75t_L g746 ( .A(n_291), .B(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_SL g680 ( .A(n_292), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g354 ( .A(n_294), .Y(n_354) );
AND2x2_ASAP7_75t_L g467 ( .A(n_294), .B(n_468), .Y(n_467) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_294), .Y(n_500) );
NOR2xp67_ASAP7_75t_SL g505 ( .A(n_294), .B(n_443), .Y(n_505) );
INVx1_ASAP7_75t_L g533 ( .A(n_294), .Y(n_533) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_304), .B1(n_313), .B2(n_319), .C(n_324), .Y(n_295) );
INVx2_ASAP7_75t_L g475 ( .A(n_296), .Y(n_475) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_300), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_298), .Y(n_387) );
AND2x2_ASAP7_75t_L g320 ( .A(n_299), .B(n_321), .Y(n_320) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_299), .Y(n_358) );
INVx2_ASAP7_75t_L g439 ( .A(n_299), .Y(n_439) );
OR2x2_ASAP7_75t_L g456 ( .A(n_299), .B(n_323), .Y(n_456) );
AND2x2_ASAP7_75t_L g539 ( .A(n_300), .B(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
BUFx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_303), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_303), .B(n_432), .Y(n_556) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
AND2x2_ASAP7_75t_L g373 ( .A(n_307), .B(n_328), .Y(n_373) );
INVx1_ASAP7_75t_L g479 ( .A(n_307), .Y(n_479) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g508 ( .A(n_308), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_309), .Y(n_509) );
INVx2_ASAP7_75t_L g551 ( .A(n_309), .Y(n_551) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx2_ASAP7_75t_L g351 ( .A(n_310), .Y(n_351) );
INVx1_ASAP7_75t_L g372 ( .A(n_310), .Y(n_372) );
INVx1_ASAP7_75t_L g406 ( .A(n_310), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_310), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g349 ( .A(n_311), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_311), .B(n_351), .Y(n_495) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g329 ( .A(n_312), .Y(n_329) );
OAI31xp33_ASAP7_75t_L g535 ( .A1(n_313), .A2(n_536), .A3(n_537), .B(n_539), .Y(n_535) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2x1_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
AND3x2_ASAP7_75t_L g347 ( .A(n_315), .B(n_348), .C(n_349), .Y(n_347) );
AND2x2_ASAP7_75t_L g360 ( .A(n_315), .B(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g368 ( .A(n_317), .B(n_349), .Y(n_368) );
INVx2_ASAP7_75t_L g468 ( .A(n_317), .Y(n_468) );
AND2x4_ASAP7_75t_L g328 ( .A(n_318), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g355 ( .A(n_319), .Y(n_355) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .Y(n_319) );
NAND2x2_ASAP7_75t_L g430 ( .A(n_320), .B(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g331 ( .A(n_321), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g357 ( .A(n_322), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g367 ( .A(n_323), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_330), .B1(n_334), .B2(n_337), .Y(n_324) );
INVx2_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
NAND2xp67_ASAP7_75t_L g403 ( .A(n_326), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g409 ( .A(n_326), .Y(n_409) );
AND2x4_ASAP7_75t_SL g326 ( .A(n_327), .B(n_328), .Y(n_326) );
INVx1_ASAP7_75t_L g424 ( .A(n_327), .Y(n_424) );
AND2x2_ASAP7_75t_L g530 ( .A(n_327), .B(n_336), .Y(n_530) );
AND2x2_ASAP7_75t_L g350 ( .A(n_328), .B(n_351), .Y(n_350) );
BUFx3_ASAP7_75t_L g384 ( .A(n_328), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_328), .B(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_329), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AOI221xp5_ASAP7_75t_L g452 ( .A1(n_331), .A2(n_350), .B1(n_453), .B2(n_457), .C(n_458), .Y(n_452) );
INVx1_ASAP7_75t_L g378 ( .A(n_333), .Y(n_378) );
INVx1_ASAP7_75t_L g518 ( .A(n_333), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
AND2x2_ASAP7_75t_L g419 ( .A(n_336), .B(n_348), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_336), .B(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_338), .Y(n_352) );
INVx2_ASAP7_75t_L g393 ( .A(n_339), .Y(n_393) );
AND2x2_ASAP7_75t_L g489 ( .A(n_339), .B(n_490), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_350), .B(n_352), .C(n_353), .Y(n_340) );
NAND3xp33_ASAP7_75t_SL g341 ( .A(n_342), .B(n_344), .C(n_346), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2x1p5_ASAP7_75t_L g435 ( .A(n_343), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g391 ( .A(n_348), .Y(n_391) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_348), .Y(n_502) );
OR2x2_ASAP7_75t_L g498 ( .A(n_349), .B(n_428), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_355), .B1(n_356), .B2(n_359), .Y(n_353) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g516 ( .A(n_358), .B(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g545 ( .A(n_361), .Y(n_545) );
OAI221xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_368), .B1(n_369), .B2(n_374), .C(n_379), .Y(n_362) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
AND2x2_ASAP7_75t_L g417 ( .A(n_367), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g462 ( .A(n_367), .Y(n_462) );
AOI21xp33_ASAP7_75t_L g513 ( .A1(n_368), .A2(n_514), .B(n_515), .Y(n_513) );
INVxp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_373), .Y(n_370) );
AND2x2_ASAP7_75t_L g380 ( .A(n_371), .B(n_381), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_371), .B(n_445), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g453 ( .A1(n_371), .A2(n_442), .B1(n_454), .B2(n_456), .Y(n_453) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g485 ( .A(n_375), .Y(n_485) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NOR2xp67_ASAP7_75t_SL g421 ( .A(n_376), .B(n_385), .Y(n_421) );
OR2x2_ASAP7_75t_L g448 ( .A(n_376), .B(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
INVx1_ASAP7_75t_L g381 ( .A(n_377), .Y(n_381) );
INVxp67_ASAP7_75t_SL g412 ( .A(n_378), .Y(n_412) );
A2O1A1Ixp33_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_382), .B(n_385), .C(n_386), .Y(n_379) );
INVx1_ASAP7_75t_L g527 ( .A(n_381), .Y(n_527) );
INVxp67_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_383), .B(n_459), .Y(n_458) );
OAI22xp33_ASAP7_75t_L g497 ( .A1(n_383), .A2(n_430), .B1(n_488), .B2(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g466 ( .A(n_385), .Y(n_466) );
AND2x2_ASAP7_75t_L g517 ( .A(n_385), .B(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g540 ( .A(n_385), .B(n_439), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B(n_394), .Y(n_386) );
INVx1_ASAP7_75t_L g490 ( .A(n_387), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_389), .B(n_392), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI221xp5_ASAP7_75t_L g463 ( .A1(n_393), .A2(n_464), .B1(n_469), .B2(n_472), .C(n_474), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_394), .B(n_439), .Y(n_529) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g473 ( .A(n_395), .B(n_439), .Y(n_473) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NAND3xp33_ASAP7_75t_SL g398 ( .A(n_399), .B(n_407), .C(n_420), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_402), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_404), .B(n_434), .Y(n_521) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AOI21x1_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_410), .B(n_416), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_419), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g541 ( .A1(n_417), .A2(n_542), .B1(n_544), .B2(n_547), .C(n_548), .Y(n_541) );
INVx2_ASAP7_75t_L g512 ( .A(n_418), .Y(n_512) );
AOI211xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_422), .B(n_425), .C(n_440), .Y(n_420) );
INVxp67_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_430), .B1(n_433), .B2(n_438), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx3_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_L g534 ( .A(n_432), .B(n_461), .Y(n_534) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AOI211xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_443), .B(n_444), .C(n_448), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g514 ( .A(n_442), .B(n_481), .Y(n_514) );
AND2x2_ASAP7_75t_L g536 ( .A(n_442), .B(n_482), .Y(n_536) );
INVx1_ASAP7_75t_L g457 ( .A(n_444), .Y(n_457) );
INVx2_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g496 ( .A(n_447), .Y(n_496) );
NOR2xp67_ASAP7_75t_L g450 ( .A(n_451), .B(n_503), .Y(n_450) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_463), .C(n_483), .Y(n_451) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_462), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_468), .B(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AOI21xp33_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B(n_477), .Y(n_474) );
NOR3xp33_ASAP7_75t_L g499 ( .A(n_475), .B(n_500), .C(n_501), .Y(n_499) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NOR3xp33_ASAP7_75t_L g483 ( .A(n_484), .B(n_497), .C(n_499), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B(n_488), .C(n_491), .Y(n_484) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_496), .Y(n_493) );
INVxp67_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NAND4xp25_ASAP7_75t_SL g503 ( .A(n_504), .B(n_519), .C(n_535), .D(n_541), .Y(n_503) );
O2A1O1Ixp33_ASAP7_75t_SL g504 ( .A1(n_505), .A2(n_506), .B(n_510), .C(n_513), .Y(n_504) );
INVxp67_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
OR2x2_ASAP7_75t_L g532 ( .A(n_508), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g525 ( .A(n_512), .Y(n_525) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AOI222xp33_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_522), .B1(n_528), .B2(n_530), .C1(n_531), .C2(n_534), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_523), .B(n_526), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g546 ( .A(n_530), .Y(n_546) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVxp67_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
INVxp67_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
AOI21xp33_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_552), .B(n_554), .Y(n_548) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AOI22xp5_ASAP7_75t_SL g557 ( .A1(n_558), .A2(n_560), .B1(n_561), .B2(n_562), .Y(n_557) );
CKINVDCx5p33_ASAP7_75t_R g558 ( .A(n_559), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_563), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVxp67_ASAP7_75t_SL g984 ( .A(n_569), .Y(n_984) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_572), .Y(n_571) );
BUFx8_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
CKINVDCx6p67_ASAP7_75t_R g575 ( .A(n_576), .Y(n_575) );
HB1xp67_ASAP7_75t_L g986 ( .A(n_576), .Y(n_986) );
NAND3xp33_ASAP7_75t_L g577 ( .A(n_578), .B(n_984), .C(n_985), .Y(n_577) );
AO22x1_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_594), .B1(n_970), .B2(n_975), .Y(n_578) );
NOR2xp33_ASAP7_75t_R g579 ( .A(n_580), .B(n_587), .Y(n_579) );
CKINVDCx20_ASAP7_75t_R g974 ( .A(n_580), .Y(n_974) );
INVx1_ASAP7_75t_L g584 ( .A(n_581), .Y(n_584) );
CKINVDCx20_ASAP7_75t_R g585 ( .A(n_586), .Y(n_585) );
NOR3xp33_ASAP7_75t_L g970 ( .A(n_587), .B(n_971), .C(n_974), .Y(n_970) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
BUFx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
BUFx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
BUFx3_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVxp67_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
BUFx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g973 ( .A(n_598), .Y(n_973) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g983 ( .A(n_601), .Y(n_983) );
NAND4xp75_ASAP7_75t_L g601 ( .A(n_602), .B(n_811), .C(n_906), .D(n_931), .Y(n_601) );
NOR2x1_ASAP7_75t_L g602 ( .A(n_603), .B(n_765), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_722), .Y(n_603) );
OAI21xp33_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_639), .B(n_665), .Y(n_604) );
INVx1_ASAP7_75t_L g915 ( .A(n_605), .Y(n_915) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_620), .Y(n_606) );
AND2x2_ASAP7_75t_L g778 ( .A(n_607), .B(n_779), .Y(n_778) );
INVx3_ASAP7_75t_L g822 ( .A(n_607), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_607), .B(n_662), .Y(n_872) );
AND2x4_ASAP7_75t_L g898 ( .A(n_607), .B(n_761), .Y(n_898) );
INVx3_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g770 ( .A(n_608), .B(n_657), .Y(n_770) );
INVx1_ASAP7_75t_L g782 ( .A(n_608), .Y(n_782) );
AND2x2_ASAP7_75t_L g809 ( .A(n_608), .B(n_629), .Y(n_809) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g664 ( .A(n_609), .Y(n_664) );
OAI21x1_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_614), .B(n_618), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g644 ( .A(n_613), .B(n_645), .Y(n_644) );
INVx4_ASAP7_75t_L g681 ( .A(n_613), .Y(n_681) );
INVx1_ASAP7_75t_L g727 ( .A(n_614), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_618), .Y(n_728) );
AND2x2_ASAP7_75t_L g892 ( .A(n_620), .B(n_769), .Y(n_892) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_629), .Y(n_620) );
INVx2_ASAP7_75t_L g657 ( .A(n_621), .Y(n_657) );
INVx3_ASAP7_75t_L g663 ( .A(n_621), .Y(n_663) );
AND2x2_ASAP7_75t_L g779 ( .A(n_621), .B(n_642), .Y(n_779) );
INVx1_ASAP7_75t_L g801 ( .A(n_621), .Y(n_801) );
HB1xp67_ASAP7_75t_L g805 ( .A(n_621), .Y(n_805) );
AND2x4_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
OR2x2_ASAP7_75t_L g758 ( .A(n_629), .B(n_726), .Y(n_758) );
AND2x4_ASAP7_75t_L g761 ( .A(n_629), .B(n_663), .Y(n_761) );
AND2x2_ASAP7_75t_L g781 ( .A(n_629), .B(n_782), .Y(n_781) );
OA21x2_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_631), .B(n_638), .Y(n_629) );
OA21x2_ASAP7_75t_L g660 ( .A1(n_630), .A2(n_631), .B(n_638), .Y(n_660) );
OAI21xp33_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_658), .B(n_661), .Y(n_639) );
AND2x2_ASAP7_75t_L g905 ( .A(n_640), .B(n_757), .Y(n_905) );
AND2x2_ASAP7_75t_L g950 ( .A(n_640), .B(n_725), .Y(n_950) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g821 ( .A(n_641), .B(n_822), .Y(n_821) );
HB1xp67_ASAP7_75t_L g869 ( .A(n_641), .Y(n_869) );
OR2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_657), .Y(n_641) );
AND2x2_ASAP7_75t_L g662 ( .A(n_642), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g738 ( .A(n_642), .B(n_659), .Y(n_738) );
INVx2_ASAP7_75t_L g769 ( .A(n_642), .Y(n_769) );
INVx1_ASAP7_75t_L g789 ( .A(n_642), .Y(n_789) );
BUFx2_ASAP7_75t_L g819 ( .A(n_642), .Y(n_819) );
INVx2_ASAP7_75t_L g854 ( .A(n_642), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_642), .B(n_660), .Y(n_921) );
INVx3_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AOI21x1_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_646), .B(n_655), .Y(n_643) );
AOI21xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_650), .B(n_651), .Y(n_646) );
AND2x4_ASAP7_75t_L g828 ( .A(n_657), .B(n_729), .Y(n_828) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_659), .B(n_789), .Y(n_806) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g729 ( .A(n_660), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .Y(n_661) );
INVx2_ASAP7_75t_L g954 ( .A(n_662), .Y(n_954) );
INVx1_ASAP7_75t_L g724 ( .A(n_663), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_663), .B(n_854), .Y(n_853) );
INVx2_ASAP7_75t_L g802 ( .A(n_664), .Y(n_802) );
OR2x2_ASAP7_75t_L g852 ( .A(n_664), .B(n_853), .Y(n_852) );
AND2x2_ASAP7_75t_L g864 ( .A(n_664), .B(n_769), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_664), .B(n_805), .Y(n_890) );
AND2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_692), .Y(n_665) );
AND2x2_ASAP7_75t_L g893 ( .A(n_666), .B(n_894), .Y(n_893) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_684), .Y(n_666) );
AND2x2_ASAP7_75t_L g741 ( .A(n_667), .B(n_695), .Y(n_741) );
INVx1_ASAP7_75t_L g901 ( .A(n_667), .Y(n_901) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_668), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_668), .B(n_695), .Y(n_764) );
AND2x4_ASAP7_75t_L g773 ( .A(n_668), .B(n_743), .Y(n_773) );
INVx1_ASAP7_75t_L g818 ( .A(n_668), .Y(n_818) );
INVx1_ASAP7_75t_L g841 ( .A(n_668), .Y(n_841) );
OR2x2_ASAP7_75t_L g862 ( .A(n_668), .B(n_710), .Y(n_862) );
HB1xp67_ASAP7_75t_L g877 ( .A(n_668), .Y(n_877) );
AND2x2_ASAP7_75t_L g904 ( .A(n_668), .B(n_710), .Y(n_904) );
AO31x2_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_675), .A3(n_680), .B(n_682), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
NOR3xp33_ASAP7_75t_L g696 ( .A(n_681), .B(n_697), .C(n_701), .Y(n_696) );
AND2x4_ASAP7_75t_L g733 ( .A(n_684), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g847 ( .A(n_684), .Y(n_847) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g742 ( .A(n_685), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g775 ( .A(n_685), .Y(n_775) );
AND2x2_ASAP7_75t_L g902 ( .A(n_685), .B(n_694), .Y(n_902) );
HB1xp67_ASAP7_75t_L g938 ( .A(n_685), .Y(n_938) );
AND2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_691), .Y(n_685) );
AND2x2_ASAP7_75t_L g752 ( .A(n_686), .B(n_753), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_687), .B(n_690), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_710), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_693), .B(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g767 ( .A(n_694), .B(n_751), .Y(n_767) );
HB1xp67_ASAP7_75t_L g836 ( .A(n_694), .Y(n_836) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g734 ( .A(n_695), .Y(n_734) );
AND2x2_ASAP7_75t_L g774 ( .A(n_695), .B(n_775), .Y(n_774) );
HB1xp67_ASAP7_75t_L g832 ( .A(n_695), .Y(n_832) );
BUFx2_ASAP7_75t_R g881 ( .A(n_695), .Y(n_881) );
AO21x2_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_706), .B(n_707), .Y(n_695) );
NAND2xp5_ASAP7_75t_SL g712 ( .A(n_706), .B(n_713), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_710), .Y(n_732) );
AND2x2_ASAP7_75t_L g817 ( .A(n_710), .B(n_818), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_710), .B(n_734), .Y(n_895) );
AND2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
AND2x2_ASAP7_75t_L g751 ( .A(n_712), .B(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
AOI211xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_730), .B(n_735), .C(n_759), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
AND2x2_ASAP7_75t_L g756 ( .A(n_724), .B(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g790 ( .A(n_725), .Y(n_790) );
INVx2_ASAP7_75t_SL g952 ( .A(n_725), .Y(n_952) );
AND2x4_ASAP7_75t_L g725 ( .A(n_726), .B(n_729), .Y(n_725) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
INVx1_ASAP7_75t_L g909 ( .A(n_732), .Y(n_909) );
AND2x2_ASAP7_75t_L g810 ( .A(n_733), .B(n_773), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_733), .B(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g949 ( .A(n_733), .Y(n_949) );
OR2x2_ASAP7_75t_L g886 ( .A(n_734), .B(n_854), .Y(n_886) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_739), .B1(n_748), .B2(n_755), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
AND2x4_ASAP7_75t_L g941 ( .A(n_738), .B(n_942), .Y(n_941) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AOI222xp33_ASAP7_75t_L g771 ( .A1(n_740), .A2(n_761), .B1(n_772), .B2(n_776), .C1(n_783), .C2(n_786), .Y(n_771) );
AND2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
INVx1_ASAP7_75t_L g785 ( .A(n_741), .Y(n_785) );
AND2x4_ASAP7_75t_L g824 ( .A(n_742), .B(n_825), .Y(n_824) );
AND2x2_ASAP7_75t_L g944 ( .A(n_742), .B(n_818), .Y(n_944) );
INVx1_ASAP7_75t_L g851 ( .A(n_743), .Y(n_851) );
OAI21x1_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_745), .B(n_746), .Y(n_743) );
HB1xp67_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g940 ( .A(n_749), .Y(n_940) );
OR2x2_ASAP7_75t_L g749 ( .A(n_750), .B(n_754), .Y(n_749) );
OR2x2_ASAP7_75t_L g960 ( .A(n_750), .B(n_818), .Y(n_960) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g763 ( .A(n_751), .Y(n_763) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
AND2x2_ASAP7_75t_L g927 ( .A(n_757), .B(n_839), .Y(n_927) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g794 ( .A(n_758), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_762), .Y(n_759) );
OR2x2_ASAP7_75t_L g795 ( .A(n_760), .B(n_796), .Y(n_795) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g863 ( .A(n_761), .B(n_864), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_761), .B(n_885), .Y(n_884) );
AND2x2_ASAP7_75t_L g913 ( .A(n_761), .B(n_822), .Y(n_913) );
OR2x2_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
OR2x2_ASAP7_75t_L g784 ( .A(n_763), .B(n_785), .Y(n_784) );
OR2x2_ASAP7_75t_L g857 ( .A(n_763), .B(n_836), .Y(n_857) );
INVx1_ASAP7_75t_L g825 ( .A(n_764), .Y(n_825) );
NAND3xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_771), .C(n_791), .Y(n_765) );
NAND2xp33_ASAP7_75t_R g766 ( .A(n_767), .B(n_768), .Y(n_766) );
OAI21xp5_ASAP7_75t_L g926 ( .A1(n_768), .A2(n_927), .B(n_928), .Y(n_926) );
AND2x2_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
INVx1_ASAP7_75t_L g798 ( .A(n_769), .Y(n_798) );
INVx1_ASAP7_75t_L g839 ( .A(n_769), .Y(n_839) );
OAI21xp5_ASAP7_75t_L g943 ( .A1(n_772), .A2(n_944), .B(n_945), .Y(n_943) );
AND2x4_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .Y(n_772) );
AND2x2_ASAP7_75t_L g830 ( .A(n_773), .B(n_831), .Y(n_830) );
INVx2_ASAP7_75t_SL g848 ( .A(n_773), .Y(n_848) );
NAND2xp33_ASAP7_75t_L g816 ( .A(n_774), .B(n_817), .Y(n_816) );
INVx2_ASAP7_75t_SL g874 ( .A(n_774), .Y(n_874) );
AND2x2_ASAP7_75t_L g903 ( .A(n_774), .B(n_904), .Y(n_903) );
NAND2xp33_ASAP7_75t_L g776 ( .A(n_777), .B(n_780), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g883 ( .A(n_778), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_779), .B(n_809), .Y(n_808) );
AND2x2_ASAP7_75t_L g911 ( .A(n_779), .B(n_822), .Y(n_911) );
INVx3_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
AND2x2_ASAP7_75t_L g858 ( .A(n_781), .B(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
OAI21xp5_ASAP7_75t_SL g896 ( .A1(n_784), .A2(n_869), .B(n_897), .Y(n_896) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
NAND3xp33_ASAP7_75t_SL g888 ( .A(n_787), .B(n_889), .C(n_891), .Y(n_888) );
OR2x2_ASAP7_75t_L g787 ( .A(n_788), .B(n_790), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
OAI31xp33_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_799), .A3(n_807), .B(n_810), .Y(n_791) );
NAND2xp33_ASAP7_75t_SL g792 ( .A(n_793), .B(n_795), .Y(n_792) );
INVx2_ASAP7_75t_SL g793 ( .A(n_794), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_794), .B(n_869), .Y(n_868) );
OAI22xp33_ASAP7_75t_L g914 ( .A1(n_795), .A2(n_840), .B1(n_848), .B2(n_915), .Y(n_914) );
OR2x2_ASAP7_75t_L g946 ( .A(n_796), .B(n_890), .Y(n_946) );
INVx2_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_800), .B(n_803), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .Y(n_800) );
NOR2xp67_ASAP7_75t_L g920 ( .A(n_801), .B(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g942 ( .A(n_801), .Y(n_942) );
AND2x4_ASAP7_75t_L g827 ( .A(n_802), .B(n_828), .Y(n_827) );
OR2x2_ASAP7_75t_L g803 ( .A(n_804), .B(n_806), .Y(n_803) );
INVxp67_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
NOR2x1_ASAP7_75t_L g811 ( .A(n_812), .B(n_865), .Y(n_811) );
NAND4xp75_ASAP7_75t_L g812 ( .A(n_813), .B(n_833), .C(n_842), .D(n_855), .Y(n_812) );
NOR2x1_ASAP7_75t_SL g813 ( .A(n_814), .B(n_820), .Y(n_813) );
AND2x2_ASAP7_75t_L g814 ( .A(n_815), .B(n_819), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
AND2x2_ASAP7_75t_L g936 ( .A(n_817), .B(n_937), .Y(n_936) );
NAND2x1p5_ASAP7_75t_L g957 ( .A(n_819), .B(n_828), .Y(n_957) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_823), .B1(n_826), .B2(n_829), .Y(n_820) );
AND2x2_ASAP7_75t_L g923 ( .A(n_822), .B(n_828), .Y(n_923) );
INVx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx2_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
AND2x2_ASAP7_75t_L g837 ( .A(n_827), .B(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
OR2x2_ASAP7_75t_L g861 ( .A(n_831), .B(n_862), .Y(n_861) );
INVx2_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
NAND3xp33_ASAP7_75t_L g833 ( .A(n_834), .B(n_837), .C(n_840), .Y(n_833) );
HB1xp67_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
HB1xp67_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_838), .B(n_898), .Y(n_965) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_839), .B(n_913), .Y(n_912) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g930 ( .A(n_841), .Y(n_930) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
O2A1O1Ixp33_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_848), .B(n_849), .C(n_852), .Y(n_843) );
AOI221x1_ASAP7_75t_L g906 ( .A1(n_844), .A2(n_907), .B1(n_914), .B2(n_916), .C(n_917), .Y(n_906) );
BUFx2_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_845), .B(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
OAI22xp5_ASAP7_75t_L g878 ( .A1(n_848), .A2(n_879), .B1(n_883), .B2(n_884), .Y(n_878) );
INVx1_ASAP7_75t_L g958 ( .A(n_849), .Y(n_958) );
NOR2xp33_ASAP7_75t_L g925 ( .A(n_850), .B(n_874), .Y(n_925) );
AOI33xp33_ASAP7_75t_L g948 ( .A1(n_850), .A2(n_944), .A3(n_949), .B1(n_950), .B2(n_951), .B3(n_953), .Y(n_948) );
INVx2_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
BUFx2_ASAP7_75t_L g859 ( .A(n_854), .Y(n_859) );
AOI22xp5_ASAP7_75t_L g855 ( .A1(n_856), .A2(n_858), .B1(n_860), .B2(n_863), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx2_ASAP7_75t_L g882 ( .A(n_862), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_866), .B(n_887), .Y(n_865) );
O2A1O1Ixp33_ASAP7_75t_L g866 ( .A1(n_867), .A2(n_870), .B(n_873), .C(n_878), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVxp67_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
BUFx2_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
NOR2xp33_ASAP7_75t_L g873 ( .A(n_874), .B(n_875), .Y(n_873) );
OR2x2_ASAP7_75t_L g963 ( .A(n_874), .B(n_900), .Y(n_963) );
INVxp67_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_880), .B(n_882), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
AOI21xp5_ASAP7_75t_L g887 ( .A1(n_888), .A2(n_893), .B(n_896), .Y(n_887) );
HB1xp67_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
INVx1_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
AOI22xp5_ASAP7_75t_L g897 ( .A1(n_898), .A2(n_899), .B1(n_903), .B2(n_905), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_898), .B(n_936), .Y(n_935) );
AND2x2_ASAP7_75t_L g899 ( .A(n_900), .B(n_902), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
BUFx2_ASAP7_75t_L g916 ( .A(n_902), .Y(n_916) );
OAI21xp33_ASAP7_75t_L g907 ( .A1(n_908), .A2(n_910), .B(n_912), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
INVxp33_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
A2O1A1Ixp33_ASAP7_75t_L g917 ( .A1(n_918), .A2(n_922), .B(n_924), .C(n_926), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
BUFx2_ASAP7_75t_SL g919 ( .A(n_920), .Y(n_919) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_923), .A2(n_956), .B1(n_958), .B2(n_959), .Y(n_955) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
NOR2xp67_ASAP7_75t_L g931 ( .A(n_932), .B(n_947), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_933), .B(n_943), .Y(n_932) );
INVxp67_ASAP7_75t_SL g933 ( .A(n_934), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_935), .B(n_939), .Y(n_934) );
INVx2_ASAP7_75t_SL g937 ( .A(n_938), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_940), .B(n_941), .Y(n_939) );
INVx1_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
NAND3xp33_ASAP7_75t_L g947 ( .A(n_948), .B(n_955), .C(n_961), .Y(n_947) );
INVx2_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
INVx2_ASAP7_75t_SL g953 ( .A(n_954), .Y(n_953) );
INVx1_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
INVx2_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
NAND2xp5_ASAP7_75t_L g961 ( .A(n_962), .B(n_964), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
INVx1_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
INVx1_ASAP7_75t_SL g966 ( .A(n_967), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
INVx2_ASAP7_75t_L g980 ( .A(n_968), .Y(n_980) );
INVx1_ASAP7_75t_SL g972 ( .A(n_973), .Y(n_972) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_976), .B(n_981), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
BUFx3_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
BUFx12f_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
CKINVDCx11_ASAP7_75t_R g979 ( .A(n_980), .Y(n_979) );
INVx1_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
HB1xp67_ASAP7_75t_SL g985 ( .A(n_986), .Y(n_985) );
INVx1_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
INVx1_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
BUFx2_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
INVx1_ASAP7_75t_L g997 ( .A(n_990), .Y(n_997) );
AND2x4_ASAP7_75t_L g990 ( .A(n_991), .B(n_993), .Y(n_990) );
CKINVDCx20_ASAP7_75t_R g991 ( .A(n_992), .Y(n_991) );
endmodule