module real_jpeg_25139_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_1),
.A2(n_49),
.B1(n_53),
.B2(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_1),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_1),
.A2(n_42),
.B1(n_43),
.B2(n_167),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_1),
.A2(n_62),
.B1(n_63),
.B2(n_167),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_167),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_2),
.A2(n_42),
.B1(n_43),
.B2(n_88),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_2),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_2),
.A2(n_62),
.B1(n_63),
.B2(n_88),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_2),
.A2(n_53),
.B1(n_88),
.B2(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_88),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_3),
.A2(n_111),
.B(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_3),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_3),
.B(n_41),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_L g233 ( 
.A1(n_3),
.A2(n_62),
.B1(n_63),
.B2(n_164),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_3),
.B(n_30),
.C(n_64),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_3),
.B(n_86),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_3),
.A2(n_27),
.B1(n_252),
.B2(n_259),
.Y(n_261)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_4),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_6),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_6),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_6),
.A2(n_42),
.B1(n_43),
.B2(n_109),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_6),
.A2(n_62),
.B1(n_63),
.B2(n_109),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_109),
.Y(n_244)
);

INVx8_ASAP7_75t_SL g47 ( 
.A(n_7),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_8),
.A2(n_42),
.B1(n_43),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_8),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_8),
.A2(n_53),
.B1(n_157),
.B2(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_8),
.A2(n_62),
.B1(n_63),
.B2(n_157),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_157),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_9),
.A2(n_62),
.B1(n_63),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_9),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_9),
.A2(n_42),
.B1(n_43),
.B2(n_69),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_69),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_10),
.A2(n_49),
.B1(n_53),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_10),
.A2(n_56),
.B1(n_62),
.B2(n_63),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_56),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_56),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_11),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_12),
.A2(n_37),
.B1(n_49),
.B2(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_12),
.A2(n_37),
.B1(n_62),
.B2(n_63),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_12),
.A2(n_37),
.B1(n_42),
.B2(n_43),
.Y(n_180)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_15),
.Y(n_99)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_15),
.Y(n_253)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_138),
.B1(n_139),
.B2(n_315),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_18),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_137),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_118),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_21),
.B(n_118),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_72),
.C(n_92),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_22),
.A2(n_23),
.B1(n_72),
.B2(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_58),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_38),
.B2(n_57),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_25),
.B(n_59),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_25),
.A2(n_57),
.B(n_58),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_25),
.A2(n_26),
.B1(n_59),
.B2(n_300),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_33),
.B(n_35),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_27),
.A2(n_148),
.B(n_150),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_27),
.A2(n_35),
.B(n_150),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_27),
.A2(n_97),
.B(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_27),
.A2(n_33),
.B1(n_249),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_28),
.B(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_28),
.A2(n_31),
.B1(n_149),
.B2(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_28),
.A2(n_248),
.B1(n_250),
.B2(n_251),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_29),
.A2(n_30),
.B1(n_64),
.B2(n_66),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_29),
.B(n_263),
.Y(n_262)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_31),
.Y(n_196)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_33),
.B(n_164),
.Y(n_263)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_36),
.B(n_98),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_51),
.B(n_54),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_39),
.A2(n_108),
.B(n_113),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_39),
.B(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_39),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_39),
.A2(n_41),
.B1(n_166),
.B2(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_39),
.A2(n_41),
.B1(n_108),
.B2(n_174),
.Y(n_287)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_48),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_40),
.B(n_52),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_40),
.A2(n_122),
.B(n_124),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_40),
.A2(n_160),
.B1(n_161),
.B2(n_165),
.Y(n_159)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_42),
.A2(n_43),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_42),
.A2(n_46),
.B(n_163),
.C(n_183),
.Y(n_182)
);

HAxp5_ASAP7_75t_SL g210 ( 
.A(n_42),
.B(n_164),
.CON(n_210),
.SN(n_210)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

NAND3xp33_ASAP7_75t_L g183 ( 
.A(n_43),
.B(n_45),
.C(n_176),
.Y(n_183)
);

OAI32xp33_ASAP7_75t_L g209 ( 
.A1(n_43),
.A2(n_63),
.A3(n_85),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_46),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_49),
.Y(n_176)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_59),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_68),
.B(n_70),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_60),
.B(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_60),
.A2(n_68),
.B1(n_104),
.B2(n_106),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_60),
.A2(n_70),
.B(n_77),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_60),
.A2(n_106),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_60),
.A2(n_75),
.B(n_216),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_60),
.A2(n_106),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_60),
.A2(n_106),
.B1(n_215),
.B2(n_234),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_67),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_61)
);

AO22x1_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_63),
.B1(n_84),
.B2(n_85),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_62),
.B(n_84),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_63),
.B(n_236),
.Y(n_235)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_67),
.A2(n_76),
.B(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_67),
.A2(n_78),
.B(n_105),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_67),
.B(n_164),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_72),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_80),
.B(n_91),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_80),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_81),
.A2(n_90),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g178 ( 
.A1(n_81),
.A2(n_158),
.B(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_81),
.A2(n_90),
.B1(n_156),
.B2(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_81),
.A2(n_132),
.B(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_82),
.B(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_82),
.A2(n_130),
.B(n_131),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_82),
.A2(n_86),
.B1(n_201),
.B2(n_210),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_86),
.B(n_117),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_86),
.B(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_87),
.A2(n_90),
.B(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

FAx1_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_119),
.CI(n_136),
.CON(n_118),
.SN(n_118)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_92),
.A2(n_93),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_107),
.C(n_114),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_94),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_102),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_95),
.A2(n_96),
.B1(n_102),
.B2(n_103),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_99),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_100),
.A2(n_187),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_101),
.B(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_107),
.A2(n_114),
.B1(n_115),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_107),
.Y(n_303)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_112),
.B(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx24_ASAP7_75t_SL g316 ( 
.A(n_118),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_126),
.B2(n_127),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_133),
.B2(n_134),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_308),
.B(n_314),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_295),
.B(n_307),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_202),
.B(n_278),
.C(n_294),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_188),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_143),
.B(n_188),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_170),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_152),
.B1(n_168),
.B2(n_169),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_145),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_145),
.B(n_169),
.C(n_170),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_146),
.B(n_147),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.C(n_159),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_153),
.A2(n_154),
.B1(n_155),
.B2(n_191),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_155),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_159),
.B(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_181),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_177),
.B2(n_178),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_173),
.B(n_177),
.C(n_181),
.Y(n_292)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_180),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_184),
.B1(n_185),
.B2(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.C(n_194),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_189),
.B(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_192),
.B(n_194),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.C(n_199),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_197),
.B1(n_198),
.B2(n_221),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_195),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_273),
.B(n_277),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_228),
.B(n_272),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_217),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_207),
.B(n_217),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.C(n_214),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_208),
.B(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_212),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_213),
.B(n_214),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_222),
.B2(n_223),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_218),
.B(n_225),
.C(n_227),
.Y(n_274)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_224),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_267),
.B(n_271),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_245),
.B(n_266),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_237),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_231),
.B(n_237),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_235),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_235),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_243),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_242),
.C(n_243),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_241),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_244),
.Y(n_250)
);

AOI21xp33_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_255),
.B(n_265),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_254),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_254),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_260),
.B(n_264),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_257),
.B(n_258),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_268),
.B(n_269),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_274),
.B(n_275),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_280),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_292),
.B2(n_293),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_284),
.C(n_293),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_291),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_288),
.C(n_291),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_292),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_296),
.B(n_297),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_306),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_301),
.B1(n_304),
.B2(n_305),
.Y(n_298)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_299),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_305),
.C(n_306),
.Y(n_309)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_301),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_309),
.B(n_310),
.Y(n_314)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);


endmodule