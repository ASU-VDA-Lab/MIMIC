module fake_jpeg_67_n_52 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_52);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_52;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_4),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

INVx4_ASAP7_75t_SL g9 ( 
.A(n_1),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

AND2x2_ASAP7_75t_L g13 ( 
.A(n_2),
.B(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_3),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_25),
.Y(n_31)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_21),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_15),
.Y(n_19)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_0),
.C(n_1),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_24),
.C(n_11),
.Y(n_33)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_3),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_8),
.Y(n_26)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_16),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_24)
);

CKINVDCx12_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_30),
.C(n_24),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_16),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_33),
.B(n_24),
.C(n_22),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_24),
.A2(n_20),
.B1(n_19),
.B2(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_12),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_35),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_29),
.A2(n_19),
.B1(n_27),
.B2(n_26),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_36),
.B(n_38),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_30),
.Y(n_41)
);

INVxp33_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_33),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_29),
.C(n_11),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_45),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_39),
.B1(n_40),
.B2(n_29),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_44),
.B(n_45),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_18),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_49),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_46),
.A2(n_10),
.B1(n_21),
.B2(n_14),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_46),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_49),
.C(n_32),
.Y(n_52)
);


endmodule