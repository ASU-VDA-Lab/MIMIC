module fake_jpeg_8290_n_317 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_36),
.B(n_37),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_38),
.B(n_23),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_19),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_28),
.Y(n_45)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_54),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_55),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_25),
.B1(n_27),
.B2(n_22),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_61),
.B1(n_36),
.B2(n_37),
.Y(n_82)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_23),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_27),
.B1(n_19),
.B2(n_17),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_56),
.A2(n_64),
.B1(n_41),
.B2(n_37),
.Y(n_76)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_62),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_27),
.B1(n_19),
.B2(n_31),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_43),
.B(n_34),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_66),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_17),
.B1(n_34),
.B2(n_26),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_36),
.A2(n_22),
.B(n_33),
.C(n_30),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_67),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_33),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_44),
.B1(n_41),
.B2(n_38),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_70),
.A2(n_21),
.B1(n_53),
.B2(n_32),
.Y(n_108)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_80),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_76),
.A2(n_79),
.B(n_91),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_77),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_41),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_66),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_82),
.B(n_89),
.Y(n_106)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_85),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_38),
.C(n_40),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_62),
.C(n_58),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_68),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_95),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_39),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_90),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_47),
.A2(n_26),
.B1(n_30),
.B2(n_29),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_39),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_92),
.B(n_0),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_31),
.Y(n_94)
);

FAx1_ASAP7_75t_SL g107 ( 
.A(n_94),
.B(n_84),
.CI(n_71),
.CON(n_107),
.SN(n_107)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_51),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_100),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_48),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_98),
.B(n_121),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_57),
.B1(n_39),
.B2(n_67),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_99),
.A2(n_102),
.B1(n_114),
.B2(n_116),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_77),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_101),
.B(n_108),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_89),
.A2(n_57),
.B1(n_39),
.B2(n_29),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_110),
.C(n_78),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_92),
.A2(n_55),
.B(n_53),
.C(n_21),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_104),
.A2(n_107),
.B(n_18),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_77),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_109),
.B(n_111),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_53),
.C(n_59),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_46),
.B1(n_32),
.B2(n_24),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_82),
.A2(n_32),
.B1(n_18),
.B2(n_9),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_18),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_118),
.B(n_18),
.Y(n_145)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_120),
.B(n_122),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_79),
.B(n_1),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_125),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_119),
.A2(n_79),
.B(n_85),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_124),
.A2(n_132),
.B(n_145),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_117),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_127),
.B(n_129),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_94),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_141),
.C(n_120),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_117),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_96),
.A2(n_75),
.B1(n_95),
.B2(n_81),
.Y(n_130)
);

OAI22x1_ASAP7_75t_L g176 ( 
.A1(n_130),
.A2(n_97),
.B1(n_115),
.B2(n_112),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_119),
.A2(n_88),
.B(n_94),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_97),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_133),
.B(n_139),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_88),
.B1(n_73),
.B2(n_74),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_137),
.A2(n_142),
.B1(n_126),
.B2(n_139),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_106),
.A2(n_81),
.B1(n_69),
.B2(n_73),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_138),
.A2(n_144),
.B1(n_97),
.B2(n_3),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_113),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_99),
.Y(n_142)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_143),
.A2(n_122),
.B(n_121),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_116),
.A2(n_69),
.B1(n_18),
.B2(n_90),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_98),
.B(n_1),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_146),
.A2(n_147),
.B(n_149),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_105),
.A2(n_90),
.B(n_78),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_105),
.B(n_16),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_148),
.B(n_9),
.Y(n_179)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_103),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_152),
.A2(n_159),
.B(n_175),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_110),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_165),
.C(n_170),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_123),
.A2(n_103),
.B1(n_107),
.B2(n_98),
.Y(n_155)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_155),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_156),
.B(n_160),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_132),
.A2(n_118),
.B(n_107),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_124),
.A2(n_107),
.B(n_114),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_164),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_167),
.Y(n_189)
);

BUFx24_ASAP7_75t_SL g164 ( 
.A(n_125),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_108),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_101),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_111),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_172),
.C(n_136),
.Y(n_204)
);

OAI32xp33_ASAP7_75t_L g173 ( 
.A1(n_149),
.A2(n_115),
.A3(n_109),
.B1(n_100),
.B2(n_12),
.Y(n_173)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_127),
.B(n_1),
.Y(n_175)
);

OA22x2_ASAP7_75t_L g198 ( 
.A1(n_176),
.A2(n_181),
.B1(n_182),
.B2(n_144),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_180),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_178),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_179),
.B(n_148),
.Y(n_197)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_137),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_136),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_153),
.B(n_150),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_185),
.B(n_6),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_145),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_187),
.B(n_195),
.C(n_204),
.Y(n_232)
);

NAND3xp33_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_129),
.C(n_134),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_188),
.B(n_197),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_178),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_191),
.B(n_199),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_146),
.Y(n_193)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_202),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_135),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_198),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_158),
.B(n_135),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_138),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_201),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_134),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_156),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_205),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_167),
.A2(n_126),
.B1(n_12),
.B2(n_5),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_206),
.A2(n_209),
.B(n_159),
.Y(n_222)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_163),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_208),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_157),
.B(n_151),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_173),
.A2(n_182),
.B1(n_174),
.B2(n_175),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_155),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_228),
.Y(n_236)
);

INVxp33_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_154),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_213),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_169),
.B(n_152),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_218),
.A2(n_221),
.B(n_198),
.Y(n_248)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_220),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_194),
.A2(n_203),
.B1(n_200),
.B2(n_209),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_165),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_206),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_203),
.A2(n_152),
.B1(n_170),
.B2(n_181),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_223),
.A2(n_231),
.B1(n_7),
.B2(n_10),
.Y(n_250)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_226),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_196),
.A2(n_175),
.B1(n_4),
.B2(n_2),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_225),
.A2(n_197),
.B1(n_198),
.B2(n_196),
.Y(n_243)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_183),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_10),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_193),
.B(n_4),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_230),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_185),
.B(n_6),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_190),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_234),
.B(n_7),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_204),
.C(n_187),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_237),
.C(n_244),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_195),
.C(n_190),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_245),
.Y(n_261)
);

NOR2xp67_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_186),
.Y(n_241)
);

NAND3xp33_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_252),
.C(n_223),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_242),
.A2(n_248),
.B(n_222),
.Y(n_260)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_243),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_228),
.C(n_218),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_198),
.C(n_8),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_250),
.A2(n_7),
.B1(n_13),
.B2(n_15),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_234),
.Y(n_262)
);

NOR2x1_ASAP7_75t_L g252 ( 
.A(n_212),
.B(n_16),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_213),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_253),
.B(n_254),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_216),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_240),
.A2(n_231),
.B1(n_215),
.B2(n_219),
.Y(n_256)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_256),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_257),
.B(n_258),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_246),
.B(n_217),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_240),
.B(n_217),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_268),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_262),
.Y(n_273)
);

FAx1_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_221),
.CI(n_227),
.CON(n_263),
.SN(n_263)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_245),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_239),
.A2(n_221),
.B1(n_224),
.B2(n_229),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_264),
.A2(n_265),
.B1(n_247),
.B2(n_251),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_239),
.A2(n_211),
.B1(n_225),
.B2(n_226),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_243),
.A2(n_230),
.B1(n_13),
.B2(n_14),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_266),
.Y(n_279)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_252),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_270),
.A2(n_247),
.B1(n_250),
.B2(n_238),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_271),
.A2(n_283),
.B1(n_263),
.B2(n_269),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_255),
.A2(n_264),
.B(n_249),
.Y(n_274)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_244),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_275),
.B(n_261),
.Y(n_286)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_265),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_263),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_249),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_280),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_261),
.Y(n_285)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_284),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_289),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_288),
.Y(n_295)
);

NOR2xp67_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_271),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_287),
.A2(n_278),
.B(n_277),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_267),
.C(n_235),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_237),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_290),
.A2(n_282),
.B(n_236),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_279),
.B(n_262),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_294),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_279),
.B(n_236),
.Y(n_294)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_297),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_276),
.Y(n_299)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_299),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_300),
.A2(n_291),
.B(n_285),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_282),
.Y(n_301)
);

OAI21x1_ASAP7_75t_L g305 ( 
.A1(n_301),
.A2(n_303),
.B(n_300),
.Y(n_305)
);

INVx11_ASAP7_75t_L g303 ( 
.A(n_284),
.Y(n_303)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_304),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_305),
.A2(n_307),
.B1(n_308),
.B2(n_303),
.Y(n_311)
);

AOI21x1_ASAP7_75t_L g307 ( 
.A1(n_301),
.A2(n_289),
.B(n_15),
.Y(n_307)
);

OA21x2_ASAP7_75t_SL g308 ( 
.A1(n_295),
.A2(n_296),
.B(n_302),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_306),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_310),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_312),
.B(n_311),
.Y(n_314)
);

AO21x1_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_309),
.B(n_298),
.Y(n_315)
);

MAJx2_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_296),
.C(n_15),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_316),
.B(n_16),
.Y(n_317)
);


endmodule