module fake_jpeg_11444_n_169 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_169);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_12),
.B(n_47),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_25),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_13),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_5),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_43),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_6),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_45),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_19),
.B(n_13),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_22),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_64),
.Y(n_80)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_70),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_49),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_77),
.Y(n_85)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

HAxp5_ASAP7_75t_SL g75 ( 
.A(n_58),
.B(n_0),
.CON(n_75),
.SN(n_75)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_76),
.Y(n_83)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_23),
.B(n_46),
.C(n_44),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_65),
.Y(n_77)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_82),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_69),
.B(n_51),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_54),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_91),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_52),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_86),
.B(n_90),
.Y(n_107)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_77),
.A2(n_65),
.B1(n_58),
.B2(n_53),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_89),
.A2(n_71),
.B1(n_68),
.B2(n_59),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_61),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_56),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_98),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_67),
.C(n_66),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_95),
.C(n_4),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_55),
.C(n_62),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_89),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_104),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_59),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_62),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_108),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_68),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_11),
.C(n_12),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_88),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_63),
.B1(n_60),
.B2(n_50),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_110),
.A2(n_87),
.B1(n_7),
.B2(n_8),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_99),
.B(n_107),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_112),
.B(n_116),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_SL g114 ( 
.A(n_106),
.B(n_48),
.C(n_2),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_132),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_87),
.B(n_21),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_31),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_101),
.B(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_94),
.B(n_1),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_120),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_93),
.B(n_3),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_122),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_3),
.B(n_4),
.C(n_7),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_124),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_127),
.Y(n_141)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_98),
.B(n_8),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_99),
.B(n_10),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_131),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_10),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_133),
.B(n_134),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_32),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_125),
.C(n_114),
.Y(n_153)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_139),
.B(n_28),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_123),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_144),
.B(n_146),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_117),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_145),
.A2(n_147),
.B1(n_124),
.B2(n_120),
.Y(n_151)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_117),
.A2(n_18),
.B1(n_26),
.B2(n_27),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_152),
.Y(n_158)
);

A2O1A1O1Ixp25_ASAP7_75t_L g152 ( 
.A1(n_135),
.A2(n_138),
.B(n_132),
.C(n_141),
.D(n_142),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_155),
.C(n_137),
.Y(n_160)
);

AOI221xp5_ASAP7_75t_L g155 ( 
.A1(n_145),
.A2(n_122),
.B1(n_115),
.B2(n_34),
.C(n_38),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_157),
.A2(n_147),
.B1(n_143),
.B2(n_154),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_159),
.A2(n_160),
.B(n_161),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_136),
.Y(n_161)
);

AOI321xp33_ASAP7_75t_L g162 ( 
.A1(n_158),
.A2(n_152),
.A3(n_149),
.B1(n_136),
.B2(n_154),
.C(n_150),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_162),
.A2(n_161),
.B(n_148),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_163),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_165),
.B(n_134),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_140),
.Y(n_167)
);

NOR3xp33_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_33),
.C(n_39),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_40),
.Y(n_169)
);


endmodule