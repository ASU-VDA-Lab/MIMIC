module fake_netlist_1_9514_n_666 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_666);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_666;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_44), .Y(n_79) );
CKINVDCx14_ASAP7_75t_R g80 ( .A(n_52), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_8), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_13), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_20), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_66), .Y(n_84) );
HB1xp67_ASAP7_75t_L g85 ( .A(n_45), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_35), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_30), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_8), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_75), .Y(n_89) );
HB1xp67_ASAP7_75t_L g90 ( .A(n_22), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_62), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_13), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_50), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_17), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_58), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_16), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_18), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_57), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_7), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_63), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_5), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_67), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_48), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_59), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_68), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_37), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_73), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_14), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_46), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_49), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_3), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_1), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_7), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_71), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_5), .Y(n_115) );
BUFx2_ASAP7_75t_L g116 ( .A(n_65), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_74), .Y(n_117) );
INVxp33_ASAP7_75t_L g118 ( .A(n_41), .Y(n_118) );
INVxp33_ASAP7_75t_SL g119 ( .A(n_27), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_77), .Y(n_120) );
CKINVDCx16_ASAP7_75t_R g121 ( .A(n_19), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_3), .Y(n_122) );
AND2x2_ASAP7_75t_L g123 ( .A(n_116), .B(n_0), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_79), .Y(n_124) );
OAI21x1_ASAP7_75t_L g125 ( .A1(n_93), .A2(n_33), .B(n_76), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_116), .B(n_0), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_85), .B(n_1), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_93), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_79), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_92), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_83), .Y(n_131) );
INVx1_ASAP7_75t_SL g132 ( .A(n_81), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_121), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_83), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_84), .Y(n_135) );
AND2x6_ASAP7_75t_L g136 ( .A(n_84), .B(n_34), .Y(n_136) );
INVx3_ASAP7_75t_L g137 ( .A(n_82), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_109), .Y(n_138) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_88), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_113), .Y(n_140) );
AND2x6_ASAP7_75t_L g141 ( .A(n_86), .B(n_32), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_86), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_118), .B(n_2), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_80), .Y(n_144) );
BUFx3_ASAP7_75t_L g145 ( .A(n_109), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_89), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_89), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_90), .B(n_2), .Y(n_148) );
INVx4_ASAP7_75t_L g149 ( .A(n_87), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_91), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g151 ( .A(n_94), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_91), .Y(n_152) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_94), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_95), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_95), .B(n_4), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_98), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_98), .Y(n_157) );
AOI22xp5_ASAP7_75t_L g158 ( .A1(n_99), .A2(n_4), .B1(n_6), .B2(n_9), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_119), .Y(n_159) );
BUFx3_ASAP7_75t_L g160 ( .A(n_136), .Y(n_160) );
AOI22xp33_ASAP7_75t_L g161 ( .A1(n_153), .A2(n_99), .B1(n_101), .B2(n_115), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_149), .B(n_105), .Y(n_162) );
CKINVDCx16_ASAP7_75t_R g163 ( .A(n_139), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_149), .B(n_114), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_123), .B(n_82), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_146), .Y(n_166) );
BUFx2_ASAP7_75t_L g167 ( .A(n_140), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_149), .B(n_97), .Y(n_168) );
INVxp67_ASAP7_75t_SL g169 ( .A(n_123), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_146), .Y(n_170) );
AND2x6_ASAP7_75t_L g171 ( .A(n_143), .B(n_107), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_125), .Y(n_172) );
CKINVDCx16_ASAP7_75t_R g173 ( .A(n_132), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_149), .B(n_103), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_133), .Y(n_175) );
NAND2xp33_ASAP7_75t_L g176 ( .A(n_136), .B(n_104), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_124), .B(n_96), .Y(n_177) );
AND2x4_ASAP7_75t_L g178 ( .A(n_124), .B(n_108), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_146), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_146), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_146), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_144), .B(n_129), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_143), .B(n_96), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_129), .B(n_100), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_131), .B(n_110), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_146), .Y(n_186) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_126), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_131), .B(n_101), .Y(n_188) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_151), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_154), .Y(n_190) );
INVx4_ASAP7_75t_L g191 ( .A(n_136), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_134), .B(n_102), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_154), .Y(n_193) );
INVx2_ASAP7_75t_SL g194 ( .A(n_134), .Y(n_194) );
INVx1_ASAP7_75t_SL g195 ( .A(n_130), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_135), .B(n_102), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_154), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_135), .B(n_111), .Y(n_198) );
NAND2x1p5_ASAP7_75t_L g199 ( .A(n_142), .B(n_106), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_125), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_154), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_159), .B(n_147), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_127), .Y(n_203) );
AND2x6_ASAP7_75t_L g204 ( .A(n_142), .B(n_106), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_194), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_194), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_173), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_180), .Y(n_208) );
INVxp67_ASAP7_75t_SL g209 ( .A(n_199), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_180), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_169), .B(n_157), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_176), .A2(n_157), .B(n_156), .Y(n_212) );
INVx4_ASAP7_75t_L g213 ( .A(n_191), .Y(n_213) );
INVx5_ASAP7_75t_L g214 ( .A(n_204), .Y(n_214) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_173), .Y(n_215) );
BUFx2_ASAP7_75t_L g216 ( .A(n_171), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_187), .B(n_156), .Y(n_217) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_160), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_199), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_202), .B(n_148), .Y(n_220) );
OR2x6_ASAP7_75t_L g221 ( .A(n_167), .B(n_155), .Y(n_221) );
NOR2x1p5_ASAP7_75t_L g222 ( .A(n_175), .B(n_115), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_191), .A2(n_150), .B(n_147), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_199), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_188), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_160), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_165), .B(n_183), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_191), .B(n_150), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_181), .Y(n_229) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_163), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_172), .Y(n_231) );
OR2x6_ASAP7_75t_L g232 ( .A(n_167), .B(n_111), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_163), .Y(n_233) );
NOR2x1_ASAP7_75t_L g234 ( .A(n_182), .B(n_145), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_203), .B(n_120), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_181), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_165), .B(n_152), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_183), .B(n_145), .Y(n_238) );
INVxp67_ASAP7_75t_SL g239 ( .A(n_188), .Y(n_239) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_172), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_203), .B(n_152), .Y(n_241) );
NOR2x1_ASAP7_75t_L g242 ( .A(n_164), .B(n_145), .Y(n_242) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_189), .Y(n_243) );
NOR3xp33_ASAP7_75t_SL g244 ( .A(n_175), .B(n_122), .C(n_112), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_188), .Y(n_245) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_195), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_186), .Y(n_247) );
BUFx4f_ASAP7_75t_SL g248 ( .A(n_171), .Y(n_248) );
INVxp67_ASAP7_75t_SL g249 ( .A(n_188), .Y(n_249) );
BUFx2_ASAP7_75t_L g250 ( .A(n_171), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_177), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_171), .A2(n_136), .B1(n_141), .B2(n_152), .Y(n_252) );
BUFx2_ASAP7_75t_L g253 ( .A(n_171), .Y(n_253) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_172), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_186), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_172), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_178), .B(n_136), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_168), .B(n_137), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_L g259 ( .A1(n_227), .A2(n_192), .B(n_198), .C(n_185), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_225), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_209), .A2(n_178), .B1(n_161), .B2(n_158), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_245), .Y(n_262) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_214), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_225), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_232), .B(n_198), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_257), .A2(n_200), .B(n_172), .Y(n_266) );
OAI22xp5_ASAP7_75t_L g267 ( .A1(n_239), .A2(n_178), .B1(n_158), .B2(n_162), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_245), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_256), .A2(n_200), .B(n_174), .Y(n_269) );
AO32x2_ASAP7_75t_L g270 ( .A1(n_231), .A2(n_200), .A3(n_171), .B1(n_136), .B2(n_141), .Y(n_270) );
BUFx2_ASAP7_75t_L g271 ( .A(n_215), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g272 ( .A1(n_249), .A2(n_177), .B1(n_171), .B2(n_196), .Y(n_272) );
O2A1O1Ixp33_ASAP7_75t_L g273 ( .A1(n_237), .A2(n_177), .B(n_108), .C(n_112), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_256), .A2(n_200), .B(n_184), .Y(n_274) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_214), .Y(n_275) );
AOI222xp33_ASAP7_75t_L g276 ( .A1(n_230), .A2(n_177), .B1(n_137), .B2(n_128), .C1(n_138), .C2(n_204), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_225), .Y(n_277) );
AOI21xp33_ASAP7_75t_L g278 ( .A1(n_220), .A2(n_200), .B(n_110), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_238), .Y(n_279) );
BUFx8_ASAP7_75t_SL g280 ( .A(n_233), .Y(n_280) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_232), .Y(n_281) );
BUFx3_ASAP7_75t_L g282 ( .A(n_233), .Y(n_282) );
AOI22xp33_ASAP7_75t_L g283 ( .A1(n_216), .A2(n_204), .B1(n_136), .B2(n_141), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_223), .A2(n_166), .B(n_201), .Y(n_284) );
O2A1O1Ixp33_ASAP7_75t_L g285 ( .A1(n_211), .A2(n_137), .B(n_128), .C(n_138), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_214), .B(n_154), .Y(n_286) );
OR2x6_ASAP7_75t_L g287 ( .A(n_232), .B(n_137), .Y(n_287) );
O2A1O1Ixp33_ASAP7_75t_L g288 ( .A1(n_217), .A2(n_107), .B(n_117), .C(n_197), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_238), .Y(n_289) );
INVx2_ASAP7_75t_SL g290 ( .A(n_232), .Y(n_290) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_214), .Y(n_291) );
BUFx8_ASAP7_75t_L g292 ( .A(n_216), .Y(n_292) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_246), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g294 ( .A1(n_250), .A2(n_204), .B1(n_141), .B2(n_154), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_241), .B(n_204), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_251), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_219), .B(n_204), .Y(n_297) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_214), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_219), .B(n_204), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_212), .A2(n_201), .B(n_197), .Y(n_300) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_224), .B(n_117), .Y(n_301) );
AO21x2_ASAP7_75t_L g302 ( .A1(n_205), .A2(n_193), .B(n_190), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_205), .A2(n_193), .B(n_190), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_224), .Y(n_304) );
INVx1_ASAP7_75t_SL g305 ( .A(n_207), .Y(n_305) );
CKINVDCx16_ASAP7_75t_R g306 ( .A(n_243), .Y(n_306) );
OAI21x1_ASAP7_75t_L g307 ( .A1(n_266), .A2(n_252), .B(n_242), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_263), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_262), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_302), .Y(n_310) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_263), .Y(n_311) );
NAND3xp33_ASAP7_75t_L g312 ( .A(n_273), .B(n_244), .C(n_258), .Y(n_312) );
OAI21xp5_ASAP7_75t_L g313 ( .A1(n_266), .A2(n_206), .B(n_228), .Y(n_313) );
OAI21x1_ASAP7_75t_L g314 ( .A1(n_269), .A2(n_206), .B(n_234), .Y(n_314) );
AO21x2_ASAP7_75t_L g315 ( .A1(n_278), .A2(n_166), .B(n_179), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_280), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_268), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_261), .A2(n_248), .B1(n_253), .B2(n_250), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g319 ( .A1(n_287), .A2(n_253), .B1(n_254), .B2(n_240), .Y(n_319) );
OAI21x1_ASAP7_75t_L g320 ( .A1(n_269), .A2(n_179), .B(n_170), .Y(n_320) );
AO21x2_ASAP7_75t_L g321 ( .A1(n_274), .A2(n_235), .B(n_229), .Y(n_321) );
OAI21x1_ASAP7_75t_L g322 ( .A1(n_274), .A2(n_170), .B(n_254), .Y(n_322) );
BUFx3_ASAP7_75t_L g323 ( .A(n_263), .Y(n_323) );
AND2x4_ASAP7_75t_L g324 ( .A(n_287), .B(n_213), .Y(n_324) );
CKINVDCx6p67_ASAP7_75t_R g325 ( .A(n_287), .Y(n_325) );
BUFx2_ASAP7_75t_L g326 ( .A(n_281), .Y(n_326) );
INVx1_ASAP7_75t_SL g327 ( .A(n_293), .Y(n_327) );
OAI21x1_ASAP7_75t_SL g328 ( .A1(n_273), .A2(n_213), .B(n_141), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_265), .B(n_221), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_296), .Y(n_330) );
OAI21x1_ASAP7_75t_L g331 ( .A1(n_285), .A2(n_170), .B(n_254), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_304), .B(n_207), .Y(n_332) );
OAI21xp5_ASAP7_75t_L g333 ( .A1(n_303), .A2(n_255), .B(n_208), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_277), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_275), .Y(n_335) );
AO21x2_ASAP7_75t_L g336 ( .A1(n_285), .A2(n_255), .B(n_229), .Y(n_336) );
OA21x2_ASAP7_75t_L g337 ( .A1(n_300), .A2(n_208), .B(n_247), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_302), .Y(n_338) );
OA21x2_ASAP7_75t_L g339 ( .A1(n_300), .A2(n_247), .B(n_236), .Y(n_339) );
A2O1A1Ixp33_ASAP7_75t_L g340 ( .A1(n_259), .A2(n_222), .B(n_240), .C(n_231), .Y(n_340) );
A2O1A1Ixp33_ASAP7_75t_L g341 ( .A1(n_312), .A2(n_259), .B(n_288), .C(n_290), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_332), .Y(n_342) );
NOR2xp67_ASAP7_75t_L g343 ( .A(n_316), .B(n_282), .Y(n_343) );
OR2x6_ASAP7_75t_L g344 ( .A(n_324), .B(n_272), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_312), .A2(n_267), .B1(n_221), .B2(n_276), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_310), .A2(n_303), .B(n_231), .Y(n_346) );
NAND2xp33_ASAP7_75t_R g347 ( .A(n_332), .B(n_271), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_318), .A2(n_221), .B1(n_305), .B2(n_279), .Y(n_348) );
OA21x2_ASAP7_75t_L g349 ( .A1(n_331), .A2(n_284), .B(n_283), .Y(n_349) );
AOI21xp33_ASAP7_75t_L g350 ( .A1(n_328), .A2(n_288), .B(n_295), .Y(n_350) );
OAI22xp33_ASAP7_75t_L g351 ( .A1(n_325), .A2(n_306), .B1(n_327), .B2(n_329), .Y(n_351) );
OAI22xp33_ASAP7_75t_L g352 ( .A1(n_325), .A2(n_221), .B1(n_289), .B2(n_299), .Y(n_352) );
BUFx4f_ASAP7_75t_SL g353 ( .A(n_327), .Y(n_353) );
INVx4_ASAP7_75t_L g354 ( .A(n_325), .Y(n_354) );
OAI211xp5_ASAP7_75t_L g355 ( .A1(n_329), .A2(n_301), .B(n_294), .C(n_264), .Y(n_355) );
AND2x4_ASAP7_75t_L g356 ( .A(n_324), .B(n_260), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_332), .B(n_270), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_330), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g359 ( .A1(n_318), .A2(n_292), .B1(n_297), .B2(n_141), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_330), .B(n_270), .Y(n_360) );
OAI22xp33_ASAP7_75t_L g361 ( .A1(n_326), .A2(n_213), .B1(n_292), .B2(n_291), .Y(n_361) );
OAI22xp33_ASAP7_75t_L g362 ( .A1(n_326), .A2(n_298), .B1(n_291), .B2(n_275), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_309), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_337), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_337), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_326), .A2(n_328), .B1(n_324), .B2(n_317), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_309), .Y(n_367) );
AOI222xp33_ASAP7_75t_L g368 ( .A1(n_317), .A2(n_141), .B1(n_286), .B2(n_291), .C1(n_275), .C2(n_298), .Y(n_368) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_353), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_347), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_363), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_342), .B(n_334), .Y(n_372) );
INVx3_ASAP7_75t_L g373 ( .A(n_364), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_364), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_357), .B(n_334), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_365), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_365), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_357), .B(n_321), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_363), .B(n_321), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_358), .B(n_310), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_367), .B(n_340), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_360), .B(n_321), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_360), .Y(n_383) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_354), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_351), .B(n_310), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_366), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_345), .B(n_321), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_349), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_356), .B(n_321), .Y(n_389) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_354), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_341), .B(n_340), .Y(n_391) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_354), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_348), .B(n_324), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_349), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_356), .B(n_338), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_349), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_344), .Y(n_397) );
BUFx2_ASAP7_75t_L g398 ( .A(n_344), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_344), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_371), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_374), .B(n_344), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_378), .B(n_338), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_375), .B(n_338), .Y(n_403) );
INVx1_ASAP7_75t_SL g404 ( .A(n_384), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_374), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_375), .B(n_336), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_395), .B(n_336), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_395), .B(n_336), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_374), .B(n_341), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_378), .B(n_336), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_376), .B(n_336), .Y(n_411) );
BUFx3_ASAP7_75t_L g412 ( .A(n_373), .Y(n_412) );
INVxp67_ASAP7_75t_L g413 ( .A(n_370), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_383), .B(n_331), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_371), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_376), .B(n_352), .Y(n_416) );
OAI21x1_ASAP7_75t_L g417 ( .A1(n_391), .A2(n_331), .B(n_322), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_376), .B(n_361), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_386), .A2(n_350), .B1(n_328), .B2(n_356), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_383), .B(n_315), .Y(n_420) );
BUFx2_ASAP7_75t_L g421 ( .A(n_373), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_383), .B(n_315), .Y(n_422) );
OAI221xp5_ASAP7_75t_L g423 ( .A1(n_393), .A2(n_359), .B1(n_355), .B2(n_343), .C(n_319), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_386), .A2(n_324), .B1(n_319), .B2(n_315), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_379), .Y(n_425) );
INVx3_ASAP7_75t_L g426 ( .A(n_373), .Y(n_426) );
NAND2x1_ASAP7_75t_L g427 ( .A(n_373), .B(n_335), .Y(n_427) );
AND2x4_ASAP7_75t_L g428 ( .A(n_397), .B(n_322), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_377), .Y(n_429) );
OR2x6_ASAP7_75t_L g430 ( .A(n_398), .B(n_346), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_377), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_377), .B(n_315), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_379), .Y(n_433) );
BUFx3_ASAP7_75t_L g434 ( .A(n_390), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_380), .B(n_315), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_380), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_382), .B(n_339), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_382), .B(n_362), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_389), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_389), .B(n_339), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_387), .B(n_339), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_381), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_400), .Y(n_443) );
NAND2x1p5_ASAP7_75t_L g444 ( .A(n_434), .B(n_398), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_404), .B(n_397), .Y(n_445) );
NOR3xp33_ASAP7_75t_SL g446 ( .A(n_423), .B(n_391), .C(n_372), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_436), .B(n_385), .Y(n_447) );
AND2x4_ASAP7_75t_L g448 ( .A(n_434), .B(n_397), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_404), .B(n_399), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_439), .B(n_399), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_400), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_415), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_415), .Y(n_453) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_436), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_413), .B(n_392), .Y(n_455) );
NAND3xp33_ASAP7_75t_L g456 ( .A(n_413), .B(n_369), .C(n_385), .Y(n_456) );
AOI221x1_ASAP7_75t_L g457 ( .A1(n_442), .A2(n_394), .B1(n_388), .B2(n_399), .C(n_387), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_434), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_439), .B(n_394), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_405), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_425), .B(n_6), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_425), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_433), .B(n_388), .Y(n_463) );
OAI211xp5_ASAP7_75t_SL g464 ( .A1(n_423), .A2(n_368), .B(n_396), .C(n_313), .Y(n_464) );
INVx3_ASAP7_75t_L g465 ( .A(n_412), .Y(n_465) );
INVxp67_ASAP7_75t_SL g466 ( .A(n_405), .Y(n_466) );
AND2x4_ASAP7_75t_L g467 ( .A(n_433), .B(n_396), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_403), .B(n_396), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_402), .B(n_9), .Y(n_469) );
NAND2x1p5_ASAP7_75t_L g470 ( .A(n_427), .B(n_323), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_405), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_403), .B(n_10), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_402), .B(n_10), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_442), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_402), .B(n_11), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_440), .B(n_11), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_440), .B(n_12), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_429), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_437), .B(n_12), .Y(n_479) );
INVxp67_ASAP7_75t_SL g480 ( .A(n_429), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_437), .B(n_14), .Y(n_481) );
INVx2_ASAP7_75t_SL g482 ( .A(n_412), .Y(n_482) );
INVxp67_ASAP7_75t_L g483 ( .A(n_421), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_406), .B(n_15), .Y(n_484) );
AND2x4_ASAP7_75t_L g485 ( .A(n_412), .B(n_322), .Y(n_485) );
AND2x4_ASAP7_75t_L g486 ( .A(n_401), .B(n_320), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_406), .B(n_15), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_429), .Y(n_488) );
NAND5xp2_ASAP7_75t_L g489 ( .A(n_419), .B(n_313), .C(n_284), .D(n_333), .E(n_16), .Y(n_489) );
INVx3_ASAP7_75t_L g490 ( .A(n_427), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_431), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_438), .B(n_17), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_438), .B(n_339), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_410), .B(n_339), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_431), .Y(n_495) );
OR2x6_ASAP7_75t_SL g496 ( .A(n_418), .B(n_270), .Y(n_496) );
NOR3xp33_ASAP7_75t_L g497 ( .A(n_418), .B(n_335), .C(n_308), .Y(n_497) );
NAND3xp33_ASAP7_75t_L g498 ( .A(n_419), .B(n_335), .C(n_308), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_431), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_443), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_451), .Y(n_501) );
NAND3xp33_ASAP7_75t_L g502 ( .A(n_456), .B(n_424), .C(n_430), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_445), .B(n_407), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_454), .B(n_401), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_462), .B(n_410), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_484), .B(n_408), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_452), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_460), .Y(n_508) );
NAND2xp33_ASAP7_75t_SL g509 ( .A(n_446), .B(n_421), .Y(n_509) );
INVxp67_ASAP7_75t_L g510 ( .A(n_454), .Y(n_510) );
INVx4_ASAP7_75t_L g511 ( .A(n_444), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_460), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_453), .Y(n_513) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_466), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_449), .B(n_407), .Y(n_515) );
OAI21xp5_ASAP7_75t_SL g516 ( .A1(n_461), .A2(n_424), .B(n_416), .Y(n_516) );
INVxp67_ASAP7_75t_SL g517 ( .A(n_466), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_447), .B(n_408), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_474), .B(n_441), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_455), .Y(n_520) );
INVx1_ASAP7_75t_SL g521 ( .A(n_476), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_455), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_494), .B(n_411), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_492), .B(n_409), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_463), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_493), .B(n_411), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_450), .B(n_441), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_459), .B(n_426), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_477), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_479), .Y(n_530) );
INVx2_ASAP7_75t_SL g531 ( .A(n_444), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_481), .Y(n_532) );
OR2x6_ASAP7_75t_L g533 ( .A(n_482), .B(n_430), .Y(n_533) );
OR2x6_ASAP7_75t_L g534 ( .A(n_490), .B(n_430), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_471), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_467), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_458), .B(n_426), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_473), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_475), .B(n_426), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_448), .B(n_426), .Y(n_540) );
AOI22xp33_ASAP7_75t_SL g541 ( .A1(n_461), .A2(n_416), .B1(n_414), .B2(n_428), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_467), .Y(n_542) );
NAND2x1p5_ASAP7_75t_L g543 ( .A(n_469), .B(n_323), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_487), .B(n_422), .Y(n_544) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_446), .A2(n_435), .B(n_409), .C(n_428), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_467), .Y(n_546) );
AND2x4_ASAP7_75t_L g547 ( .A(n_465), .B(n_430), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_448), .B(n_422), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_478), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_471), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_472), .B(n_420), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_489), .B(n_435), .Y(n_552) );
OAI21xp5_ASAP7_75t_L g553 ( .A1(n_498), .A2(n_417), .B(n_432), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_495), .Y(n_554) );
OAI21xp33_ASAP7_75t_L g555 ( .A1(n_483), .A2(n_430), .B(n_420), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_488), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_509), .A2(n_480), .B(n_497), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_500), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_516), .A2(n_497), .B1(n_486), .B2(n_464), .Y(n_559) );
OAI21xp33_ASAP7_75t_L g560 ( .A1(n_541), .A2(n_483), .B(n_464), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_514), .Y(n_561) );
AOI21xp33_ASAP7_75t_L g562 ( .A1(n_502), .A2(n_490), .B(n_485), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_509), .A2(n_480), .B(n_457), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_525), .B(n_491), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_552), .A2(n_541), .B1(n_524), .B2(n_520), .Y(n_565) );
CKINVDCx14_ASAP7_75t_R g566 ( .A(n_527), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_501), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_503), .B(n_465), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_552), .A2(n_486), .B1(n_485), .B2(n_428), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_507), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_518), .B(n_468), .Y(n_571) );
AOI222xp33_ASAP7_75t_L g572 ( .A1(n_524), .A2(n_486), .B1(n_485), .B2(n_414), .C1(n_428), .C2(n_432), .Y(n_572) );
A2O1A1Ixp33_ASAP7_75t_L g573 ( .A1(n_545), .A2(n_496), .B(n_499), .C(n_495), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_522), .A2(n_499), .B1(n_470), .B2(n_417), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_521), .B(n_470), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_513), .Y(n_576) );
OAI222xp33_ASAP7_75t_L g577 ( .A1(n_538), .A2(n_308), .B1(n_335), .B2(n_417), .C1(n_323), .C2(n_270), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_529), .A2(n_335), .B1(n_308), .B2(n_314), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_510), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_545), .A2(n_337), .B(n_308), .Y(n_580) );
AOI22x1_ASAP7_75t_SL g581 ( .A1(n_511), .A2(n_21), .B1(n_23), .B2(n_24), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_510), .Y(n_582) );
XNOR2xp5_ASAP7_75t_L g583 ( .A(n_551), .B(n_314), .Y(n_583) );
NOR4xp25_ASAP7_75t_SL g584 ( .A(n_517), .B(n_25), .C(n_26), .D(n_28), .Y(n_584) );
OAI322xp33_ASAP7_75t_L g585 ( .A1(n_530), .A2(n_311), .A3(n_254), .B1(n_231), .B2(n_240), .C1(n_307), .C2(n_314), .Y(n_585) );
INVxp67_ASAP7_75t_L g586 ( .A(n_504), .Y(n_586) );
OAI22xp33_ASAP7_75t_L g587 ( .A1(n_511), .A2(n_311), .B1(n_337), .B2(n_333), .Y(n_587) );
INVx1_ASAP7_75t_SL g588 ( .A(n_528), .Y(n_588) );
NOR2xp67_ASAP7_75t_L g589 ( .A(n_514), .B(n_29), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_532), .A2(n_337), .B1(n_307), .B2(n_320), .Y(n_590) );
INVx3_ASAP7_75t_SL g591 ( .A(n_531), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_506), .B(n_505), .Y(n_592) );
INVxp67_ASAP7_75t_L g593 ( .A(n_537), .Y(n_593) );
OAI21xp33_ASAP7_75t_SL g594 ( .A1(n_517), .A2(n_320), .B(n_307), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_508), .Y(n_595) );
OAI21xp5_ASAP7_75t_SL g596 ( .A1(n_543), .A2(n_311), .B(n_298), .Y(n_596) );
NOR4xp25_ASAP7_75t_SL g597 ( .A(n_555), .B(n_31), .C(n_36), .D(n_38), .Y(n_597) );
OAI211xp5_ASAP7_75t_L g598 ( .A1(n_553), .A2(n_311), .B(n_254), .C(n_240), .Y(n_598) );
OAI221xp5_ASAP7_75t_L g599 ( .A1(n_543), .A2(n_311), .B1(n_240), .B2(n_231), .C(n_43), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_579), .B(n_556), .Y(n_600) );
AOI211xp5_ASAP7_75t_L g601 ( .A1(n_591), .A2(n_547), .B(n_544), .C(n_539), .Y(n_601) );
INVxp67_ASAP7_75t_L g602 ( .A(n_582), .Y(n_602) );
O2A1O1Ixp33_ASAP7_75t_L g603 ( .A1(n_562), .A2(n_534), .B(n_519), .C(n_533), .Y(n_603) );
INVxp67_ASAP7_75t_SL g604 ( .A(n_561), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_564), .Y(n_605) );
NOR4xp25_ASAP7_75t_L g606 ( .A(n_565), .B(n_536), .C(n_542), .D(n_546), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_564), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_558), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_567), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_566), .A2(n_533), .B1(n_534), .B2(n_547), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_570), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g612 ( .A1(n_573), .A2(n_534), .B(n_533), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_592), .B(n_515), .Y(n_613) );
OAI221xp5_ASAP7_75t_L g614 ( .A1(n_560), .A2(n_526), .B1(n_523), .B2(n_549), .C(n_512), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_586), .B(n_547), .Y(n_615) );
OAI211xp5_ASAP7_75t_SL g616 ( .A1(n_562), .A2(n_559), .B(n_569), .C(n_572), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_576), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_571), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_575), .A2(n_548), .B1(n_512), .B2(n_508), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_595), .B(n_554), .Y(n_620) );
NOR3xp33_ASAP7_75t_SL g621 ( .A(n_577), .B(n_599), .C(n_557), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_568), .Y(n_622) );
NAND2xp33_ASAP7_75t_SL g623 ( .A(n_597), .B(n_540), .Y(n_623) );
XOR2x2_ASAP7_75t_L g624 ( .A(n_588), .B(n_39), .Y(n_624) );
XOR2x2_ASAP7_75t_L g625 ( .A(n_589), .B(n_40), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_605), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_607), .B(n_593), .Y(n_627) );
AOI222xp33_ASAP7_75t_L g628 ( .A1(n_616), .A2(n_583), .B1(n_594), .B2(n_587), .C1(n_578), .C2(n_599), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_606), .B(n_602), .Y(n_629) );
INVx3_ASAP7_75t_L g630 ( .A(n_624), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_618), .B(n_574), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_610), .A2(n_557), .B(n_563), .Y(n_632) );
OAI21xp33_ASAP7_75t_L g633 ( .A1(n_621), .A2(n_598), .B(n_596), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_600), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_615), .B(n_535), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_601), .B(n_535), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_608), .B(n_554), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_609), .B(n_550), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_600), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_623), .A2(n_581), .B1(n_550), .B2(n_590), .Y(n_640) );
INVx1_ASAP7_75t_SL g641 ( .A(n_625), .Y(n_641) );
AOI322xp5_ASAP7_75t_L g642 ( .A1(n_629), .A2(n_613), .A3(n_622), .B1(n_604), .B2(n_617), .C1(n_611), .C2(n_620), .Y(n_642) );
AOI211xp5_ASAP7_75t_L g643 ( .A1(n_633), .A2(n_603), .B(n_614), .C(n_612), .Y(n_643) );
AOI32xp33_ASAP7_75t_L g644 ( .A1(n_641), .A2(n_619), .A3(n_620), .B1(n_584), .B2(n_585), .Y(n_644) );
AOI211xp5_ASAP7_75t_L g645 ( .A1(n_632), .A2(n_580), .B(n_311), .C(n_51), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_627), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g647 ( .A1(n_631), .A2(n_311), .B1(n_236), .B2(n_210), .C(n_54), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_634), .A2(n_210), .B1(n_47), .B2(n_53), .C(n_55), .Y(n_648) );
OAI211xp5_ASAP7_75t_SL g649 ( .A1(n_628), .A2(n_42), .B(n_56), .C(n_60), .Y(n_649) );
OAI211xp5_ASAP7_75t_SL g650 ( .A1(n_640), .A2(n_61), .B(n_64), .C(n_69), .Y(n_650) );
NAND4xp75_ASAP7_75t_L g651 ( .A(n_644), .B(n_646), .C(n_649), .D(n_647), .Y(n_651) );
OAI222xp33_ASAP7_75t_L g652 ( .A1(n_643), .A2(n_630), .B1(n_636), .B2(n_627), .C1(n_639), .C2(n_626), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_642), .B(n_630), .Y(n_653) );
AND2x4_ASAP7_75t_L g654 ( .A(n_650), .B(n_635), .Y(n_654) );
OAI31xp33_ASAP7_75t_L g655 ( .A1(n_645), .A2(n_638), .A3(n_637), .B(n_78), .Y(n_655) );
NOR3xp33_ASAP7_75t_SL g656 ( .A(n_652), .B(n_648), .C(n_638), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_653), .Y(n_657) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_651), .Y(n_658) );
AOI21x1_ASAP7_75t_L g659 ( .A1(n_658), .A2(n_654), .B(n_655), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_657), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_660), .Y(n_661) );
OAI31xp33_ASAP7_75t_SL g662 ( .A1(n_659), .A2(n_657), .A3(n_656), .B(n_654), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_661), .Y(n_663) );
OAI321xp33_ASAP7_75t_L g664 ( .A1(n_663), .A2(n_662), .A3(n_72), .B1(n_70), .B2(n_226), .C(n_218), .Y(n_664) );
AOI322xp5_ASAP7_75t_L g665 ( .A1(n_664), .A2(n_218), .A3(n_226), .B1(n_658), .B2(n_657), .C1(n_663), .C2(n_660), .Y(n_665) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_665), .A2(n_218), .B(n_226), .Y(n_666) );
endmodule