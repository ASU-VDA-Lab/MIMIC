module real_jpeg_7444_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_0),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_0),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_0),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_0),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_0),
.B(n_269),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_0),
.B(n_311),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_0),
.B(n_290),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_0),
.B(n_390),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_1),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_1),
.B(n_76),
.Y(n_180)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_1),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_1),
.B(n_276),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_1),
.B(n_311),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_1),
.B(n_328),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_1),
.B(n_392),
.Y(n_391)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_2),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_2),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_2),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_3),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_3),
.Y(n_104)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_3),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_3),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_3),
.Y(n_208)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_3),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_4),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_4),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_4),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_4),
.B(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_4),
.B(n_166),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g213 ( 
.A(n_4),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_5),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_5),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_5),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_5),
.B(n_320),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_5),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_5),
.B(n_367),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_5),
.B(n_382),
.Y(n_381)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_6),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_6),
.Y(n_118)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_6),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g175 ( 
.A(n_6),
.Y(n_175)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_7),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_8),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_8),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_8),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_8),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_8),
.B(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_9),
.Y(n_274)
);

BUFx5_ASAP7_75t_L g296 ( 
.A(n_9),
.Y(n_296)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_11),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_11),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_12),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_12),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_12),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_12),
.B(n_294),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_12),
.B(n_309),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_12),
.B(n_266),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_12),
.B(n_362),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_12),
.B(n_82),
.Y(n_388)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_14),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_15),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_15),
.B(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_15),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_15),
.B(n_143),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_15),
.B(n_196),
.Y(n_195)
);

AND2x2_ASAP7_75t_SL g265 ( 
.A(n_15),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_15),
.B(n_311),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_15),
.B(n_211),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_16),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_16),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_16),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_16),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_16),
.B(n_253),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_16),
.B(n_272),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_16),
.B(n_214),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_17),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_17),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_17),
.B(n_290),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_17),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_17),
.B(n_333),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_17),
.B(n_369),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_17),
.B(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_18),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_18),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_18),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_18),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_18),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_18),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_18),
.B(n_241),
.Y(n_240)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_474),
.B(n_477),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_182),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_181),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_152),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_25),
.B(n_152),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_108),
.B2(n_151),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_74),
.C(n_89),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_28),
.B(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_47),
.C(n_62),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_29),
.B(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_34),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_30),
.B(n_36),
.C(n_40),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_32),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_32),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_32),
.Y(n_367)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_33),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_33),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_40),
.B2(n_46),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_35),
.A2(n_36),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_35),
.B(n_112),
.C(n_115),
.Y(n_133)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_39),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_40),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_40),
.B(n_92),
.C(n_96),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_40),
.A2(n_46),
.B1(n_96),
.B2(n_97),
.Y(n_161)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_44),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_47),
.B(n_62),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_53),
.C(n_57),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_48),
.B(n_57),
.Y(n_168)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_51),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_51),
.Y(n_369)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_52),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_53),
.B(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_56),
.Y(n_266)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_60),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_60),
.Y(n_392)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_61),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_61),
.Y(n_321)
);

BUFx5_ASAP7_75t_L g334 ( 
.A(n_61),
.Y(n_334)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_61),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_71),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_64),
.B(n_67),
.C(n_71),
.Y(n_120)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_74),
.A2(n_89),
.B1(n_90),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_75),
.B(n_78),
.C(n_88),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_88),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_100),
.C(n_105),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_91),
.B(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_92),
.B(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_96),
.A2(n_97),
.B1(n_165),
.B2(n_202),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_97),
.B(n_163),
.C(n_165),
.Y(n_162)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_99),
.Y(n_215)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_99),
.Y(n_241)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_99),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_100),
.A2(n_101),
.B1(n_105),
.B2(n_106),
.Y(n_170)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_105),
.A2(n_106),
.B1(n_179),
.B2(n_180),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_106),
.B(n_172),
.C(n_179),
.Y(n_171)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_121),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_119),
.C(n_120),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_115),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_113),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_120),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_132),
.B2(n_150),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_131),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_126),
.Y(n_194)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_127),
.Y(n_250)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_127),
.Y(n_382)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_148),
.B2(n_149),
.Y(n_132)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_139),
.B1(n_140),
.B2(n_147),
.Y(n_134)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_144),
.B(n_255),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_146),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.C(n_158),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_153),
.B(n_156),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_158),
.B(n_470),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_169),
.C(n_171),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_159),
.B(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.C(n_167),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_160),
.B(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_162),
.B(n_167),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_201),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_165),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_169),
.B(n_171),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_204),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.C(n_178),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_178),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_176),
.B(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AO21x1_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_467),
.B(n_472),
.Y(n_182)
);

OAI21x1_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_278),
.B(n_466),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_226),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_185),
.B(n_226),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_221),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_186),
.B(n_222),
.C(n_224),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_203),
.C(n_205),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_187),
.B(n_229),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.C(n_200),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_188),
.B(n_451),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_190),
.A2(n_191),
.B1(n_200),
.B2(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.C(n_198),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_192),
.B(n_198),
.Y(n_441)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_195),
.B(n_441),
.Y(n_440)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_200),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_205),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_216),
.C(n_219),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_206),
.B(n_258),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.C(n_213),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_207),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_213),
.Y(n_238)
);

BUFx8_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx5_ASAP7_75t_L g253 ( 
.A(n_212),
.Y(n_253)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_216),
.B(n_219),
.Y(n_258)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_230),
.C(n_233),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_228),
.B(n_231),
.Y(n_461)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_233),
.B(n_461),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_256),
.C(n_259),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_235),
.B(n_454),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.C(n_246),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_236),
.A2(n_237),
.B1(n_432),
.B2(n_433),
.Y(n_431)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_239),
.A2(n_240),
.B(n_242),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_239),
.B(n_246),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

MAJx2_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_251),
.C(n_254),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_247),
.A2(n_248),
.B1(n_251),
.B2(n_252),
.Y(n_409)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_254),
.B(n_409),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_255),
.B(n_350),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g454 ( 
.A1(n_256),
.A2(n_257),
.B1(n_259),
.B2(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_259),
.Y(n_455)
);

MAJx2_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_271),
.C(n_275),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_261),
.B(n_443),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.C(n_267),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_262),
.B(n_421),
.Y(n_420)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_265),
.A2(n_267),
.B1(n_268),
.B2(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_265),
.Y(n_422)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_271),
.B(n_275),
.Y(n_443)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx8_ASAP7_75t_L g390 ( 
.A(n_273),
.Y(n_390)
);

BUFx5_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_274),
.Y(n_317)
);

INVx4_ASAP7_75t_L g380 ( 
.A(n_276),
.Y(n_380)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

AOI21x1_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_459),
.B(n_465),
.Y(n_278)
);

OAI21x1_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_446),
.B(n_458),
.Y(n_279)
);

AOI21x1_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_428),
.B(n_445),
.Y(n_280)
);

OAI21x1_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_402),
.B(n_427),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_373),
.B(n_401),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_342),
.B(n_372),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_323),
.B(n_341),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_303),
.B(n_322),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_297),
.B(n_302),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_295),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_295),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_293),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_298),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_293),
.Y(n_304)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_292),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_292),
.Y(n_328)
);

INVx4_ASAP7_75t_SL g350 ( 
.A(n_296),
.Y(n_350)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_305),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_312),
.B2(n_313),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_306),
.B(n_315),
.C(n_318),
.Y(n_340)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_310),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_308),
.B(n_310),
.Y(n_330)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_318),
.B2(n_319),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_340),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_324),
.B(n_340),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_331),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_330),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_326),
.B(n_330),
.C(n_344),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_329),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_327),
.B(n_329),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_331),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_335),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_332),
.B(n_358),
.C(n_359),
.Y(n_357)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_339),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_336),
.Y(n_358)
);

INVx6_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_339),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_345),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_343),
.B(n_345),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_356),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_346),
.B(n_357),
.C(n_360),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_347),
.B(n_349),
.C(n_351),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_351),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_352),
.A2(n_353),
.B1(n_354),
.B2(n_355),
.Y(n_351)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_352),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_353),
.B(n_355),
.Y(n_383)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_360),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_365),
.Y(n_360)
);

MAJx2_ASAP7_75t_L g399 ( 
.A(n_361),
.B(n_368),
.C(n_370),
.Y(n_399)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_366),
.A2(n_368),
.B1(n_370),
.B2(n_371),
.Y(n_365)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_366),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_368),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_374),
.B(n_400),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_374),
.B(n_400),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_375),
.B(n_385),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_384),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_376),
.B(n_384),
.C(n_426),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_383),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_381),
.Y(n_377)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_378),
.Y(n_416)
);

INVx5_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_381),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_383),
.B(n_416),
.C(n_417),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_385),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_393),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_386),
.B(n_395),
.C(n_398),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_391),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

MAJx2_ASAP7_75t_L g413 ( 
.A(n_388),
.B(n_389),
.C(n_391),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_394),
.A2(n_395),
.B1(n_398),
.B2(n_399),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_396),
.B(n_397),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_399),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_425),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_403),
.B(n_425),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_414),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_406),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_405),
.B(n_406),
.C(n_414),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_407),
.A2(n_408),
.B1(n_410),
.B2(n_411),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_407),
.B(n_437),
.C(n_438),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_413),
.Y(n_411)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_412),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_413),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_SL g414 ( 
.A(n_415),
.B(n_418),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_415),
.B(n_419),
.C(n_424),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_419),
.A2(n_420),
.B1(n_423),
.B2(n_424),
.Y(n_418)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_419),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_420),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_429),
.B(n_444),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_429),
.B(n_444),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_430),
.B(n_435),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_434),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_431),
.B(n_434),
.C(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_432),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_435),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_436),
.B(n_439),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_436),
.B(n_440),
.C(n_442),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_442),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_447),
.B(n_456),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_447),
.B(n_456),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_449),
.Y(n_447)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_448),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_453),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_450),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_453),
.B(n_463),
.C(n_464),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_460),
.B(n_462),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_460),
.B(n_462),
.Y(n_465)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_469),
.B(n_471),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_469),
.B(n_471),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

BUFx12f_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx5_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx13_ASAP7_75t_L g479 ( 
.A(n_476),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_480),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);


endmodule