module fake_netlist_6_497_n_2111 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_507, n_580, n_209, n_367, n_465, n_590, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_557, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_555, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_522, n_466, n_506, n_56, n_360, n_119, n_235, n_536, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_581, n_428, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_323, n_393, n_411, n_503, n_152, n_92, n_513, n_321, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_95, n_311, n_10, n_403, n_253, n_583, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_560, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_582, n_4, n_199, n_138, n_266, n_296, n_571, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2111);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_590;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_557;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_536;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_583;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_560;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_571;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2111;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_1380;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1930;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_830;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_699;
wire n_1986;
wire n_824;
wire n_686;
wire n_757;
wire n_1641;
wire n_1918;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_1970;
wire n_608;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2073;
wire n_792;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_2031;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_702;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_851;
wire n_644;
wire n_682;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_765;
wire n_1492;
wire n_987;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_2069;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_683;
wire n_811;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_889;
wire n_1478;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_1440;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_1993;
wire n_1427;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_1060;
wire n_1951;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_1520;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_1731;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_613;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2016;
wire n_1905;
wire n_793;
wire n_1593;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_607;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_952;
wire n_725;
wire n_999;
wire n_1254;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_1997;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2037;
wire n_782;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1640;
wire n_804;
wire n_1846;
wire n_806;
wire n_879;
wire n_959;
wire n_1343;
wire n_1522;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_652;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_1373;
wire n_1292;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_672;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_655;
wire n_1045;
wire n_706;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1949;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1929;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_1848;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_1922;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_1276;
wire n_2015;
wire n_1148;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_924;
wire n_1582;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_1218;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_985;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_1996;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_849;
wire n_753;
wire n_1753;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_2091;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_1025;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_316),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_39),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_292),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_534),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_76),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_74),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_128),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_105),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_191),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_181),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_275),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_393),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_78),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_283),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_550),
.Y(n_609)
);

BUFx2_ASAP7_75t_L g610 ( 
.A(n_496),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_242),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_527),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_190),
.Y(n_613)
);

BUFx10_ASAP7_75t_L g614 ( 
.A(n_580),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_570),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_532),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_195),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_290),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_92),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_298),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_343),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_22),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_83),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_15),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_471),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_399),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_20),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_431),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_308),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_554),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_141),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_581),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_196),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_237),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_374),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_592),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_335),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_578),
.Y(n_638)
);

HB1xp67_ASAP7_75t_L g639 ( 
.A(n_81),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_338),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_461),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_543),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_224),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_587),
.Y(n_644)
);

BUFx10_ASAP7_75t_L g645 ( 
.A(n_280),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_526),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_110),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_129),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_133),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_390),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_502),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_225),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_186),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_328),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_428),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_498),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_81),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_146),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_382),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_282),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_56),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_545),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_388),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_312),
.Y(n_664)
);

BUFx10_ASAP7_75t_L g665 ( 
.A(n_232),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_500),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_159),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_58),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_175),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_401),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_152),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_572),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_99),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_495),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_28),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_172),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_408),
.Y(n_677)
);

BUFx2_ASAP7_75t_SL g678 ( 
.A(n_453),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_14),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_229),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_208),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_266),
.Y(n_682)
);

BUFx8_ASAP7_75t_SL g683 ( 
.A(n_557),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_56),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_560),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_12),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_192),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_273),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_499),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_482),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_67),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_515),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_173),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_78),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_454),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_586),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_504),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_188),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_381),
.Y(n_699)
);

CKINVDCx16_ASAP7_75t_R g700 ( 
.A(n_370),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_100),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_121),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_248),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_575),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_304),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_246),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_555),
.Y(n_707)
);

BUFx2_ASAP7_75t_L g708 ( 
.A(n_429),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_562),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_513),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_549),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_569),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_288),
.Y(n_713)
);

CKINVDCx20_ASAP7_75t_R g714 ( 
.A(n_577),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_334),
.Y(n_715)
);

CKINVDCx16_ASAP7_75t_R g716 ( 
.A(n_548),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_62),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_244),
.Y(n_718)
);

CKINVDCx16_ASAP7_75t_R g719 ( 
.A(n_536),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_300),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_394),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_62),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_327),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_573),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_377),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_583),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_341),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_241),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_472),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_187),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_508),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_574),
.Y(n_732)
);

INVx1_ASAP7_75t_SL g733 ( 
.A(n_77),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_530),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_74),
.Y(n_735)
);

CKINVDCx20_ASAP7_75t_R g736 ( 
.A(n_143),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_144),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_520),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_439),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_269),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_571),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_591),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_497),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_485),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_391),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_50),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_329),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_271),
.Y(n_748)
);

CKINVDCx20_ASAP7_75t_R g749 ( 
.A(n_579),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_50),
.Y(n_750)
);

BUFx2_ASAP7_75t_R g751 ( 
.A(n_470),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_293),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_262),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_22),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_210),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_94),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_193),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_72),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_325),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_576),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_245),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_228),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_568),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_128),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_315),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_363),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_417),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_220),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_161),
.Y(n_769)
);

CKINVDCx20_ASAP7_75t_R g770 ( 
.A(n_364),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_622),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_683),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_622),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_622),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_623),
.Y(n_775)
);

BUFx2_ASAP7_75t_L g776 ( 
.A(n_639),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_668),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_673),
.Y(n_778)
);

CKINVDCx20_ASAP7_75t_R g779 ( 
.A(n_629),
.Y(n_779)
);

CKINVDCx20_ASAP7_75t_R g780 ( 
.A(n_664),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_595),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_702),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_735),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_692),
.Y(n_784)
);

CKINVDCx20_ASAP7_75t_R g785 ( 
.A(n_696),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_714),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_750),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_754),
.Y(n_788)
);

BUFx2_ASAP7_75t_L g789 ( 
.A(n_596),
.Y(n_789)
);

CKINVDCx16_ASAP7_75t_R g790 ( 
.A(n_700),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_600),
.Y(n_791)
);

BUFx2_ASAP7_75t_SL g792 ( 
.A(n_718),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_647),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_603),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_608),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_615),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_618),
.Y(n_797)
);

INVxp67_ASAP7_75t_SL g798 ( 
.A(n_756),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_637),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_642),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_653),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_680),
.Y(n_802)
);

INVxp33_ASAP7_75t_SL g803 ( 
.A(n_599),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_681),
.Y(n_804)
);

BUFx10_ASAP7_75t_L g805 ( 
.A(n_601),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_687),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_597),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_695),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_697),
.Y(n_809)
);

INVxp67_ASAP7_75t_L g810 ( 
.A(n_758),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_698),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_709),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_598),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_713),
.Y(n_814)
);

CKINVDCx16_ASAP7_75t_R g815 ( 
.A(n_716),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_721),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_726),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_604),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_605),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_606),
.Y(n_820)
);

CKINVDCx16_ASAP7_75t_R g821 ( 
.A(n_719),
.Y(n_821)
);

CKINVDCx16_ASAP7_75t_R g822 ( 
.A(n_736),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_729),
.Y(n_823)
);

CKINVDCx16_ASAP7_75t_R g824 ( 
.A(n_749),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_731),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_734),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_742),
.Y(n_827)
);

INVxp33_ASAP7_75t_SL g828 ( 
.A(n_602),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_748),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_755),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_761),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_609),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_765),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_733),
.Y(n_834)
);

HB1xp67_ASAP7_75t_L g835 ( 
.A(n_619),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_766),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_612),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_688),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_723),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_611),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_613),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_614),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_621),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_616),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_651),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_636),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_720),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_617),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_732),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_636),
.Y(n_850)
);

INVx1_ASAP7_75t_SL g851 ( 
.A(n_607),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_610),
.B(n_0),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_614),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_620),
.Y(n_854)
);

CKINVDCx16_ASAP7_75t_R g855 ( 
.A(n_770),
.Y(n_855)
);

INVxp67_ASAP7_75t_SL g856 ( 
.A(n_636),
.Y(n_856)
);

INVxp33_ASAP7_75t_SL g857 ( 
.A(n_624),
.Y(n_857)
);

INVxp33_ASAP7_75t_SL g858 ( 
.A(n_627),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_753),
.Y(n_859)
);

CKINVDCx20_ASAP7_75t_R g860 ( 
.A(n_625),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_646),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_646),
.Y(n_862)
);

INVxp67_ASAP7_75t_SL g863 ( 
.A(n_646),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_656),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_656),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_656),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_739),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_739),
.Y(n_868)
);

INVxp33_ASAP7_75t_L g869 ( 
.A(n_708),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_739),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_768),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_781),
.B(n_807),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_846),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_856),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_805),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_834),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_842),
.B(n_659),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_856),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_846),
.Y(n_879)
);

AND2x6_ASAP7_75t_L g880 ( 
.A(n_843),
.B(n_768),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_863),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_846),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_863),
.Y(n_883)
);

OAI22x1_ASAP7_75t_SL g884 ( 
.A1(n_851),
.A2(n_649),
.B1(n_657),
.B2(n_648),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_850),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_771),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_773),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_774),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_861),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_868),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_813),
.Y(n_891)
);

OA21x2_ASAP7_75t_L g892 ( 
.A1(n_794),
.A2(n_740),
.B(n_677),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_862),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_835),
.B(n_869),
.Y(n_894)
);

INVx4_ASAP7_75t_L g895 ( 
.A(n_818),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_790),
.B(n_645),
.Y(n_896)
);

OA21x2_ASAP7_75t_L g897 ( 
.A1(n_795),
.A2(n_743),
.B(n_628),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_864),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_865),
.Y(n_899)
);

BUFx12f_ASAP7_75t_L g900 ( 
.A(n_772),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_866),
.Y(n_901)
);

NOR2x1_ASAP7_75t_L g902 ( 
.A(n_842),
.B(n_678),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_867),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_L g904 ( 
.A1(n_834),
.A2(n_675),
.B1(n_679),
.B2(n_661),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_870),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_859),
.B(n_737),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_871),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_775),
.Y(n_908)
);

OAI21x1_ASAP7_75t_L g909 ( 
.A1(n_796),
.A2(n_799),
.B(n_797),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_815),
.A2(n_686),
.B1(n_691),
.B2(n_684),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_821),
.B(n_645),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_788),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_803),
.B(n_665),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_791),
.Y(n_914)
);

AOI22x1_ASAP7_75t_SL g915 ( 
.A1(n_779),
.A2(n_701),
.B1(n_717),
.B2(n_694),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_800),
.Y(n_916)
);

OA22x2_ASAP7_75t_SL g917 ( 
.A1(n_798),
.A2(n_751),
.B1(n_2),
.B2(n_0),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_819),
.B(n_747),
.Y(n_918)
);

OA21x2_ASAP7_75t_L g919 ( 
.A1(n_801),
.A2(n_804),
.B(n_802),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_828),
.B(n_665),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_853),
.B(n_768),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_777),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_820),
.B(n_832),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_782),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_SL g925 ( 
.A1(n_822),
.A2(n_746),
.B1(n_764),
.B2(n_722),
.Y(n_925)
);

BUFx8_ASAP7_75t_L g926 ( 
.A(n_789),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_837),
.B(n_626),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_806),
.Y(n_928)
);

CKINVDCx20_ASAP7_75t_R g929 ( 
.A(n_780),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_840),
.B(n_760),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_841),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_808),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_783),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_809),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_844),
.B(n_762),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_811),
.Y(n_936)
);

BUFx8_ASAP7_75t_L g937 ( 
.A(n_776),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_787),
.Y(n_938)
);

CKINVDCx6p67_ASAP7_75t_R g939 ( 
.A(n_792),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_812),
.Y(n_940)
);

OA21x2_ASAP7_75t_L g941 ( 
.A1(n_814),
.A2(n_631),
.B(n_630),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_845),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_838),
.B(n_632),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_816),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_852),
.A2(n_634),
.B1(n_635),
.B2(n_633),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_839),
.Y(n_946)
);

OA21x2_ASAP7_75t_L g947 ( 
.A1(n_817),
.A2(n_640),
.B(n_638),
.Y(n_947)
);

OA22x2_ASAP7_75t_L g948 ( 
.A1(n_778),
.A2(n_810),
.B1(n_798),
.B2(n_793),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_848),
.B(n_730),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_805),
.Y(n_950)
);

BUFx2_ASAP7_75t_L g951 ( 
.A(n_854),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_823),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_825),
.Y(n_953)
);

AND2x6_ASAP7_75t_L g954 ( 
.A(n_847),
.B(n_135),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_826),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_849),
.Y(n_956)
);

NAND2xp33_ASAP7_75t_L g957 ( 
.A(n_778),
.B(n_641),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_885),
.Y(n_958)
);

AOI21x1_ASAP7_75t_L g959 ( 
.A1(n_916),
.A2(n_829),
.B(n_827),
.Y(n_959)
);

CKINVDCx6p67_ASAP7_75t_R g960 ( 
.A(n_900),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_874),
.B(n_830),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_877),
.B(n_857),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_921),
.B(n_878),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_881),
.B(n_858),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_877),
.B(n_643),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_885),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_873),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_882),
.Y(n_968)
);

NOR2x1p5_ASAP7_75t_L g969 ( 
.A(n_950),
.B(n_644),
.Y(n_969)
);

INVx2_ASAP7_75t_SL g970 ( 
.A(n_894),
.Y(n_970)
);

INVx11_ASAP7_75t_L g971 ( 
.A(n_926),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_928),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_902),
.B(n_650),
.Y(n_973)
);

AO21x2_ASAP7_75t_L g974 ( 
.A1(n_918),
.A2(n_833),
.B(n_831),
.Y(n_974)
);

AND3x2_ASAP7_75t_L g975 ( 
.A(n_876),
.B(n_810),
.C(n_793),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_914),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_932),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_890),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_879),
.Y(n_979)
);

INVx1_ASAP7_75t_SL g980 ( 
.A(n_929),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_934),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_906),
.B(n_652),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_879),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_912),
.Y(n_984)
);

NAND3xp33_ASAP7_75t_L g985 ( 
.A(n_897),
.B(n_836),
.C(n_655),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_936),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_883),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_901),
.Y(n_988)
);

INVx2_ASAP7_75t_SL g989 ( 
.A(n_943),
.Y(n_989)
);

XOR2xp5_ASAP7_75t_L g990 ( 
.A(n_915),
.B(n_784),
.Y(n_990)
);

OR2x6_ASAP7_75t_L g991 ( 
.A(n_875),
.B(n_824),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_908),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_903),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_906),
.B(n_654),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_919),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_907),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_944),
.Y(n_997)
);

AND3x2_ASAP7_75t_L g998 ( 
.A(n_913),
.B(n_9),
.C(n_1),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_908),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_937),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_952),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_951),
.B(n_921),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_945),
.B(n_658),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_886),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_940),
.Y(n_1005)
);

INVxp67_ASAP7_75t_SL g1006 ( 
.A(n_919),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_887),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_888),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_889),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_940),
.Y(n_1010)
);

NAND3xp33_ASAP7_75t_L g1011 ( 
.A(n_897),
.B(n_662),
.C(n_660),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_927),
.B(n_663),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_953),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_951),
.B(n_860),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_892),
.B(n_666),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_953),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_955),
.Y(n_1017)
);

INVx4_ASAP7_75t_L g1018 ( 
.A(n_955),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_893),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_933),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_909),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_898),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_933),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_899),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_922),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_924),
.Y(n_1026)
);

NOR2x1p5_ASAP7_75t_L g1027 ( 
.A(n_939),
.B(n_667),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_927),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_905),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_956),
.Y(n_1030)
);

INVx2_ASAP7_75t_SL g1031 ( 
.A(n_948),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_938),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_946),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_930),
.B(n_669),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_942),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_920),
.B(n_670),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_942),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_892),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_941),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_941),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_947),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_947),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_880),
.Y(n_1043)
);

AOI21x1_ASAP7_75t_L g1044 ( 
.A1(n_935),
.A2(n_672),
.B(n_671),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_891),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_949),
.B(n_674),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_880),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_957),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_880),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_954),
.Y(n_1050)
);

OR2x2_ASAP7_75t_L g1051 ( 
.A(n_910),
.B(n_855),
.Y(n_1051)
);

XNOR2x1_ASAP7_75t_L g1052 ( 
.A(n_990),
.B(n_904),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_970),
.B(n_931),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_972),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_977),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_981),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_1035),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_1002),
.B(n_923),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_986),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_997),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1001),
.Y(n_1061)
);

INVx2_ASAP7_75t_SL g1062 ( 
.A(n_999),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_1045),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_964),
.B(n_872),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1037),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_984),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_976),
.Y(n_1067)
);

NAND2xp33_ASAP7_75t_R g1068 ( 
.A(n_1051),
.B(n_915),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_978),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_958),
.B(n_966),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_1030),
.Y(n_1071)
);

INVxp33_ASAP7_75t_SL g1072 ( 
.A(n_1045),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1025),
.Y(n_1073)
);

NOR2xp67_ASAP7_75t_L g1074 ( 
.A(n_1011),
.B(n_895),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1026),
.Y(n_1075)
);

INVx1_ASAP7_75t_SL g1076 ( 
.A(n_980),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_964),
.B(n_1036),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1032),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_1036),
.B(n_896),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_987),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_988),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_1014),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_993),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_996),
.Y(n_1084)
);

NAND2xp33_ASAP7_75t_R g1085 ( 
.A(n_975),
.B(n_676),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1034),
.B(n_954),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_963),
.Y(n_1087)
);

BUFx3_ASAP7_75t_L g1088 ( 
.A(n_1020),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_963),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1004),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_1007),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1008),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1009),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_SL g1094 ( 
.A(n_991),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1019),
.Y(n_1095)
);

INVxp33_ASAP7_75t_L g1096 ( 
.A(n_962),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1022),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1024),
.Y(n_1098)
);

INVxp33_ASAP7_75t_SL g1099 ( 
.A(n_980),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_989),
.B(n_785),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1029),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_967),
.Y(n_1102)
);

CKINVDCx20_ASAP7_75t_R g1103 ( 
.A(n_960),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_SL g1104 ( 
.A(n_998),
.B(n_954),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_968),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_1048),
.B(n_911),
.Y(n_1106)
);

NOR2xp67_ASAP7_75t_L g1107 ( 
.A(n_1011),
.B(n_136),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_971),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_1018),
.B(n_786),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_961),
.Y(n_1110)
);

INVx4_ASAP7_75t_L g1111 ( 
.A(n_1020),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_961),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1033),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1005),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_979),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1010),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1013),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1016),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1006),
.A2(n_685),
.B(n_682),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1017),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_982),
.B(n_925),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1023),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_959),
.Y(n_1123)
);

XNOR2xp5_ASAP7_75t_L g1124 ( 
.A(n_1027),
.B(n_884),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1018),
.B(n_689),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_983),
.Y(n_1126)
);

INVxp67_ASAP7_75t_SL g1127 ( 
.A(n_992),
.Y(n_1127)
);

XOR2xp5_ASAP7_75t_L g1128 ( 
.A(n_1000),
.B(n_690),
.Y(n_1128)
);

INVx2_ASAP7_75t_SL g1129 ( 
.A(n_958),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1020),
.B(n_693),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_966),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_992),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1028),
.B(n_699),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_991),
.Y(n_1134)
);

CKINVDCx20_ASAP7_75t_R g1135 ( 
.A(n_991),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_992),
.Y(n_1136)
);

XOR2xp5_ASAP7_75t_L g1137 ( 
.A(n_985),
.B(n_703),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1006),
.Y(n_1138)
);

INVx1_ASAP7_75t_SL g1139 ( 
.A(n_975),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1021),
.Y(n_1140)
);

CKINVDCx20_ASAP7_75t_R g1141 ( 
.A(n_1046),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1038),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_995),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_982),
.B(n_926),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_995),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1015),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1015),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_962),
.B(n_994),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_994),
.B(n_704),
.Y(n_1149)
);

AND2x6_ASAP7_75t_SL g1150 ( 
.A(n_1034),
.B(n_917),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_1077),
.B(n_1046),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_1063),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1110),
.B(n_974),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_1064),
.B(n_1003),
.Y(n_1154)
);

INVx2_ASAP7_75t_SL g1155 ( 
.A(n_1053),
.Y(n_1155)
);

OAI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1143),
.A2(n_1041),
.B(n_1039),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1142),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1058),
.B(n_1112),
.Y(n_1158)
);

AND2x6_ASAP7_75t_SL g1159 ( 
.A(n_1121),
.B(n_998),
.Y(n_1159)
);

INVxp67_ASAP7_75t_L g1160 ( 
.A(n_1100),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_1072),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_1091),
.Y(n_1162)
);

NOR3xp33_ASAP7_75t_L g1163 ( 
.A(n_1079),
.B(n_1003),
.C(n_1012),
.Y(n_1163)
);

BUFx4_ASAP7_75t_L g1164 ( 
.A(n_1099),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1146),
.B(n_974),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1054),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1055),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_1106),
.B(n_1031),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1145),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1056),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_SL g1171 ( 
.A(n_1104),
.B(n_1144),
.Y(n_1171)
);

OAI221xp5_ASAP7_75t_L g1172 ( 
.A1(n_1137),
.A2(n_1012),
.B1(n_965),
.B2(n_985),
.C(n_973),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1147),
.B(n_1138),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1066),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1059),
.B(n_1040),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1067),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1060),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_1148),
.B(n_973),
.Y(n_1178)
);

OR2x6_ASAP7_75t_SL g1179 ( 
.A(n_1108),
.B(n_705),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1071),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1061),
.Y(n_1181)
);

AND2x6_ASAP7_75t_SL g1182 ( 
.A(n_1109),
.B(n_937),
.Y(n_1182)
);

NOR3xp33_ASAP7_75t_L g1183 ( 
.A(n_1082),
.B(n_965),
.C(n_1044),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1057),
.B(n_1065),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1069),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1087),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1089),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1096),
.B(n_1042),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_1080),
.B(n_1049),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1149),
.B(n_1050),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1073),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_1074),
.B(n_1049),
.Y(n_1192)
);

NOR3xp33_ASAP7_75t_L g1193 ( 
.A(n_1082),
.B(n_1076),
.C(n_1139),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1150),
.B(n_1139),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1074),
.B(n_1043),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1133),
.B(n_1130),
.Y(n_1196)
);

AND2x2_ASAP7_75t_SL g1197 ( 
.A(n_1104),
.B(n_1047),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_1088),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1081),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1107),
.A2(n_969),
.B1(n_707),
.B2(n_710),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1075),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1140),
.B(n_706),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1078),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1141),
.B(n_711),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1083),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1084),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1111),
.B(n_712),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1102),
.Y(n_1208)
);

NAND2xp33_ASAP7_75t_L g1209 ( 
.A(n_1086),
.B(n_715),
.Y(n_1209)
);

BUFx3_ASAP7_75t_L g1210 ( 
.A(n_1103),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1125),
.B(n_724),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1090),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1123),
.B(n_725),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1092),
.B(n_727),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_1070),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1093),
.B(n_728),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1150),
.B(n_738),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1095),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1097),
.B(n_741),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1113),
.B(n_744),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1132),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1098),
.Y(n_1222)
);

INVx2_ASAP7_75t_SL g1223 ( 
.A(n_1070),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1101),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1114),
.B(n_745),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_1111),
.B(n_752),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1105),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1116),
.B(n_757),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1117),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1107),
.A2(n_763),
.B1(n_767),
.B2(n_759),
.Y(n_1230)
);

BUFx4f_ASAP7_75t_L g1231 ( 
.A(n_1198),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1158),
.B(n_1119),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1157),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1169),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_R g1235 ( 
.A(n_1161),
.B(n_1068),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_1152),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1154),
.B(n_1052),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1174),
.Y(n_1238)
);

INVx2_ASAP7_75t_SL g1239 ( 
.A(n_1155),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1160),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1196),
.B(n_1127),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_1198),
.Y(n_1242)
);

NOR3xp33_ASAP7_75t_SL g1243 ( 
.A(n_1194),
.B(n_1085),
.C(n_1124),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1166),
.Y(n_1244)
);

INVx2_ASAP7_75t_SL g1245 ( 
.A(n_1164),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1176),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1180),
.Y(n_1247)
);

BUFx4f_ASAP7_75t_L g1248 ( 
.A(n_1198),
.Y(n_1248)
);

OR2x2_ASAP7_75t_SL g1249 ( 
.A(n_1159),
.B(n_1118),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1163),
.B(n_1062),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1191),
.Y(n_1251)
);

BUFx3_ASAP7_75t_L g1252 ( 
.A(n_1210),
.Y(n_1252)
);

INVx5_ASAP7_75t_L g1253 ( 
.A(n_1215),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_R g1254 ( 
.A(n_1171),
.B(n_1134),
.Y(n_1254)
);

NOR3xp33_ASAP7_75t_SL g1255 ( 
.A(n_1217),
.B(n_769),
.C(n_1136),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1182),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_1179),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1201),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_R g1259 ( 
.A(n_1171),
.B(n_1135),
.Y(n_1259)
);

AOI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1151),
.A2(n_1122),
.B1(n_1120),
.B2(n_1131),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1167),
.Y(n_1261)
);

INVx3_ASAP7_75t_L g1262 ( 
.A(n_1215),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1172),
.A2(n_1126),
.B1(n_1129),
.B2(n_1115),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_R g1264 ( 
.A(n_1159),
.B(n_1094),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1173),
.A2(n_1094),
.B1(n_1128),
.B2(n_138),
.Y(n_1265)
);

BUFx3_ASAP7_75t_L g1266 ( 
.A(n_1223),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1170),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_1197),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1203),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1177),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1221),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1168),
.B(n_1),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1153),
.B(n_2),
.Y(n_1273)
);

AND2x4_ASAP7_75t_SL g1274 ( 
.A(n_1193),
.B(n_137),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1199),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1181),
.Y(n_1276)
);

AND2x4_ASAP7_75t_L g1277 ( 
.A(n_1186),
.B(n_139),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1187),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1229),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1188),
.B(n_3),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_1182),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_1190),
.B(n_140),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1208),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1212),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_1162),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1165),
.B(n_3),
.Y(n_1286)
);

BUFx3_ASAP7_75t_L g1287 ( 
.A(n_1218),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1211),
.B(n_4),
.Y(n_1288)
);

INVx2_ASAP7_75t_SL g1289 ( 
.A(n_1227),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1162),
.Y(n_1290)
);

NAND2xp33_ASAP7_75t_R g1291 ( 
.A(n_1175),
.B(n_142),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1204),
.B(n_4),
.Y(n_1292)
);

AOI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1183),
.A2(n_147),
.B1(n_148),
.B2(n_145),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1185),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_1184),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1222),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1224),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1205),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1206),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1213),
.Y(n_1300)
);

BUFx2_ASAP7_75t_L g1301 ( 
.A(n_1214),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1178),
.B(n_1202),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1213),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1202),
.B(n_5),
.Y(n_1304)
);

BUFx4f_ASAP7_75t_L g1305 ( 
.A(n_1207),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1302),
.A2(n_1156),
.B(n_1195),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1300),
.B(n_1220),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_SL g1308 ( 
.A1(n_1232),
.A2(n_1192),
.B(n_1156),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1303),
.A2(n_1209),
.B(n_1226),
.Y(n_1309)
);

BUFx4f_ASAP7_75t_L g1310 ( 
.A(n_1242),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1241),
.A2(n_1200),
.B(n_1216),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1250),
.A2(n_1219),
.B(n_1189),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1282),
.A2(n_1230),
.B(n_1228),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1273),
.A2(n_1225),
.B(n_150),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1286),
.A2(n_151),
.B(n_149),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_1231),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1301),
.A2(n_154),
.B(n_153),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1301),
.B(n_5),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1268),
.B(n_6),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1237),
.B(n_6),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1260),
.A2(n_156),
.B(n_155),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1268),
.B(n_7),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1248),
.Y(n_1323)
);

AO31x2_ASAP7_75t_L g1324 ( 
.A1(n_1280),
.A2(n_158),
.A3(n_160),
.B(n_157),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1288),
.A2(n_163),
.B(n_162),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1263),
.A2(n_165),
.B(n_164),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1240),
.Y(n_1327)
);

AOI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1304),
.A2(n_167),
.B(n_166),
.Y(n_1328)
);

NAND2x1p5_ASAP7_75t_L g1329 ( 
.A(n_1242),
.B(n_168),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1268),
.B(n_7),
.Y(n_1330)
);

AND2x6_ASAP7_75t_SL g1331 ( 
.A(n_1292),
.B(n_8),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1252),
.Y(n_1332)
);

AOI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1244),
.A2(n_170),
.B(n_169),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1233),
.A2(n_174),
.B(n_171),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1272),
.B(n_8),
.Y(n_1335)
);

INVx3_ASAP7_75t_L g1336 ( 
.A(n_1236),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1295),
.B(n_9),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1275),
.A2(n_177),
.B(n_176),
.Y(n_1338)
);

INVx2_ASAP7_75t_SL g1339 ( 
.A(n_1240),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1283),
.A2(n_179),
.B(n_178),
.Y(n_1340)
);

AO31x2_ASAP7_75t_L g1341 ( 
.A1(n_1261),
.A2(n_182),
.A3(n_183),
.B(n_180),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1234),
.A2(n_185),
.B(n_184),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1262),
.A2(n_194),
.B(n_189),
.Y(n_1343)
);

CKINVDCx11_ASAP7_75t_R g1344 ( 
.A(n_1257),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1295),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_1345)
);

O2A1O1Ixp5_ASAP7_75t_L g1346 ( 
.A1(n_1305),
.A2(n_13),
.B(n_10),
.C(n_11),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1284),
.B(n_13),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1251),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1258),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1287),
.B(n_14),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1254),
.B(n_15),
.Y(n_1351)
);

BUFx4f_ASAP7_75t_L g1352 ( 
.A(n_1245),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1294),
.A2(n_198),
.B(n_197),
.Y(n_1353)
);

BUFx8_ASAP7_75t_L g1354 ( 
.A(n_1239),
.Y(n_1354)
);

AO31x2_ASAP7_75t_L g1355 ( 
.A1(n_1267),
.A2(n_200),
.A3(n_201),
.B(n_199),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1238),
.A2(n_203),
.B(n_202),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1266),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1297),
.B(n_16),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1295),
.B(n_16),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_L g1360 ( 
.A(n_1299),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_SL g1361 ( 
.A1(n_1293),
.A2(n_205),
.B(n_204),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1269),
.B(n_17),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1270),
.B(n_17),
.Y(n_1363)
);

INVx1_ASAP7_75t_SL g1364 ( 
.A(n_1271),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1246),
.A2(n_207),
.B(n_206),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1249),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1276),
.B(n_18),
.Y(n_1367)
);

BUFx3_ASAP7_75t_L g1368 ( 
.A(n_1285),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1279),
.B(n_18),
.Y(n_1369)
);

OAI22x1_ASAP7_75t_L g1370 ( 
.A1(n_1277),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_SL g1371 ( 
.A(n_1259),
.B(n_19),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_SL g1372 ( 
.A(n_1296),
.B(n_21),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1247),
.A2(n_211),
.B(n_209),
.Y(n_1373)
);

BUFx2_ASAP7_75t_L g1374 ( 
.A(n_1298),
.Y(n_1374)
);

INVx2_ASAP7_75t_SL g1375 ( 
.A(n_1235),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1253),
.A2(n_213),
.B(n_212),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1243),
.B(n_23),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1296),
.B(n_23),
.Y(n_1378)
);

OAI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1278),
.A2(n_215),
.B(n_214),
.Y(n_1379)
);

OAI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1289),
.A2(n_217),
.B(n_216),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1253),
.A2(n_219),
.B(n_218),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1296),
.Y(n_1382)
);

A2O1A1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1277),
.A2(n_26),
.B(n_24),
.C(n_25),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1348),
.Y(n_1384)
);

AO21x1_ASAP7_75t_L g1385 ( 
.A1(n_1335),
.A2(n_1291),
.B(n_1265),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1320),
.B(n_1274),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1321),
.A2(n_1255),
.B(n_1253),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1314),
.A2(n_1290),
.B(n_1285),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1311),
.A2(n_1290),
.B(n_1285),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1327),
.Y(n_1390)
);

OAI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1307),
.A2(n_1281),
.B(n_1256),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1364),
.B(n_1290),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1306),
.A2(n_222),
.B(n_221),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1349),
.Y(n_1394)
);

BUFx10_ASAP7_75t_L g1395 ( 
.A(n_1323),
.Y(n_1395)
);

AO31x2_ASAP7_75t_L g1396 ( 
.A1(n_1309),
.A2(n_1312),
.A3(n_1315),
.B(n_1325),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1356),
.A2(n_226),
.B(n_223),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_SL g1398 ( 
.A1(n_1379),
.A2(n_1264),
.B(n_230),
.Y(n_1398)
);

AO21x1_ASAP7_75t_L g1399 ( 
.A1(n_1380),
.A2(n_24),
.B(n_25),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1374),
.B(n_26),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1308),
.A2(n_594),
.B(n_231),
.Y(n_1401)
);

NAND2x1p5_ASAP7_75t_L g1402 ( 
.A(n_1336),
.B(n_227),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1362),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1377),
.B(n_27),
.Y(n_1404)
);

INVx3_ASAP7_75t_L g1405 ( 
.A(n_1332),
.Y(n_1405)
);

OAI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1313),
.A2(n_27),
.B(n_28),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1317),
.A2(n_234),
.B(n_233),
.Y(n_1407)
);

BUFx10_ASAP7_75t_L g1408 ( 
.A(n_1323),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1374),
.B(n_29),
.Y(n_1409)
);

A2O1A1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1383),
.A2(n_31),
.B(n_29),
.C(n_30),
.Y(n_1410)
);

INVx3_ASAP7_75t_L g1411 ( 
.A(n_1357),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_SL g1412 ( 
.A(n_1352),
.B(n_1375),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1365),
.A2(n_236),
.B(n_235),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_SL g1414 ( 
.A(n_1310),
.B(n_238),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1319),
.B(n_30),
.Y(n_1415)
);

O2A1O1Ixp33_ASAP7_75t_SL g1416 ( 
.A1(n_1372),
.A2(n_33),
.B(n_31),
.C(n_32),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1327),
.B(n_32),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1339),
.B(n_33),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1363),
.Y(n_1419)
);

AO31x2_ASAP7_75t_L g1420 ( 
.A1(n_1370),
.A2(n_240),
.A3(n_243),
.B(n_239),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1318),
.B(n_34),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1360),
.B(n_34),
.Y(n_1422)
);

A2O1A1Ixp33_ASAP7_75t_L g1423 ( 
.A1(n_1326),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1322),
.B(n_35),
.Y(n_1424)
);

A2O1A1Ixp33_ASAP7_75t_L g1425 ( 
.A1(n_1346),
.A2(n_38),
.B(n_36),
.C(n_37),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_SL g1426 ( 
.A(n_1360),
.B(n_38),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1351),
.B(n_247),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1373),
.A2(n_250),
.B(n_249),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1376),
.A2(n_593),
.B(n_252),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1367),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1334),
.A2(n_1340),
.B(n_1338),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1381),
.A2(n_590),
.B(n_253),
.Y(n_1432)
);

AO31x2_ASAP7_75t_L g1433 ( 
.A1(n_1345),
.A2(n_254),
.A3(n_255),
.B(n_251),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1330),
.B(n_39),
.Y(n_1434)
);

O2A1O1Ixp33_ASAP7_75t_L g1435 ( 
.A1(n_1371),
.A2(n_42),
.B(n_40),
.C(n_41),
.Y(n_1435)
);

INVxp67_ASAP7_75t_L g1436 ( 
.A(n_1357),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1316),
.Y(n_1437)
);

BUFx2_ASAP7_75t_L g1438 ( 
.A(n_1354),
.Y(n_1438)
);

A2O1A1Ixp33_ASAP7_75t_L g1439 ( 
.A1(n_1378),
.A2(n_42),
.B(n_40),
.C(n_41),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1369),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1342),
.A2(n_257),
.B(n_256),
.Y(n_1441)
);

AOI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1366),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_1368),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1361),
.A2(n_259),
.B(n_258),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1361),
.A2(n_1343),
.B(n_1353),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1337),
.A2(n_261),
.B(n_260),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1333),
.A2(n_264),
.B(n_263),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1359),
.B(n_43),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1382),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1328),
.A2(n_267),
.B(n_265),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1328),
.A2(n_270),
.B(n_268),
.Y(n_1451)
);

OAI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1347),
.A2(n_44),
.B(n_45),
.Y(n_1452)
);

AOI221x1_ASAP7_75t_L g1453 ( 
.A1(n_1350),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.C(n_49),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1358),
.A2(n_1329),
.B1(n_1331),
.B2(n_1344),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1324),
.Y(n_1455)
);

BUFx2_ASAP7_75t_L g1456 ( 
.A(n_1324),
.Y(n_1456)
);

AO32x2_ASAP7_75t_L g1457 ( 
.A1(n_1341),
.A2(n_48),
.A3(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_1457)
);

AOI221x1_ASAP7_75t_L g1458 ( 
.A1(n_1341),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.C(n_54),
.Y(n_1458)
);

BUFx6f_ASAP7_75t_SL g1459 ( 
.A(n_1355),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1355),
.B(n_51),
.Y(n_1460)
);

AOI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1311),
.A2(n_274),
.B(n_272),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1307),
.B(n_276),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1348),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1348),
.Y(n_1464)
);

A2O1A1Ixp33_ASAP7_75t_L g1465 ( 
.A1(n_1307),
.A2(n_54),
.B(n_52),
.C(n_53),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1332),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1311),
.A2(n_278),
.B(n_277),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_SL g1468 ( 
.A(n_1323),
.B(n_279),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1307),
.B(n_55),
.Y(n_1469)
);

OAI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1311),
.A2(n_55),
.B(n_57),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1311),
.A2(n_284),
.B(n_281),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1311),
.A2(n_286),
.B(n_285),
.Y(n_1472)
);

BUFx2_ASAP7_75t_L g1473 ( 
.A(n_1327),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1348),
.Y(n_1474)
);

CKINVDCx20_ASAP7_75t_R g1475 ( 
.A(n_1344),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1348),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_1344),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1415),
.B(n_287),
.Y(n_1478)
);

CKINVDCx11_ASAP7_75t_R g1479 ( 
.A(n_1475),
.Y(n_1479)
);

BUFx12f_ASAP7_75t_L g1480 ( 
.A(n_1395),
.Y(n_1480)
);

AOI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1385),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1390),
.B(n_289),
.Y(n_1482)
);

INVx5_ASAP7_75t_L g1483 ( 
.A(n_1443),
.Y(n_1483)
);

INVx4_ASAP7_75t_L g1484 ( 
.A(n_1437),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1452),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1384),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_SL g1487 ( 
.A1(n_1470),
.A2(n_63),
.B1(n_60),
.B2(n_61),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_SL g1488 ( 
.A1(n_1454),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_1473),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1394),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1474),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1427),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1463),
.Y(n_1493)
);

INVx1_ASAP7_75t_SL g1494 ( 
.A(n_1405),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1464),
.Y(n_1495)
);

CKINVDCx6p67_ASAP7_75t_R g1496 ( 
.A(n_1408),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1399),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1443),
.Y(n_1498)
);

AOI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1386),
.A2(n_1462),
.B1(n_1419),
.B2(n_1440),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_SL g1500 ( 
.A1(n_1460),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_1500)
);

OAI22xp33_ASAP7_75t_SL g1501 ( 
.A1(n_1442),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1404),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1424),
.B(n_291),
.Y(n_1503)
);

INVxp67_ASAP7_75t_SL g1504 ( 
.A(n_1449),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1476),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1455),
.Y(n_1506)
);

AOI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1398),
.A2(n_295),
.B(n_294),
.Y(n_1507)
);

OAI21xp5_ASAP7_75t_SL g1508 ( 
.A1(n_1453),
.A2(n_73),
.B(n_75),
.Y(n_1508)
);

OAI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1414),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_1437),
.Y(n_1510)
);

CKINVDCx6p67_ASAP7_75t_R g1511 ( 
.A(n_1438),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1430),
.Y(n_1512)
);

OAI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1403),
.A2(n_82),
.B1(n_79),
.B2(n_80),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1469),
.B(n_79),
.Y(n_1514)
);

INVx6_ASAP7_75t_L g1515 ( 
.A(n_1417),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1391),
.A2(n_1422),
.B1(n_1426),
.B2(n_1434),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1457),
.Y(n_1517)
);

OAI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1468),
.A2(n_83),
.B1(n_80),
.B2(n_82),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1448),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1457),
.Y(n_1520)
);

CKINVDCx11_ASAP7_75t_R g1521 ( 
.A(n_1477),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1388),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1456),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1456),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1459),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1406),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_1411),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_SL g1528 ( 
.A1(n_1421),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_1528)
);

INVx1_ASAP7_75t_SL g1529 ( 
.A(n_1466),
.Y(n_1529)
);

INVx2_ASAP7_75t_SL g1530 ( 
.A(n_1392),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1444),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1450),
.Y(n_1532)
);

INVx6_ASAP7_75t_L g1533 ( 
.A(n_1418),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1451),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1400),
.B(n_90),
.Y(n_1535)
);

INVx6_ASAP7_75t_L g1536 ( 
.A(n_1412),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1409),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1446),
.A2(n_1407),
.B1(n_1472),
.B2(n_1471),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1458),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1467),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1439),
.B(n_1465),
.Y(n_1541)
);

INVx1_ASAP7_75t_SL g1542 ( 
.A(n_1389),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_SL g1543 ( 
.A1(n_1402),
.A2(n_94),
.B1(n_91),
.B2(n_93),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1420),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1401),
.A2(n_96),
.B1(n_93),
.B2(n_95),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1410),
.B(n_95),
.Y(n_1546)
);

INVx1_ASAP7_75t_SL g1547 ( 
.A(n_1436),
.Y(n_1547)
);

CKINVDCx11_ASAP7_75t_R g1548 ( 
.A(n_1416),
.Y(n_1548)
);

BUFx3_ASAP7_75t_L g1549 ( 
.A(n_1387),
.Y(n_1549)
);

INVx6_ASAP7_75t_L g1550 ( 
.A(n_1435),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_1429),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_SL g1552 ( 
.A1(n_1432),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1445),
.A2(n_1393),
.B1(n_1447),
.B2(n_1413),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1420),
.Y(n_1554)
);

CKINVDCx11_ASAP7_75t_R g1555 ( 
.A(n_1423),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1397),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1461),
.Y(n_1557)
);

OAI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1425),
.A2(n_102),
.B1(n_100),
.B2(n_101),
.Y(n_1558)
);

OAI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1431),
.A2(n_101),
.B(n_102),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1428),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.Y(n_1560)
);

CKINVDCx11_ASAP7_75t_R g1561 ( 
.A(n_1433),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1441),
.A2(n_106),
.B1(n_103),
.B2(n_104),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1433),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1396),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_SL g1565 ( 
.A1(n_1396),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1384),
.Y(n_1566)
);

BUFx2_ASAP7_75t_L g1567 ( 
.A(n_1390),
.Y(n_1567)
);

CKINVDCx11_ASAP7_75t_R g1568 ( 
.A(n_1475),
.Y(n_1568)
);

BUFx12f_ASAP7_75t_L g1569 ( 
.A(n_1395),
.Y(n_1569)
);

INVx8_ASAP7_75t_L g1570 ( 
.A(n_1443),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1384),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1384),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1490),
.Y(n_1573)
);

OA21x2_ASAP7_75t_L g1574 ( 
.A1(n_1563),
.A2(n_109),
.B(n_110),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1567),
.B(n_111),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1504),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1493),
.Y(n_1577)
);

BUFx2_ASAP7_75t_L g1578 ( 
.A(n_1525),
.Y(n_1578)
);

INVx2_ASAP7_75t_SL g1579 ( 
.A(n_1483),
.Y(n_1579)
);

OR2x6_ASAP7_75t_L g1580 ( 
.A(n_1536),
.B(n_296),
.Y(n_1580)
);

BUFx3_ASAP7_75t_L g1581 ( 
.A(n_1570),
.Y(n_1581)
);

NOR2x1_ASAP7_75t_L g1582 ( 
.A(n_1512),
.B(n_111),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1515),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1537),
.B(n_112),
.Y(n_1584)
);

OAI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1507),
.A2(n_1487),
.B(n_1508),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1506),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1495),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1524),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1523),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1505),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1486),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1489),
.B(n_112),
.Y(n_1592)
);

INVx4_ASAP7_75t_L g1593 ( 
.A(n_1483),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1499),
.B(n_113),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1491),
.Y(n_1595)
);

BUFx3_ASAP7_75t_L g1596 ( 
.A(n_1570),
.Y(n_1596)
);

OAI21x1_ASAP7_75t_L g1597 ( 
.A1(n_1553),
.A2(n_299),
.B(n_297),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1566),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1530),
.B(n_113),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_SL g1600 ( 
.A(n_1527),
.Y(n_1600)
);

OAI21x1_ASAP7_75t_L g1601 ( 
.A1(n_1557),
.A2(n_302),
.B(n_301),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1544),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1571),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1572),
.Y(n_1604)
);

INVx3_ASAP7_75t_L g1605 ( 
.A(n_1549),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1554),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1517),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1520),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1522),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1539),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1542),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1515),
.B(n_114),
.Y(n_1612)
);

AND2x6_ASAP7_75t_SL g1613 ( 
.A(n_1535),
.B(n_114),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1533),
.Y(n_1614)
);

INVx3_ASAP7_75t_L g1615 ( 
.A(n_1536),
.Y(n_1615)
);

BUFx6f_ASAP7_75t_L g1616 ( 
.A(n_1510),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1533),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1532),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_SL g1619 ( 
.A(n_1498),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1534),
.Y(n_1620)
);

OA21x2_ASAP7_75t_L g1621 ( 
.A1(n_1559),
.A2(n_115),
.B(n_116),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1516),
.B(n_115),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1561),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1546),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1514),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1482),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1481),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1482),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1494),
.B(n_116),
.Y(n_1629)
);

BUFx6f_ASAP7_75t_L g1630 ( 
.A(n_1510),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1541),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1550),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1478),
.B(n_117),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1550),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1529),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1513),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1547),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1565),
.Y(n_1638)
);

AOI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1538),
.A2(n_305),
.B(n_303),
.Y(n_1639)
);

INVx3_ASAP7_75t_L g1640 ( 
.A(n_1483),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1558),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1503),
.B(n_117),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1551),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1510),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1484),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1484),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1555),
.Y(n_1647)
);

AOI222xp33_ASAP7_75t_L g1648 ( 
.A1(n_1485),
.A2(n_1543),
.B1(n_1526),
.B2(n_1492),
.C1(n_1497),
.C2(n_1519),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1548),
.Y(n_1649)
);

INVx3_ASAP7_75t_L g1650 ( 
.A(n_1480),
.Y(n_1650)
);

INVx3_ASAP7_75t_L g1651 ( 
.A(n_1569),
.Y(n_1651)
);

OAI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1540),
.A2(n_307),
.B(n_306),
.Y(n_1652)
);

OR2x6_ASAP7_75t_L g1653 ( 
.A(n_1479),
.B(n_309),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1564),
.Y(n_1654)
);

BUFx2_ASAP7_75t_L g1655 ( 
.A(n_1511),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1501),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1552),
.Y(n_1657)
);

AO21x1_ASAP7_75t_SL g1658 ( 
.A1(n_1531),
.A2(n_118),
.B(n_119),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1500),
.B(n_118),
.Y(n_1659)
);

CKINVDCx20_ASAP7_75t_R g1660 ( 
.A(n_1568),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1556),
.B(n_119),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1488),
.B(n_120),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1560),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1562),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1528),
.Y(n_1665)
);

OAI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1545),
.A2(n_311),
.B(n_310),
.Y(n_1666)
);

OAI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1502),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1496),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1518),
.B(n_122),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1509),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1521),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1506),
.Y(n_1672)
);

AO21x1_ASAP7_75t_SL g1673 ( 
.A1(n_1517),
.A2(n_123),
.B(n_124),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1504),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1567),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1490),
.Y(n_1676)
);

INVx5_ASAP7_75t_L g1677 ( 
.A(n_1550),
.Y(n_1677)
);

OAI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1507),
.A2(n_314),
.B(n_313),
.Y(n_1678)
);

OR2x6_ASAP7_75t_L g1679 ( 
.A(n_1536),
.B(n_317),
.Y(n_1679)
);

OAI21x1_ASAP7_75t_L g1680 ( 
.A1(n_1553),
.A2(n_319),
.B(n_318),
.Y(n_1680)
);

INVxp67_ASAP7_75t_L g1681 ( 
.A(n_1567),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1490),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1490),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1573),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1675),
.B(n_123),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1577),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1623),
.B(n_124),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1589),
.Y(n_1688)
);

OAI21xp33_ASAP7_75t_SL g1689 ( 
.A1(n_1582),
.A2(n_125),
.B(n_126),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1583),
.B(n_125),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1672),
.Y(n_1691)
);

OA21x2_ASAP7_75t_L g1692 ( 
.A1(n_1610),
.A2(n_126),
.B(n_127),
.Y(n_1692)
);

AO21x2_ASAP7_75t_L g1693 ( 
.A1(n_1643),
.A2(n_127),
.B(n_129),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1672),
.Y(n_1694)
);

AND2x4_ASAP7_75t_L g1695 ( 
.A(n_1605),
.B(n_130),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1590),
.Y(n_1696)
);

HB1xp67_ASAP7_75t_L g1697 ( 
.A(n_1602),
.Y(n_1697)
);

HB1xp67_ASAP7_75t_L g1698 ( 
.A(n_1588),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1587),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1586),
.Y(n_1700)
);

INVx2_ASAP7_75t_SL g1701 ( 
.A(n_1616),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1681),
.B(n_1614),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1576),
.B(n_130),
.Y(n_1703)
);

BUFx2_ASAP7_75t_L g1704 ( 
.A(n_1578),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1676),
.Y(n_1705)
);

AO21x1_ASAP7_75t_SL g1706 ( 
.A1(n_1585),
.A2(n_131),
.B(n_132),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1606),
.Y(n_1707)
);

INVx3_ASAP7_75t_SL g1708 ( 
.A(n_1660),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1682),
.Y(n_1709)
);

AO21x2_ASAP7_75t_L g1710 ( 
.A1(n_1620),
.A2(n_131),
.B(n_132),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1617),
.B(n_133),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1683),
.Y(n_1712)
);

AO21x2_ASAP7_75t_L g1713 ( 
.A1(n_1609),
.A2(n_134),
.B(n_320),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1615),
.B(n_134),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1674),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1607),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1608),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1598),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1611),
.B(n_321),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1603),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1591),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1595),
.Y(n_1722)
);

INVx1_ASAP7_75t_SL g1723 ( 
.A(n_1632),
.Y(n_1723)
);

NOR2x1_ASAP7_75t_SL g1724 ( 
.A(n_1677),
.B(n_322),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1615),
.B(n_323),
.Y(n_1725)
);

OAI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1678),
.A2(n_324),
.B(n_326),
.Y(n_1726)
);

BUFx6f_ASAP7_75t_L g1727 ( 
.A(n_1616),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1647),
.B(n_330),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1604),
.Y(n_1729)
);

NAND2x1_ASAP7_75t_L g1730 ( 
.A(n_1605),
.B(n_331),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1618),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1627),
.A2(n_336),
.B1(n_332),
.B2(n_333),
.Y(n_1732)
);

OAI21x1_ASAP7_75t_L g1733 ( 
.A1(n_1597),
.A2(n_337),
.B(n_339),
.Y(n_1733)
);

BUFx2_ASAP7_75t_L g1734 ( 
.A(n_1640),
.Y(n_1734)
);

BUFx6f_ASAP7_75t_L g1735 ( 
.A(n_1616),
.Y(n_1735)
);

CKINVDCx20_ASAP7_75t_R g1736 ( 
.A(n_1655),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1574),
.Y(n_1737)
);

OAI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1652),
.A2(n_1666),
.B(n_1639),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1637),
.B(n_340),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1624),
.B(n_342),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1635),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1644),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1645),
.B(n_344),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1574),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1646),
.Y(n_1745)
);

OR2x6_ASAP7_75t_L g1746 ( 
.A(n_1580),
.B(n_345),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1625),
.B(n_346),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1634),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1656),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1631),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1584),
.Y(n_1751)
);

BUFx3_ASAP7_75t_L g1752 ( 
.A(n_1640),
.Y(n_1752)
);

AO21x2_ASAP7_75t_L g1753 ( 
.A1(n_1622),
.A2(n_347),
.B(n_348),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1621),
.Y(n_1754)
);

BUFx3_ASAP7_75t_L g1755 ( 
.A(n_1677),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1630),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1601),
.Y(n_1757)
);

HB1xp67_ASAP7_75t_L g1758 ( 
.A(n_1621),
.Y(n_1758)
);

BUFx2_ASAP7_75t_L g1759 ( 
.A(n_1593),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1677),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1707),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1707),
.Y(n_1762)
);

AND2x4_ASAP7_75t_L g1763 ( 
.A(n_1752),
.B(n_1579),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1716),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1717),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1723),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1738),
.A2(n_1648),
.B1(n_1654),
.B2(n_1657),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1723),
.Y(n_1768)
);

BUFx3_ASAP7_75t_L g1769 ( 
.A(n_1708),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1698),
.B(n_1592),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1704),
.B(n_1698),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1752),
.B(n_1760),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1734),
.B(n_1649),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1691),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1694),
.Y(n_1775)
);

INVx3_ASAP7_75t_L g1776 ( 
.A(n_1755),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1688),
.B(n_1629),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1688),
.B(n_1594),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1748),
.Y(n_1779)
);

INVx3_ASAP7_75t_L g1780 ( 
.A(n_1755),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1738),
.A2(n_1670),
.B1(n_1665),
.B2(n_1638),
.Y(n_1781)
);

HB1xp67_ASAP7_75t_L g1782 ( 
.A(n_1697),
.Y(n_1782)
);

AOI21xp5_ASAP7_75t_L g1783 ( 
.A1(n_1726),
.A2(n_1679),
.B(n_1580),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1760),
.B(n_1650),
.Y(n_1784)
);

OAI221xp5_ASAP7_75t_L g1785 ( 
.A1(n_1689),
.A2(n_1659),
.B1(n_1669),
.B2(n_1661),
.C(n_1662),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1749),
.B(n_1671),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1697),
.Y(n_1787)
);

NOR2x1_ASAP7_75t_L g1788 ( 
.A(n_1736),
.B(n_1668),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1702),
.B(n_1650),
.Y(n_1789)
);

NAND4xp25_ASAP7_75t_SL g1790 ( 
.A(n_1726),
.B(n_1613),
.C(n_1641),
.D(n_1633),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1684),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1715),
.B(n_1636),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1745),
.B(n_1651),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1684),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1699),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1700),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1754),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1741),
.B(n_1651),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1705),
.Y(n_1799)
);

HB1xp67_ASAP7_75t_L g1800 ( 
.A(n_1754),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1742),
.B(n_1575),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1709),
.Y(n_1802)
);

INVx2_ASAP7_75t_SL g1803 ( 
.A(n_1727),
.Y(n_1803)
);

AND2x4_ASAP7_75t_L g1804 ( 
.A(n_1759),
.B(n_1686),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1720),
.Y(n_1805)
);

BUFx3_ASAP7_75t_L g1806 ( 
.A(n_1708),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1718),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_SL g1808 ( 
.A(n_1758),
.B(n_1626),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1696),
.Y(n_1809)
);

BUFx2_ASAP7_75t_L g1810 ( 
.A(n_1756),
.Y(n_1810)
);

OAI211xp5_ASAP7_75t_L g1811 ( 
.A1(n_1758),
.A2(n_1692),
.B(n_1663),
.C(n_1664),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1712),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1721),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1722),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1729),
.B(n_1628),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1751),
.B(n_1612),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1731),
.B(n_1581),
.Y(n_1817)
);

HB1xp67_ASAP7_75t_L g1818 ( 
.A(n_1737),
.Y(n_1818)
);

AOI221xp5_ASAP7_75t_L g1819 ( 
.A1(n_1703),
.A2(n_1667),
.B1(n_1599),
.B2(n_1642),
.C(n_1596),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1731),
.Y(n_1820)
);

BUFx3_ASAP7_75t_L g1821 ( 
.A(n_1736),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1750),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1761),
.B(n_1762),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1771),
.B(n_1744),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1773),
.B(n_1701),
.Y(n_1825)
);

OR2x6_ASAP7_75t_L g1826 ( 
.A(n_1783),
.B(n_1746),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1782),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1782),
.B(n_1703),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1774),
.Y(n_1829)
);

NOR2x1_ASAP7_75t_SL g1830 ( 
.A(n_1808),
.B(n_1673),
.Y(n_1830)
);

BUFx2_ASAP7_75t_L g1831 ( 
.A(n_1788),
.Y(n_1831)
);

AOI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1783),
.A2(n_1746),
.B(n_1693),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1784),
.B(n_1776),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1775),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1818),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1818),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1804),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1787),
.Y(n_1838)
);

BUFx6f_ASAP7_75t_L g1839 ( 
.A(n_1806),
.Y(n_1839)
);

BUFx2_ASAP7_75t_L g1840 ( 
.A(n_1821),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1764),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1797),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1804),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1772),
.Y(n_1844)
);

AND2x4_ASAP7_75t_L g1845 ( 
.A(n_1784),
.B(n_1757),
.Y(n_1845)
);

BUFx8_ASAP7_75t_L g1846 ( 
.A(n_1806),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1777),
.B(n_1757),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1765),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1772),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1795),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1796),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1791),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1776),
.B(n_1685),
.Y(n_1853)
);

HB1xp67_ASAP7_75t_L g1854 ( 
.A(n_1797),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1794),
.Y(n_1855)
);

AOI322xp5_ASAP7_75t_L g1856 ( 
.A1(n_1767),
.A2(n_1687),
.A3(n_1690),
.B1(n_1714),
.B2(n_1695),
.C1(n_1740),
.C2(n_1711),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1800),
.B(n_1692),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1805),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1780),
.B(n_1695),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1820),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1780),
.B(n_1727),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1842),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1833),
.B(n_1786),
.Y(n_1863)
);

NOR2xp33_ASAP7_75t_L g1864 ( 
.A(n_1839),
.B(n_1769),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1844),
.B(n_1849),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1828),
.B(n_1770),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1831),
.B(n_1837),
.Y(n_1867)
);

OR2x2_ASAP7_75t_L g1868 ( 
.A(n_1828),
.B(n_1778),
.Y(n_1868)
);

OR2x2_ASAP7_75t_L g1869 ( 
.A(n_1847),
.B(n_1778),
.Y(n_1869)
);

AND2x4_ASAP7_75t_SL g1870 ( 
.A(n_1839),
.B(n_1746),
.Y(n_1870)
);

NOR2xp33_ASAP7_75t_L g1871 ( 
.A(n_1839),
.B(n_1821),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1842),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1829),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1843),
.B(n_1789),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1845),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1823),
.B(n_1792),
.Y(n_1876)
);

HB1xp67_ASAP7_75t_L g1877 ( 
.A(n_1854),
.Y(n_1877)
);

INVx5_ASAP7_75t_SL g1878 ( 
.A(n_1826),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1845),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1840),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1852),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1827),
.B(n_1800),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1861),
.B(n_1859),
.Y(n_1883)
);

AND2x4_ASAP7_75t_L g1884 ( 
.A(n_1826),
.B(n_1763),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1826),
.B(n_1853),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1855),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_L g1887 ( 
.A(n_1846),
.B(n_1790),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1824),
.B(n_1825),
.Y(n_1888)
);

AND2x4_ASAP7_75t_L g1889 ( 
.A(n_1830),
.B(n_1763),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1835),
.B(n_1822),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1834),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1823),
.B(n_1838),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1860),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1841),
.B(n_1793),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1848),
.B(n_1798),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1850),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1883),
.B(n_1817),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1866),
.B(n_1868),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1873),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1873),
.Y(n_1900)
);

OR2x2_ASAP7_75t_L g1901 ( 
.A(n_1880),
.B(n_1832),
.Y(n_1901)
);

OAI21xp33_ASAP7_75t_L g1902 ( 
.A1(n_1887),
.A2(n_1832),
.B(n_1767),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1894),
.B(n_1856),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1863),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1885),
.B(n_1810),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1878),
.B(n_1856),
.Y(n_1906)
);

INVx3_ASAP7_75t_L g1907 ( 
.A(n_1889),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1891),
.Y(n_1908)
);

HB1xp67_ASAP7_75t_L g1909 ( 
.A(n_1877),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1891),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1896),
.Y(n_1911)
);

NAND2x1p5_ASAP7_75t_L g1912 ( 
.A(n_1889),
.B(n_1593),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1896),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1862),
.Y(n_1914)
);

INVxp67_ASAP7_75t_L g1915 ( 
.A(n_1871),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1888),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1878),
.B(n_1801),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1867),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_L g1919 ( 
.A(n_1915),
.B(n_1864),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1909),
.B(n_1865),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1906),
.B(n_1895),
.Y(n_1921)
);

NOR2x1_ASAP7_75t_L g1922 ( 
.A(n_1907),
.B(n_1862),
.Y(n_1922)
);

INVxp33_ASAP7_75t_L g1923 ( 
.A(n_1917),
.Y(n_1923)
);

AOI22xp5_ASAP7_75t_L g1924 ( 
.A1(n_1902),
.A2(n_1790),
.B1(n_1884),
.B2(n_1870),
.Y(n_1924)
);

AO221x2_ASAP7_75t_L g1925 ( 
.A1(n_1903),
.A2(n_1872),
.B1(n_1846),
.B2(n_1857),
.C(n_1875),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1916),
.B(n_1881),
.Y(n_1926)
);

OAI221xp5_ASAP7_75t_L g1927 ( 
.A1(n_1912),
.A2(n_1781),
.B1(n_1785),
.B2(n_1819),
.C(n_1872),
.Y(n_1927)
);

OAI22xp33_ASAP7_75t_L g1928 ( 
.A1(n_1907),
.A2(n_1901),
.B1(n_1898),
.B2(n_1918),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1904),
.B(n_1886),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1897),
.B(n_1884),
.Y(n_1930)
);

OAI22xp33_ASAP7_75t_L g1931 ( 
.A1(n_1914),
.A2(n_1785),
.B1(n_1857),
.B2(n_1879),
.Y(n_1931)
);

CKINVDCx14_ASAP7_75t_R g1932 ( 
.A(n_1905),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1900),
.B(n_1893),
.Y(n_1933)
);

OAI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1911),
.A2(n_1876),
.B1(n_1869),
.B2(n_1892),
.Y(n_1934)
);

AOI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1913),
.A2(n_1811),
.B1(n_1781),
.B2(n_1693),
.Y(n_1935)
);

OR2x2_ASAP7_75t_L g1936 ( 
.A(n_1920),
.B(n_1882),
.Y(n_1936)
);

INVx2_ASAP7_75t_SL g1937 ( 
.A(n_1922),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1933),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1932),
.B(n_1874),
.Y(n_1939)
);

OAI32xp33_ASAP7_75t_L g1940 ( 
.A1(n_1927),
.A2(n_1908),
.A3(n_1910),
.B1(n_1899),
.B2(n_1882),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_SL g1941 ( 
.A(n_1931),
.B(n_1890),
.Y(n_1941)
);

NAND2x1_ASAP7_75t_L g1942 ( 
.A(n_1924),
.B(n_1930),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1923),
.B(n_1899),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1921),
.B(n_1926),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1919),
.B(n_1908),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1929),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1925),
.Y(n_1947)
);

INVx1_ASAP7_75t_SL g1948 ( 
.A(n_1935),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1925),
.Y(n_1949)
);

AOI32xp33_ASAP7_75t_L g1950 ( 
.A1(n_1934),
.A2(n_1910),
.A3(n_1819),
.B1(n_1836),
.B2(n_1768),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1928),
.Y(n_1951)
);

AOI21xp5_ASAP7_75t_L g1952 ( 
.A1(n_1941),
.A2(n_1811),
.B(n_1890),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1939),
.B(n_1816),
.Y(n_1953)
);

OAI21xp33_ASAP7_75t_L g1954 ( 
.A1(n_1950),
.A2(n_1792),
.B(n_1851),
.Y(n_1954)
);

OAI21xp5_ASAP7_75t_SL g1955 ( 
.A1(n_1948),
.A2(n_1728),
.B(n_1732),
.Y(n_1955)
);

NOR2xp33_ASAP7_75t_L g1956 ( 
.A(n_1947),
.B(n_1600),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1951),
.B(n_1858),
.Y(n_1957)
);

INVx1_ASAP7_75t_SL g1958 ( 
.A(n_1937),
.Y(n_1958)
);

OAI322xp33_ASAP7_75t_L g1959 ( 
.A1(n_1942),
.A2(n_1808),
.A3(n_1740),
.B1(n_1732),
.B2(n_1766),
.C1(n_1747),
.C2(n_1673),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1943),
.Y(n_1960)
);

OAI21xp5_ASAP7_75t_L g1961 ( 
.A1(n_1940),
.A2(n_1653),
.B(n_1719),
.Y(n_1961)
);

INVxp67_ASAP7_75t_L g1962 ( 
.A(n_1942),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1946),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1949),
.B(n_1706),
.Y(n_1964)
);

OAI211xp5_ASAP7_75t_L g1965 ( 
.A1(n_1962),
.A2(n_1945),
.B(n_1938),
.C(n_1944),
.Y(n_1965)
);

INVx2_ASAP7_75t_SL g1966 ( 
.A(n_1958),
.Y(n_1966)
);

INVx2_ASAP7_75t_SL g1967 ( 
.A(n_1953),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1960),
.B(n_1936),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1957),
.Y(n_1969)
);

AOI211xp5_ASAP7_75t_L g1970 ( 
.A1(n_1952),
.A2(n_1739),
.B(n_1725),
.C(n_1719),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1963),
.Y(n_1971)
);

OAI22x1_ASAP7_75t_L g1972 ( 
.A1(n_1956),
.A2(n_1803),
.B1(n_1619),
.B2(n_1743),
.Y(n_1972)
);

OAI22xp5_ASAP7_75t_L g1973 ( 
.A1(n_1955),
.A2(n_1961),
.B1(n_1964),
.B2(n_1954),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1959),
.B(n_1653),
.Y(n_1974)
);

OAI21xp33_ASAP7_75t_L g1975 ( 
.A1(n_1959),
.A2(n_1679),
.B(n_1799),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1958),
.B(n_1802),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1966),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1968),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1967),
.B(n_1779),
.Y(n_1979)
);

AOI322xp5_ASAP7_75t_L g1980 ( 
.A1(n_1974),
.A2(n_1730),
.A3(n_1814),
.B1(n_1809),
.B2(n_1807),
.C1(n_1815),
.C2(n_1812),
.Y(n_1980)
);

OAI31xp33_ASAP7_75t_L g1981 ( 
.A1(n_1965),
.A2(n_1724),
.A3(n_1658),
.B(n_1710),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1973),
.B(n_1813),
.Y(n_1982)
);

O2A1O1Ixp33_ASAP7_75t_SL g1983 ( 
.A1(n_1976),
.A2(n_1710),
.B(n_1713),
.C(n_1658),
.Y(n_1983)
);

AOI22xp5_ASAP7_75t_L g1984 ( 
.A1(n_1975),
.A2(n_1753),
.B1(n_1713),
.B2(n_1630),
.Y(n_1984)
);

AOI32xp33_ASAP7_75t_L g1985 ( 
.A1(n_1970),
.A2(n_1733),
.A3(n_1680),
.B1(n_1753),
.B2(n_1630),
.Y(n_1985)
);

AOI222xp33_ASAP7_75t_L g1986 ( 
.A1(n_1969),
.A2(n_1735),
.B1(n_1727),
.B2(n_351),
.C1(n_352),
.C2(n_353),
.Y(n_1986)
);

OAI22xp5_ASAP7_75t_L g1987 ( 
.A1(n_1971),
.A2(n_1735),
.B1(n_354),
.B2(n_349),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1977),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1979),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1978),
.Y(n_1990)
);

CKINVDCx20_ASAP7_75t_R g1991 ( 
.A(n_1982),
.Y(n_1991)
);

HB1xp67_ASAP7_75t_L g1992 ( 
.A(n_1987),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1984),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1983),
.Y(n_1994)
);

INVxp33_ASAP7_75t_SL g1995 ( 
.A(n_1986),
.Y(n_1995)
);

INVxp33_ASAP7_75t_SL g1996 ( 
.A(n_1985),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1980),
.B(n_1972),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1981),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1977),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1977),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1977),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1977),
.Y(n_2002)
);

NOR2xp33_ASAP7_75t_L g2003 ( 
.A(n_1977),
.B(n_1735),
.Y(n_2003)
);

INVx1_ASAP7_75t_SL g2004 ( 
.A(n_1977),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1988),
.Y(n_2005)
);

NOR2xp33_ASAP7_75t_L g2006 ( 
.A(n_1995),
.B(n_350),
.Y(n_2006)
);

AOI211x1_ASAP7_75t_L g2007 ( 
.A1(n_1998),
.A2(n_357),
.B(n_355),
.C(n_356),
.Y(n_2007)
);

NAND4xp75_ASAP7_75t_L g2008 ( 
.A(n_2000),
.B(n_360),
.C(n_358),
.D(n_359),
.Y(n_2008)
);

NOR2x1_ASAP7_75t_L g2009 ( 
.A(n_2004),
.B(n_361),
.Y(n_2009)
);

NOR3x1_ASAP7_75t_L g2010 ( 
.A(n_2001),
.B(n_362),
.C(n_365),
.Y(n_2010)
);

AOI221xp5_ASAP7_75t_L g2011 ( 
.A1(n_2004),
.A2(n_366),
.B1(n_367),
.B2(n_368),
.C(n_369),
.Y(n_2011)
);

NOR3xp33_ASAP7_75t_L g2012 ( 
.A(n_2002),
.B(n_371),
.C(n_372),
.Y(n_2012)
);

NOR3xp33_ASAP7_75t_L g2013 ( 
.A(n_1999),
.B(n_1993),
.C(n_1990),
.Y(n_2013)
);

INVxp67_ASAP7_75t_L g2014 ( 
.A(n_2003),
.Y(n_2014)
);

AOI22xp5_ASAP7_75t_L g2015 ( 
.A1(n_1996),
.A2(n_376),
.B1(n_373),
.B2(n_375),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_SL g2016 ( 
.A(n_1994),
.B(n_378),
.Y(n_2016)
);

AOI22xp5_ASAP7_75t_L g2017 ( 
.A1(n_1991),
.A2(n_383),
.B1(n_379),
.B2(n_380),
.Y(n_2017)
);

HB1xp67_ASAP7_75t_L g2018 ( 
.A(n_1992),
.Y(n_2018)
);

OAI221xp5_ASAP7_75t_L g2019 ( 
.A1(n_2013),
.A2(n_1989),
.B1(n_1997),
.B2(n_386),
.C(n_387),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_2018),
.Y(n_2020)
);

INVx1_ASAP7_75t_SL g2021 ( 
.A(n_2009),
.Y(n_2021)
);

AOI21xp33_ASAP7_75t_SL g2022 ( 
.A1(n_2005),
.A2(n_384),
.B(n_385),
.Y(n_2022)
);

AOI22xp5_ASAP7_75t_L g2023 ( 
.A1(n_2006),
.A2(n_395),
.B1(n_389),
.B2(n_392),
.Y(n_2023)
);

NAND4xp25_ASAP7_75t_L g2024 ( 
.A(n_2007),
.B(n_398),
.C(n_396),
.D(n_397),
.Y(n_2024)
);

NAND4xp25_ASAP7_75t_SL g2025 ( 
.A(n_2015),
.B(n_400),
.C(n_402),
.D(n_403),
.Y(n_2025)
);

OAI211xp5_ASAP7_75t_SL g2026 ( 
.A1(n_2014),
.A2(n_404),
.B(n_405),
.C(n_406),
.Y(n_2026)
);

INVx1_ASAP7_75t_SL g2027 ( 
.A(n_2016),
.Y(n_2027)
);

AOI322xp5_ASAP7_75t_L g2028 ( 
.A1(n_2012),
.A2(n_2011),
.A3(n_2010),
.B1(n_2017),
.B2(n_2008),
.C1(n_412),
.C2(n_413),
.Y(n_2028)
);

NAND4xp75_ASAP7_75t_L g2029 ( 
.A(n_2020),
.B(n_407),
.C(n_409),
.D(n_410),
.Y(n_2029)
);

AOI22xp5_ASAP7_75t_L g2030 ( 
.A1(n_2027),
.A2(n_411),
.B1(n_414),
.B2(n_415),
.Y(n_2030)
);

OAI211xp5_ASAP7_75t_L g2031 ( 
.A1(n_2019),
.A2(n_416),
.B(n_418),
.C(n_419),
.Y(n_2031)
);

OR5x1_ASAP7_75t_L g2032 ( 
.A(n_2024),
.B(n_2025),
.C(n_2026),
.D(n_2021),
.E(n_2028),
.Y(n_2032)
);

NAND3x1_ASAP7_75t_L g2033 ( 
.A(n_2023),
.B(n_420),
.C(n_421),
.Y(n_2033)
);

NAND4xp75_ASAP7_75t_L g2034 ( 
.A(n_2022),
.B(n_422),
.C(n_423),
.D(n_424),
.Y(n_2034)
);

NOR3xp33_ASAP7_75t_L g2035 ( 
.A(n_2019),
.B(n_425),
.C(n_426),
.Y(n_2035)
);

NOR2xp67_ASAP7_75t_L g2036 ( 
.A(n_2020),
.B(n_427),
.Y(n_2036)
);

NAND2x1p5_ASAP7_75t_L g2037 ( 
.A(n_2021),
.B(n_430),
.Y(n_2037)
);

NOR2x1_ASAP7_75t_L g2038 ( 
.A(n_2020),
.B(n_432),
.Y(n_2038)
);

OAI211xp5_ASAP7_75t_SL g2039 ( 
.A1(n_2019),
.A2(n_433),
.B(n_434),
.C(n_435),
.Y(n_2039)
);

NOR3xp33_ASAP7_75t_L g2040 ( 
.A(n_2019),
.B(n_436),
.C(n_437),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_2037),
.B(n_438),
.Y(n_2041)
);

AOI211xp5_ASAP7_75t_L g2042 ( 
.A1(n_2031),
.A2(n_440),
.B(n_441),
.C(n_442),
.Y(n_2042)
);

INVx2_ASAP7_75t_SL g2043 ( 
.A(n_2038),
.Y(n_2043)
);

NOR3xp33_ASAP7_75t_SL g2044 ( 
.A(n_2039),
.B(n_589),
.C(n_443),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_2036),
.Y(n_2045)
);

NOR4xp75_ASAP7_75t_L g2046 ( 
.A(n_2033),
.B(n_444),
.C(n_445),
.D(n_446),
.Y(n_2046)
);

AOI221xp5_ASAP7_75t_L g2047 ( 
.A1(n_2035),
.A2(n_447),
.B1(n_448),
.B2(n_449),
.C(n_450),
.Y(n_2047)
);

AOI211xp5_ASAP7_75t_L g2048 ( 
.A1(n_2040),
.A2(n_451),
.B(n_452),
.C(n_455),
.Y(n_2048)
);

AOI22xp5_ASAP7_75t_L g2049 ( 
.A1(n_2034),
.A2(n_456),
.B1(n_457),
.B2(n_458),
.Y(n_2049)
);

NAND3xp33_ASAP7_75t_SL g2050 ( 
.A(n_2030),
.B(n_459),
.C(n_460),
.Y(n_2050)
);

NAND3xp33_ASAP7_75t_L g2051 ( 
.A(n_2032),
.B(n_462),
.C(n_463),
.Y(n_2051)
);

AND2x4_ASAP7_75t_L g2052 ( 
.A(n_2029),
.B(n_464),
.Y(n_2052)
);

NOR4xp25_ASAP7_75t_L g2053 ( 
.A(n_2031),
.B(n_465),
.C(n_466),
.D(n_467),
.Y(n_2053)
);

NOR2x1p5_ASAP7_75t_L g2054 ( 
.A(n_2034),
.B(n_468),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2043),
.Y(n_2055)
);

AOI211xp5_ASAP7_75t_L g2056 ( 
.A1(n_2053),
.A2(n_469),
.B(n_473),
.C(n_474),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_2045),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_2052),
.B(n_475),
.Y(n_2058)
);

XNOR2xp5_ASAP7_75t_L g2059 ( 
.A(n_2046),
.B(n_476),
.Y(n_2059)
);

AOI21xp5_ASAP7_75t_L g2060 ( 
.A1(n_2051),
.A2(n_477),
.B(n_478),
.Y(n_2060)
);

INVx2_ASAP7_75t_SL g2061 ( 
.A(n_2041),
.Y(n_2061)
);

XNOR2xp5_ASAP7_75t_L g2062 ( 
.A(n_2054),
.B(n_479),
.Y(n_2062)
);

BUFx3_ASAP7_75t_L g2063 ( 
.A(n_2049),
.Y(n_2063)
);

AND2x4_ASAP7_75t_L g2064 ( 
.A(n_2044),
.B(n_480),
.Y(n_2064)
);

OR2x2_ASAP7_75t_L g2065 ( 
.A(n_2050),
.B(n_481),
.Y(n_2065)
);

AND2x4_ASAP7_75t_L g2066 ( 
.A(n_2042),
.B(n_483),
.Y(n_2066)
);

XNOR2xp5_ASAP7_75t_L g2067 ( 
.A(n_2048),
.B(n_484),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_2047),
.B(n_486),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_2041),
.B(n_487),
.Y(n_2069)
);

NOR2x1_ASAP7_75t_L g2070 ( 
.A(n_2051),
.B(n_588),
.Y(n_2070)
);

OR2x2_ASAP7_75t_L g2071 ( 
.A(n_2043),
.B(n_488),
.Y(n_2071)
);

NAND3x1_ASAP7_75t_L g2072 ( 
.A(n_2045),
.B(n_489),
.C(n_490),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_2055),
.B(n_2070),
.Y(n_2073)
);

NAND3x1_ASAP7_75t_L g2074 ( 
.A(n_2057),
.B(n_491),
.C(n_492),
.Y(n_2074)
);

OAI221xp5_ASAP7_75t_L g2075 ( 
.A1(n_2056),
.A2(n_493),
.B1(n_494),
.B2(n_501),
.C(n_503),
.Y(n_2075)
);

XOR2xp5_ASAP7_75t_L g2076 ( 
.A(n_2059),
.B(n_585),
.Y(n_2076)
);

OAI221xp5_ASAP7_75t_L g2077 ( 
.A1(n_2062),
.A2(n_505),
.B1(n_506),
.B2(n_507),
.C(n_509),
.Y(n_2077)
);

HB1xp67_ASAP7_75t_L g2078 ( 
.A(n_2072),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2061),
.B(n_2058),
.Y(n_2079)
);

XOR2xp5_ASAP7_75t_L g2080 ( 
.A(n_2067),
.B(n_510),
.Y(n_2080)
);

AO22x2_ASAP7_75t_L g2081 ( 
.A1(n_2071),
.A2(n_511),
.B1(n_512),
.B2(n_514),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_2064),
.B(n_516),
.Y(n_2082)
);

OAI221xp5_ASAP7_75t_L g2083 ( 
.A1(n_2060),
.A2(n_517),
.B1(n_518),
.B2(n_519),
.C(n_521),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_2066),
.B(n_522),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_2081),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2078),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2076),
.Y(n_2087)
);

AOI22xp5_ASAP7_75t_L g2088 ( 
.A1(n_2073),
.A2(n_2068),
.B1(n_2080),
.B2(n_2063),
.Y(n_2088)
);

AO22x2_ASAP7_75t_L g2089 ( 
.A1(n_2082),
.A2(n_2069),
.B1(n_2065),
.B2(n_525),
.Y(n_2089)
);

AOI31xp33_ASAP7_75t_L g2090 ( 
.A1(n_2079),
.A2(n_584),
.A3(n_524),
.B(n_528),
.Y(n_2090)
);

HB1xp67_ASAP7_75t_L g2091 ( 
.A(n_2074),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_2081),
.Y(n_2092)
);

AOI22xp5_ASAP7_75t_L g2093 ( 
.A1(n_2075),
.A2(n_523),
.B1(n_529),
.B2(n_531),
.Y(n_2093)
);

AOI21xp5_ASAP7_75t_L g2094 ( 
.A1(n_2086),
.A2(n_2084),
.B(n_2083),
.Y(n_2094)
);

XNOR2xp5_ASAP7_75t_L g2095 ( 
.A(n_2088),
.B(n_2077),
.Y(n_2095)
);

AOI211x1_ASAP7_75t_L g2096 ( 
.A1(n_2087),
.A2(n_533),
.B(n_535),
.C(n_537),
.Y(n_2096)
);

XNOR2xp5_ASAP7_75t_L g2097 ( 
.A(n_2089),
.B(n_538),
.Y(n_2097)
);

OAI22xp33_ASAP7_75t_L g2098 ( 
.A1(n_2094),
.A2(n_2092),
.B1(n_2085),
.B2(n_2091),
.Y(n_2098)
);

OA21x2_ASAP7_75t_L g2099 ( 
.A1(n_2095),
.A2(n_2093),
.B(n_2090),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2099),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_2098),
.Y(n_2101)
);

AOI21xp33_ASAP7_75t_SL g2102 ( 
.A1(n_2101),
.A2(n_2097),
.B(n_2096),
.Y(n_2102)
);

AOI222xp33_ASAP7_75t_L g2103 ( 
.A1(n_2100),
.A2(n_539),
.B1(n_540),
.B2(n_541),
.C1(n_542),
.C2(n_544),
.Y(n_2103)
);

OAI22xp5_ASAP7_75t_L g2104 ( 
.A1(n_2102),
.A2(n_546),
.B1(n_547),
.B2(n_551),
.Y(n_2104)
);

AOI22xp5_ASAP7_75t_L g2105 ( 
.A1(n_2103),
.A2(n_552),
.B1(n_553),
.B2(n_556),
.Y(n_2105)
);

AOI21xp33_ASAP7_75t_SL g2106 ( 
.A1(n_2104),
.A2(n_558),
.B(n_559),
.Y(n_2106)
);

NOR2xp33_ASAP7_75t_L g2107 ( 
.A(n_2105),
.B(n_561),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2107),
.Y(n_2108)
);

OR2x2_ASAP7_75t_L g2109 ( 
.A(n_2106),
.B(n_582),
.Y(n_2109)
);

AOI22xp5_ASAP7_75t_L g2110 ( 
.A1(n_2108),
.A2(n_563),
.B1(n_564),
.B2(n_565),
.Y(n_2110)
);

AOI211xp5_ASAP7_75t_L g2111 ( 
.A1(n_2110),
.A2(n_2109),
.B(n_566),
.C(n_567),
.Y(n_2111)
);


endmodule