module fake_jpeg_11613_n_146 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_146);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

AND2x2_ASAP7_75t_SL g34 ( 
.A(n_27),
.B(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_34),
.B(n_35),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_3),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_3),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_36),
.B(n_39),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_37),
.B(n_47),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_12),
.B(n_4),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_4),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_12),
.B(n_28),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_52),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_23),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_11),
.B(n_21),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_54),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_55),
.A2(n_56),
.B1(n_16),
.B2(n_18),
.Y(n_57)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

AO22x2_ASAP7_75t_L g60 ( 
.A1(n_34),
.A2(n_18),
.B1(n_20),
.B2(n_6),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_60),
.A2(n_79),
.B1(n_82),
.B2(n_77),
.Y(n_100)
);

NOR2x1_ASAP7_75t_L g69 ( 
.A(n_35),
.B(n_20),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_68),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_33),
.A2(n_22),
.B1(n_26),
.B2(n_21),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_72),
.A2(n_74),
.B1(n_75),
.B2(n_77),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_36),
.A2(n_39),
.B1(n_54),
.B2(n_50),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_59),
.B1(n_60),
.B2(n_75),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_22),
.B1(n_26),
.B2(n_23),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_28),
.B1(n_6),
.B2(n_5),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_44),
.A2(n_5),
.B1(n_7),
.B2(n_41),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_51),
.A2(n_34),
.B1(n_38),
.B2(n_54),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_44),
.A2(n_19),
.B1(n_29),
.B2(n_33),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_82),
.A2(n_43),
.B1(n_51),
.B2(n_57),
.Y(n_86)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_SL g112 ( 
.A1(n_86),
.A2(n_65),
.B(n_76),
.C(n_80),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_69),
.B(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_87),
.B(n_90),
.Y(n_103)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_70),
.B(n_68),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_92),
.B(n_94),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_78),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_67),
.B1(n_58),
.B2(n_78),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_97),
.Y(n_111)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_62),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_98),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_72),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_100),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_60),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_100),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_108),
.A2(n_112),
.B1(n_88),
.B2(n_93),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_58),
.C(n_76),
.Y(n_110)
);

FAx1_ASAP7_75t_SL g113 ( 
.A(n_110),
.B(n_91),
.CI(n_86),
.CON(n_113),
.SN(n_113)
);

AOI21x1_ASAP7_75t_L g126 ( 
.A1(n_113),
.A2(n_112),
.B(n_106),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_121),
.B(n_112),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_104),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_117),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_116),
.B(n_119),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_110),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_95),
.B1(n_88),
.B2(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_100),
.B1(n_67),
.B2(n_80),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_102),
.A2(n_65),
.B1(n_96),
.B2(n_108),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_122),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_65),
.B(n_111),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_105),
.B(n_103),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_109),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_127),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_129),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_130),
.A2(n_120),
.B1(n_115),
.B2(n_122),
.Y(n_137)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_127),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_132),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_125),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_134),
.B(n_117),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_133),
.A2(n_128),
.B1(n_123),
.B2(n_114),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_119),
.C(n_118),
.Y(n_141)
);

OAI21x1_ASAP7_75t_SL g139 ( 
.A1(n_136),
.A2(n_137),
.B(n_133),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_140),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_138),
.A2(n_130),
.B(n_134),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_141),
.B(n_135),
.Y(n_143)
);

OAI21x1_ASAP7_75t_SL g144 ( 
.A1(n_143),
.A2(n_136),
.B(n_113),
.Y(n_144)
);

OAI21x1_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_142),
.B(n_124),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_124),
.C(n_112),
.Y(n_146)
);


endmodule