module real_jpeg_20507_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx13_ASAP7_75t_L g88 ( 
.A(n_0),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_1),
.A2(n_37),
.B1(n_75),
.B2(n_76),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_1),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_2),
.A2(n_72),
.B1(n_78),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_2),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_2),
.A2(n_75),
.B1(n_76),
.B2(n_81),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_81),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_2),
.A2(n_40),
.B1(n_41),
.B2(n_81),
.Y(n_194)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_3),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_L g152 ( 
.A1(n_3),
.A2(n_14),
.B(n_30),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_3),
.A2(n_40),
.B1(n_41),
.B2(n_102),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_3),
.A2(n_60),
.B1(n_64),
.B2(n_161),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_3),
.B(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_3),
.B(n_76),
.Y(n_186)
);

AOI21xp33_ASAP7_75t_L g190 ( 
.A1(n_3),
.A2(n_76),
.B(n_186),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_3),
.B(n_74),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_4),
.A2(n_31),
.B1(n_40),
.B2(n_41),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_4),
.A2(n_31),
.B1(n_75),
.B2(n_76),
.Y(n_95)
);

BUFx16f_ASAP7_75t_L g72 ( 
.A(n_5),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_6),
.A2(n_72),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_6),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_6),
.A2(n_75),
.B1(n_76),
.B2(n_79),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_79),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_6),
.A2(n_40),
.B1(n_41),
.B2(n_79),
.Y(n_177)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_9),
.A2(n_72),
.B1(n_78),
.B2(n_114),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_9),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_9),
.A2(n_40),
.B1(n_41),
.B2(n_114),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_114),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_9),
.A2(n_75),
.B1(n_76),
.B2(n_114),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_11),
.A2(n_40),
.B1(n_41),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_11),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_49),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_12),
.A2(n_40),
.B1(n_41),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_12),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_47),
.Y(n_104)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_13),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_13),
.A2(n_71),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_14),
.A2(n_40),
.B(n_43),
.C(n_44),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_14),
.B(n_40),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_45),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_15),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_134),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_133),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_116),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_20),
.B(n_116),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_97),
.B2(n_115),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_50),
.B2(n_51),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_38),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_35),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_26),
.A2(n_64),
.B(n_104),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_32),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_28),
.B(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_29),
.B(n_165),
.Y(n_164)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_32),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_32),
.A2(n_36),
.B(n_63),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_34),
.A2(n_60),
.B1(n_145),
.B2(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_35),
.A2(n_60),
.B(n_148),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_44),
.B1(n_46),
.B2(n_48),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_39),
.A2(n_125),
.B(n_127),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_39),
.A2(n_44),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_39),
.A2(n_44),
.B1(n_156),
.B2(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_39),
.A2(n_44),
.B1(n_177),
.B2(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_39),
.A2(n_194),
.B(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_40),
.A2(n_41),
.B1(n_87),
.B2(n_91),
.Y(n_90)
);

AOI32xp33_ASAP7_75t_L g185 ( 
.A1(n_40),
.A2(n_75),
.A3(n_91),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_41),
.A2(n_45),
.B(n_102),
.C(n_152),
.Y(n_151)
);

NAND2xp33_ASAP7_75t_SL g187 ( 
.A(n_41),
.B(n_87),
.Y(n_187)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_46),
.B(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_44),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_44),
.B(n_102),
.Y(n_159)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_65),
.B1(n_66),
.B2(n_96),
.Y(n_51)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_58),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_53),
.A2(n_54),
.B1(n_58),
.B2(n_59),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_56),
.B(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B(n_62),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_60),
.A2(n_61),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_64),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_64),
.B(n_102),
.Y(n_165)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_83),
.B2(n_84),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_77),
.B1(n_80),
.B2(n_82),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_69),
.A2(n_77),
.B1(n_82),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_70),
.A2(n_74),
.B1(n_101),
.B2(n_113),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B(n_73),
.C(n_74),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_72),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_76),
.Y(n_100)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

HAxp5_ASAP7_75t_SL g101 ( 
.A(n_72),
.B(n_102),
.CON(n_101),
.SN(n_101)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_73),
.A2(n_75),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_74),
.Y(n_82)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_87),
.B(n_89),
.C(n_90),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_87),
.Y(n_89)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_92),
.B(n_94),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_85),
.A2(n_107),
.B(n_109),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_85),
.A2(n_174),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_86),
.A2(n_90),
.B1(n_108),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_86),
.A2(n_90),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_93),
.Y(n_109)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_90),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_97),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_106),
.C(n_110),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_99),
.B(n_103),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_106),
.A2(n_110),
.B1(n_111),
.B2(n_120),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_106),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.C(n_122),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_117),
.A2(n_118),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_121),
.B(n_122),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_129),
.C(n_132),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_123),
.A2(n_124),
.B1(n_129),
.B2(n_130),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_126),
.B(n_128),
.Y(n_216)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_131),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_132),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_234),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_229),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_218),
.B(n_228),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_199),
.B(n_217),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_180),
.B(n_198),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_168),
.B(n_179),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_157),
.B(n_167),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_149),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_149),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_153),
.B2(n_154),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_151),
.B(n_153),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_162),
.B(n_166),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_160),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_169),
.B(n_170),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_178),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_176),
.C(n_178),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_182),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_188),
.B1(n_196),
.B2(n_197),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_183),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_185),
.Y(n_214)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_192),
.B1(n_193),
.B2(n_195),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_189),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_191),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_195),
.C(n_196),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_200),
.B(n_201),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_212),
.B2(n_213),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_214),
.C(n_215),
.Y(n_219)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_209),
.C(n_210),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_219),
.B(n_220),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_226),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_225),
.C(n_226),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_224),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_231),
.Y(n_235)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);


endmodule