module fake_jpeg_3013_n_526 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_526);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_526;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_5),
.B(n_9),
.Y(n_25)
);

BUFx4f_ASAP7_75t_SL g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_53),
.Y(n_136)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_54),
.Y(n_142)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_56),
.Y(n_122)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_57),
.Y(n_137)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_63),
.Y(n_153)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_65),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_66),
.B(n_71),
.Y(n_115)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_67),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_68),
.Y(n_161)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_47),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_73),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_74),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_34),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_75),
.A2(n_25),
.B1(n_45),
.B2(n_44),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_15),
.Y(n_76)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_81),
.Y(n_163)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_16),
.Y(n_84)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_16),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_16),
.Y(n_86)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_25),
.B(n_14),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_87),
.B(n_41),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_88),
.Y(n_156)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_16),
.Y(n_89)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_90),
.Y(n_164)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_94),
.Y(n_166)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_95),
.Y(n_167)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_97),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

NAND2xp33_ASAP7_75t_SL g116 ( 
.A(n_99),
.B(n_101),
.Y(n_116)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_21),
.Y(n_100)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_21),
.Y(n_103)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_103),
.Y(n_158)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_26),
.Y(n_104)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_105),
.Y(n_169)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_26),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_106),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_38),
.Y(n_107)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_107),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_128),
.A2(n_132),
.B1(n_162),
.B2(n_22),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_87),
.A2(n_38),
.B1(n_28),
.B2(n_17),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_103),
.B(n_17),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_139),
.B(n_141),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_56),
.B(n_28),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_143),
.B(n_151),
.Y(n_209)
);

AOI21xp33_ASAP7_75t_SL g144 ( 
.A1(n_57),
.A2(n_41),
.B(n_20),
.Y(n_144)
);

AND2x2_ASAP7_75t_SL g215 ( 
.A(n_144),
.B(n_107),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_98),
.B(n_50),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_146),
.B(n_149),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_53),
.B(n_50),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_93),
.A2(n_26),
.B1(n_44),
.B2(n_24),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_150),
.A2(n_159),
.B1(n_92),
.B2(n_73),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_56),
.B(n_24),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_59),
.A2(n_22),
.B1(n_38),
.B2(n_33),
.Y(n_157)
);

OAI22x1_ASAP7_75t_L g195 ( 
.A1(n_157),
.A2(n_59),
.B1(n_76),
.B2(n_106),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_63),
.A2(n_22),
.B1(n_33),
.B2(n_32),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_94),
.A2(n_38),
.B1(n_32),
.B2(n_45),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_115),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_173),
.B(n_175),
.Y(n_255)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_109),
.Y(n_174)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_174),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_177),
.Y(n_248)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_178),
.Y(n_250)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_170),
.Y(n_179)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_179),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_163),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_180),
.Y(n_258)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_120),
.Y(n_181)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_181),
.Y(n_254)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_154),
.Y(n_182)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_182),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_183),
.Y(n_244)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_184),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_185),
.Y(n_235)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_186),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_163),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_187),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_137),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_188),
.A2(n_195),
.B1(n_197),
.B2(n_207),
.Y(n_253)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_137),
.Y(n_189)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_189),
.Y(n_229)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_138),
.Y(n_190)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_190),
.Y(n_228)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_112),
.Y(n_191)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_191),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_122),
.Y(n_192)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_192),
.Y(n_230)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_122),
.Y(n_194)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_194),
.Y(n_251)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_155),
.Y(n_196)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_196),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_159),
.A2(n_75),
.B1(n_65),
.B2(n_68),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_198),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_243)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_113),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_199),
.B(n_211),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_152),
.Y(n_200)
);

BUFx4f_ASAP7_75t_SL g201 ( 
.A(n_145),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_118),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_117),
.B(n_37),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_210),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_125),
.A2(n_88),
.B1(n_74),
.B2(n_80),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_208),
.Y(n_259)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_124),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_126),
.Y(n_206)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_134),
.Y(n_208)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_110),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_172),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_119),
.B(n_20),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_213),
.Y(n_231)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_129),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_111),
.B(n_76),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_217),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_215),
.A2(n_218),
.B(n_157),
.Y(n_232)
);

INVx3_ASAP7_75t_SL g216 ( 
.A(n_108),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_216),
.A2(n_171),
.B1(n_136),
.B2(n_161),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_145),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_121),
.A2(n_37),
.B1(n_90),
.B2(n_83),
.Y(n_218)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_171),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_153),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_148),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_220),
.B(n_221),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_148),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_222),
.A2(n_136),
.B1(n_161),
.B2(n_160),
.Y(n_241)
);

OAI21xp33_ASAP7_75t_SL g288 ( 
.A1(n_232),
.A2(n_202),
.B(n_208),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_131),
.C(n_167),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_236),
.B(n_213),
.C(n_199),
.Y(n_271)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_237),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_193),
.B(n_168),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_247),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_241),
.A2(n_216),
.B1(n_181),
.B2(n_179),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_222),
.A2(n_135),
.B1(n_140),
.B2(n_160),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_245),
.A2(n_249),
.B1(n_216),
.B2(n_156),
.Y(n_269)
);

O2A1O1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_215),
.A2(n_116),
.B(n_145),
.C(n_127),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_246),
.A2(n_123),
.B(n_127),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_193),
.B(n_168),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_203),
.A2(n_142),
.B1(n_153),
.B2(n_97),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_176),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_261),
.B(n_267),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_226),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_263),
.B(n_274),
.Y(n_308)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_234),
.Y(n_265)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_265),
.Y(n_296)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_266),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_212),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_231),
.A2(n_195),
.B1(n_187),
.B2(n_180),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_268),
.A2(n_283),
.B1(n_253),
.B2(n_276),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_269),
.B(n_276),
.Y(n_298)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_270),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_271),
.B(n_250),
.C(n_225),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_186),
.Y(n_272)
);

AND2x2_ASAP7_75t_SL g310 ( 
.A(n_272),
.B(n_284),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_209),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_273),
.B(n_278),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_226),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_248),
.Y(n_275)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_275),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_225),
.Y(n_277)
);

NAND2xp33_ASAP7_75t_SL g301 ( 
.A(n_277),
.B(n_279),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_227),
.B(n_173),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_247),
.B(n_174),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_281),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_227),
.B(n_257),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_190),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_282),
.B(n_285),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_241),
.A2(n_142),
.B1(n_177),
.B2(n_178),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_256),
.B(n_182),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_196),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_232),
.A2(n_191),
.B1(n_123),
.B2(n_210),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_286),
.A2(n_290),
.B1(n_269),
.B2(n_189),
.Y(n_294)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_230),
.Y(n_287)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_287),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_288),
.A2(n_289),
.B(n_258),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_206),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_246),
.A2(n_205),
.B1(n_192),
.B2(n_194),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_265),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_291),
.B(n_305),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_279),
.A2(n_246),
.B(n_258),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_292),
.A2(n_294),
.B(n_300),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_284),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_293),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_288),
.A2(n_236),
.B1(n_253),
.B2(n_239),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_304),
.A2(n_309),
.B1(n_318),
.B2(n_277),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_284),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_306),
.A2(n_316),
.B1(n_272),
.B2(n_268),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_282),
.A2(n_238),
.B(n_254),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_307),
.A2(n_289),
.B(n_284),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_264),
.A2(n_254),
.B1(n_252),
.B2(n_250),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_271),
.B(n_238),
.C(n_252),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_311),
.B(n_313),
.C(n_270),
.Y(n_339)
);

OAI32xp33_ASAP7_75t_L g315 ( 
.A1(n_260),
.A2(n_198),
.A3(n_223),
.B1(n_200),
.B2(n_259),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_315),
.B(n_290),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_260),
.A2(n_228),
.B1(n_108),
.B2(n_114),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_264),
.A2(n_228),
.B1(n_233),
.B2(n_242),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_266),
.Y(n_319)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_319),
.Y(n_335)
);

NAND2xp67_ASAP7_75t_L g320 ( 
.A(n_292),
.B(n_274),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_320),
.A2(n_342),
.B1(n_346),
.B2(n_322),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_302),
.B(n_261),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_321),
.B(n_312),
.Y(n_364)
);

INVx3_ASAP7_75t_SL g322 ( 
.A(n_298),
.Y(n_322)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_322),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_323),
.A2(n_331),
.B1(n_338),
.B2(n_343),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_313),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_324),
.B(n_330),
.C(n_334),
.Y(n_353)
);

INVxp33_ASAP7_75t_L g326 ( 
.A(n_307),
.Y(n_326)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_326),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_311),
.B(n_273),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_327),
.B(n_333),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_309),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_328),
.B(n_332),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_302),
.B(n_271),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_306),
.A2(n_304),
.B1(n_300),
.B2(n_298),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_318),
.Y(n_332)
);

XOR2x2_ASAP7_75t_L g333 ( 
.A(n_303),
.B(n_281),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_303),
.B(n_278),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_303),
.B(n_267),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_336),
.B(n_339),
.C(n_340),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_298),
.A2(n_280),
.B1(n_263),
.B2(n_268),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_314),
.B(n_285),
.C(n_275),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_299),
.B(n_314),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_341),
.B(n_310),
.C(n_317),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_298),
.A2(n_272),
.B1(n_262),
.B2(n_283),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_344),
.Y(n_365)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_291),
.Y(n_345)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_345),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_299),
.A2(n_286),
.B1(n_272),
.B2(n_262),
.Y(n_347)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_347),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_308),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_348),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_324),
.B(n_314),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_350),
.B(n_356),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_328),
.A2(n_308),
.B1(n_305),
.B2(n_293),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_351),
.A2(n_361),
.B1(n_362),
.B2(n_363),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_341),
.B(n_315),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g399 ( 
.A(n_359),
.B(n_371),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_339),
.B(n_310),
.C(n_317),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_360),
.B(n_372),
.C(n_376),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_342),
.A2(n_316),
.B1(n_294),
.B2(n_291),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_338),
.A2(n_291),
.B1(n_301),
.B2(n_319),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_364),
.A2(n_366),
.B1(n_367),
.B2(n_375),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_322),
.A2(n_301),
.B1(n_312),
.B2(n_297),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_331),
.A2(n_297),
.B1(n_296),
.B2(n_310),
.Y(n_367)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_335),
.Y(n_369)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_369),
.Y(n_379)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_335),
.Y(n_370)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_370),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_330),
.B(n_296),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_327),
.B(n_310),
.C(n_235),
.Y(n_372)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_325),
.Y(n_374)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_374),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_348),
.A2(n_295),
.B1(n_277),
.B2(n_287),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_336),
.B(n_235),
.C(n_251),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_325),
.Y(n_377)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_377),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_378),
.B(n_329),
.Y(n_380)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_380),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_360),
.B(n_334),
.Y(n_383)
);

CKINVDCx14_ASAP7_75t_R g410 ( 
.A(n_383),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_358),
.A2(n_323),
.B1(n_344),
.B2(n_343),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_385),
.A2(n_394),
.B1(n_404),
.B2(n_361),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_354),
.B(n_345),
.Y(n_386)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_386),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_355),
.B(n_340),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_387),
.Y(n_430)
);

OA21x2_ASAP7_75t_L g388 ( 
.A1(n_349),
.A2(n_337),
.B(n_320),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_388),
.B(n_407),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_365),
.A2(n_337),
.B(n_333),
.Y(n_389)
);

AO21x1_ASAP7_75t_L g414 ( 
.A1(n_389),
.A2(n_396),
.B(n_402),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_355),
.B(n_295),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_391),
.B(n_405),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_353),
.B(n_251),
.C(n_229),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_392),
.B(n_393),
.C(n_356),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_353),
.B(n_224),
.C(n_229),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_349),
.A2(n_287),
.B1(n_233),
.B2(n_230),
.Y(n_394)
);

A2O1A1Ixp33_ASAP7_75t_SL g396 ( 
.A1(n_363),
.A2(n_243),
.B(n_201),
.C(n_224),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_373),
.B(n_223),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_400),
.B(n_406),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_376),
.B(n_352),
.Y(n_401)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_401),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_351),
.A2(n_242),
.B(n_244),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_375),
.B(n_219),
.Y(n_403)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_403),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_357),
.A2(n_201),
.B1(n_244),
.B2(n_183),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_350),
.B(n_175),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_373),
.B(n_105),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_367),
.A2(n_184),
.B(n_14),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_409),
.B(n_419),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_380),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_413),
.B(n_418),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_382),
.B(n_371),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_416),
.B(n_427),
.Y(n_432)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_386),
.Y(n_417)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_417),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_393),
.B(n_372),
.C(n_359),
.Y(n_418)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_379),
.Y(n_420)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_420),
.Y(n_447)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_381),
.Y(n_421)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_421),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_384),
.B(n_362),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g442 ( 
.A(n_422),
.B(n_426),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_392),
.B(n_366),
.C(n_368),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_424),
.B(n_396),
.Y(n_446)
);

MAJx2_ASAP7_75t_L g425 ( 
.A(n_399),
.B(n_368),
.C(n_30),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_425),
.B(n_407),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_395),
.B(n_164),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_382),
.B(n_164),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_397),
.A2(n_156),
.B1(n_114),
.B2(n_54),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_428),
.A2(n_394),
.B1(n_404),
.B2(n_403),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_409),
.B(n_390),
.C(n_400),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_433),
.B(n_434),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_427),
.B(n_390),
.C(n_406),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_418),
.B(n_385),
.C(n_389),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_435),
.B(n_438),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_424),
.B(n_402),
.C(n_398),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_416),
.B(n_408),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_439),
.B(n_443),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_410),
.B(n_388),
.C(n_399),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_440),
.B(n_450),
.C(n_451),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_441),
.A2(n_39),
.B1(n_31),
.B2(n_43),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_431),
.B(n_388),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_449),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_446),
.B(n_419),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_430),
.A2(n_396),
.B(n_10),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_448),
.A2(n_414),
.B(n_421),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_429),
.B(n_396),
.C(n_39),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_408),
.B(n_39),
.C(n_31),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_417),
.B(n_31),
.C(n_39),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_445),
.A2(n_412),
.B1(n_411),
.B2(n_423),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_453),
.A2(n_468),
.B1(n_469),
.B2(n_471),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_454),
.B(n_457),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_442),
.A2(n_412),
.B(n_414),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_455),
.A2(n_459),
.B(n_2),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_433),
.B(n_436),
.C(n_438),
.Y(n_457)
);

AO21x1_ASAP7_75t_L g458 ( 
.A1(n_442),
.A2(n_422),
.B(n_415),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g478 ( 
.A(n_458),
.B(n_453),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_437),
.A2(n_415),
.B(n_428),
.Y(n_459)
);

XNOR2x1_ASAP7_75t_L g485 ( 
.A(n_464),
.B(n_2),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_436),
.B(n_439),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_465),
.B(n_467),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_434),
.B(n_425),
.C(n_426),
.Y(n_466)
);

NOR2xp67_ASAP7_75t_SL g486 ( 
.A(n_466),
.B(n_18),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_440),
.B(n_432),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_447),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_452),
.A2(n_420),
.B1(n_443),
.B2(n_435),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_43),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_470),
.B(n_1),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_462),
.B(n_39),
.C(n_31),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_472),
.B(n_473),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_457),
.B(n_31),
.C(n_30),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_467),
.B(n_18),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_474),
.B(n_477),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_455),
.A2(n_13),
.B1(n_11),
.B2(n_10),
.Y(n_476)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_476),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_464),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_478),
.B(n_479),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_463),
.B(n_13),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_458),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_480),
.B(n_482),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_465),
.B(n_18),
.C(n_15),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_483),
.B(n_485),
.Y(n_499)
);

AOI21x1_ASAP7_75t_L g496 ( 
.A1(n_484),
.A2(n_2),
.B(n_3),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_486),
.B(n_461),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_477),
.B(n_466),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_489),
.B(n_490),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_475),
.B(n_460),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_481),
.B(n_456),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_491),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_481),
.B(n_456),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_494),
.A2(n_495),
.B1(n_498),
.B2(n_500),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_478),
.B(n_487),
.Y(n_495)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_496),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_483),
.A2(n_471),
.B1(n_461),
.B2(n_470),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_497),
.A2(n_485),
.B(n_482),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_502),
.A2(n_509),
.B(n_4),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_492),
.B(n_18),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_505),
.B(n_508),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_493),
.B(n_501),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_499),
.B(n_9),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_498),
.B(n_488),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_510),
.B(n_511),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_499),
.B(n_3),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_507),
.B(n_496),
.Y(n_512)
);

NAND3xp33_ASAP7_75t_L g519 ( 
.A(n_512),
.B(n_513),
.C(n_516),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_503),
.B(n_510),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_504),
.B(n_3),
.C(n_4),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_515),
.A2(n_506),
.B(n_511),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_518),
.A2(n_520),
.B(n_521),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_517),
.B(n_505),
.C(n_5),
.Y(n_520)
);

NAND2xp33_ASAP7_75t_L g521 ( 
.A(n_517),
.B(n_4),
.Y(n_521)
);

OAI321xp33_ASAP7_75t_L g523 ( 
.A1(n_519),
.A2(n_514),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_523)
);

AOI31xp33_ASAP7_75t_L g524 ( 
.A1(n_523),
.A2(n_5),
.A3(n_6),
.B(n_8),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_522),
.C(n_6),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_8),
.C(n_380),
.Y(n_526)
);


endmodule