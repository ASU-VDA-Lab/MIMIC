module real_aes_257_n_7 (n_4, n_0, n_3, n_5, n_2, n_6, n_1, n_7);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_6;
input n_1;
output n_7;
wire n_16;
wire n_17;
wire n_13;
wire n_18;
wire n_15;
wire n_8;
wire n_9;
wire n_12;
wire n_14;
wire n_10;
wire n_11;
OAI22xp5_ASAP7_75t_L g14 ( .A1(n_0), .A2(n_4), .B1(n_15), .B2(n_16), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_0), .Y(n_16) );
CKINVDCx16_ASAP7_75t_R g18 ( .A(n_1), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_2), .B(n_18), .Y(n_17) );
BUFx2_ASAP7_75t_SL g10 ( .A(n_3), .Y(n_10) );
INVx1_ASAP7_75t_L g15 ( .A(n_4), .Y(n_15) );
AOI221xp5_ASAP7_75t_L g7 ( .A1(n_5), .A2(n_8), .B1(n_13), .B2(n_14), .C(n_17), .Y(n_7) );
CKINVDCx16_ASAP7_75t_R g12 ( .A(n_6), .Y(n_12) );
INVx1_ASAP7_75t_SL g13 ( .A(n_8), .Y(n_13) );
NOR2xp33_ASAP7_75t_SL g8 ( .A(n_9), .B(n_11), .Y(n_8) );
CKINVDCx8_ASAP7_75t_R g9 ( .A(n_10), .Y(n_9) );
CKINVDCx16_ASAP7_75t_R g11 ( .A(n_12), .Y(n_11) );
endmodule