module fake_jpeg_30130_n_483 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_483);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_483;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_SL g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_16),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_49),
.B(n_82),
.Y(n_101)
);

BUFx12f_ASAP7_75t_SL g50 ( 
.A(n_39),
.Y(n_50)
);

NAND2x1_ASAP7_75t_SL g120 ( 
.A(n_50),
.B(n_19),
.Y(n_120)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_55),
.Y(n_135)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_56),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_46),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_58),
.B(n_59),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_16),
.Y(n_59)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx4f_ASAP7_75t_SL g150 ( 
.A(n_60),
.Y(n_150)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_62),
.B(n_70),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_64),
.Y(n_115)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx11_ASAP7_75t_L g136 ( 
.A(n_65),
.Y(n_136)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_69),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_15),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx5_ASAP7_75t_SL g112 ( 
.A(n_72),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_15),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_77),
.Y(n_119)
);

BUFx16f_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

BUFx16f_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_75),
.Y(n_153)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_46),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g154 ( 
.A(n_78),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_20),
.B(n_15),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_81),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_17),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_46),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_20),
.B(n_25),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_85),
.B(n_89),
.Y(n_130)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_23),
.B(n_14),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_88),
.B(n_32),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_23),
.B(n_14),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_46),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_97),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_25),
.B(n_34),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_74),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_102),
.B(n_133),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_50),
.A2(n_47),
.B1(n_29),
.B2(n_28),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_117),
.A2(n_121),
.B1(n_72),
.B2(n_54),
.Y(n_203)
);

NAND2xp33_ASAP7_75t_SL g159 ( 
.A(n_120),
.B(n_96),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_59),
.A2(n_86),
.B1(n_95),
.B2(n_57),
.Y(n_121)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_63),
.A2(n_24),
.B1(n_43),
.B2(n_29),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_129),
.A2(n_92),
.B1(n_91),
.B2(n_87),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_66),
.A2(n_34),
.B1(n_45),
.B2(n_26),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_132),
.B(n_149),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_74),
.Y(n_133)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_75),
.B(n_40),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_141),
.B(n_155),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_60),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_152),
.Y(n_158)
);

CKINVDCx12_ASAP7_75t_R g144 ( 
.A(n_60),
.Y(n_144)
);

CKINVDCx12_ASAP7_75t_R g187 ( 
.A(n_144),
.Y(n_187)
);

AOI21xp33_ASAP7_75t_L g149 ( 
.A1(n_78),
.A2(n_32),
.B(n_45),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_78),
.B(n_40),
.Y(n_152)
);

BUFx4f_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

INVx3_ASAP7_75t_SL g215 ( 
.A(n_156),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_116),
.A2(n_93),
.B1(n_83),
.B2(n_98),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_157),
.A2(n_112),
.B1(n_114),
.B2(n_145),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_159),
.B(n_169),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_106),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_161),
.B(n_168),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_104),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_162),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_104),
.Y(n_164)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_164),
.Y(n_246)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_165),
.Y(n_218)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_166),
.Y(n_211)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_118),
.Y(n_167)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_167),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_134),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_114),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_108),
.Y(n_171)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_171),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_106),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_172),
.B(n_179),
.Y(n_238)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_173),
.Y(n_236)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_99),
.Y(n_174)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_174),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_175),
.Y(n_239)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_176),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_177),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_178),
.A2(n_183),
.B1(n_192),
.B2(n_208),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_110),
.B(n_119),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_107),
.Y(n_181)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_182),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_126),
.A2(n_80),
.B1(n_137),
.B2(n_116),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_125),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_184),
.B(n_189),
.Y(n_249)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_118),
.Y(n_185)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_185),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_123),
.Y(n_186)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_146),
.Y(n_188)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_188),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_120),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_123),
.Y(n_190)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_130),
.B(n_105),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_191),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_126),
.A2(n_47),
.B1(n_29),
.B2(n_68),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_101),
.B(n_85),
.Y(n_193)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_193),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_128),
.B(n_85),
.Y(n_194)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_194),
.Y(n_248)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_109),
.Y(n_197)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_197),
.Y(n_243)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_100),
.Y(n_198)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_198),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_103),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_115),
.B(n_26),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_43),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_109),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_202),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_65),
.Y(n_240)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_140),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_204),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_122),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_205),
.A2(n_206),
.B1(n_138),
.B2(n_113),
.Y(n_242)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_139),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_131),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_207),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_137),
.A2(n_24),
.B1(n_43),
.B2(n_47),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_113),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_209),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_157),
.A2(n_139),
.B1(n_122),
.B2(n_142),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_214),
.A2(n_217),
.B1(n_231),
.B2(n_252),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_221),
.B(n_171),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_180),
.A2(n_117),
.B1(n_56),
.B2(n_55),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_223),
.A2(n_240),
.B1(n_136),
.B2(n_197),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_180),
.A2(n_145),
.B1(n_142),
.B2(n_135),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_124),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_156),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_242),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_192),
.A2(n_24),
.B1(n_111),
.B2(n_136),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_158),
.B(n_150),
.C(n_61),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_177),
.C(n_153),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_196),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_254),
.B(n_257),
.Y(n_293)
);

OAI22xp33_ASAP7_75t_L g255 ( 
.A1(n_212),
.A2(n_185),
.B1(n_206),
.B2(n_167),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_255),
.A2(n_251),
.B1(n_239),
.B2(n_229),
.Y(n_314)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_211),
.Y(n_256)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_256),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_233),
.B(n_163),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_258),
.B(n_259),
.Y(n_297)
);

AO22x1_ASAP7_75t_SL g259 ( 
.A1(n_240),
.A2(n_156),
.B1(n_183),
.B2(n_202),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_260),
.B(n_265),
.Y(n_322)
);

O2A1O1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_232),
.A2(n_169),
.B(n_187),
.C(n_200),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_261),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_228),
.B(n_176),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_262),
.B(n_226),
.C(n_216),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_210),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_263),
.B(n_264),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_249),
.B(n_13),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_221),
.B(n_188),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_228),
.A2(n_160),
.B(n_170),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_266),
.A2(n_271),
.B(n_281),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_220),
.B(n_160),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_267),
.B(n_268),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_238),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_207),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_270),
.B(n_274),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_228),
.A2(n_170),
.B(n_165),
.Y(n_271)
);

INVx13_ASAP7_75t_L g272 ( 
.A(n_236),
.Y(n_272)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_236),
.Y(n_273)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_273),
.Y(n_326)
);

AND2x6_ASAP7_75t_L g274 ( 
.A(n_223),
.B(n_19),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_241),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_275),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_213),
.B(n_173),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_276),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_240),
.B(n_186),
.Y(n_277)
);

FAx1_ASAP7_75t_SL g310 ( 
.A(n_277),
.B(n_280),
.CI(n_247),
.CON(n_310),
.SN(n_310)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_219),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_278),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_227),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_241),
.B(n_190),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_231),
.A2(n_111),
.B(n_150),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_244),
.Y(n_282)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_282),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_225),
.B(n_153),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_284),
.A2(n_286),
.B(n_290),
.Y(n_325)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_244),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_285),
.A2(n_287),
.B1(n_289),
.B2(n_246),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_234),
.B(n_153),
.Y(n_286)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_230),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_288),
.A2(n_290),
.B1(n_291),
.B2(n_259),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_212),
.A2(n_205),
.B1(n_175),
.B2(n_164),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_250),
.A2(n_41),
.B1(n_22),
.B2(n_44),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_SL g291 ( 
.A(n_253),
.B(n_44),
.C(n_150),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_291),
.A2(n_232),
.B(n_215),
.Y(n_298)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_211),
.Y(n_292)
);

BUFx5_ASAP7_75t_L g309 ( 
.A(n_292),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_295),
.B(n_299),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_288),
.A2(n_217),
.B1(n_252),
.B2(n_243),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_296),
.A2(n_318),
.B1(n_320),
.B2(n_321),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_298),
.Y(n_348)
);

XOR2x2_ASAP7_75t_L g299 ( 
.A(n_262),
.B(n_224),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_301),
.B(n_310),
.Y(n_328)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_302),
.Y(n_334)
);

OAI32xp33_ASAP7_75t_L g304 ( 
.A1(n_254),
.A2(n_250),
.A3(n_226),
.B1(n_216),
.B2(n_222),
.Y(n_304)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_304),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_277),
.A2(n_215),
.B(n_247),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_307),
.A2(n_235),
.B(n_272),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_283),
.A2(n_243),
.B1(n_239),
.B2(n_229),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_313),
.B(n_286),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_314),
.A2(n_315),
.B1(n_287),
.B2(n_292),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_269),
.A2(n_251),
.B1(n_246),
.B2(n_162),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_258),
.B(n_279),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_282),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_265),
.A2(n_230),
.B1(n_235),
.B2(n_245),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_274),
.A2(n_259),
.B1(n_269),
.B2(n_260),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_259),
.A2(n_281),
.B1(n_257),
.B2(n_263),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_323),
.B(n_272),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_266),
.B(n_271),
.C(n_268),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_284),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_329),
.Y(n_371)
);

O2A1O1Ixp33_ASAP7_75t_L g330 ( 
.A1(n_297),
.A2(n_280),
.B(n_275),
.C(n_285),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_330),
.B(n_344),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_331),
.B(n_358),
.Y(n_379)
);

NAND3xp33_ASAP7_75t_L g332 ( 
.A(n_311),
.B(n_264),
.C(n_270),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_332),
.B(n_351),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_293),
.B(n_278),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_333),
.B(n_340),
.Y(n_368)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_309),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_335),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_319),
.A2(n_261),
.B(n_276),
.Y(n_336)
);

AO21x1_ASAP7_75t_L g363 ( 
.A1(n_336),
.A2(n_353),
.B(n_298),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_338),
.B(n_347),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_293),
.B(n_218),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_324),
.Y(n_341)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_341),
.Y(n_372)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_324),
.Y(n_342)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_342),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_343),
.A2(n_355),
.B1(n_296),
.B2(n_320),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_322),
.B(n_261),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_322),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_345),
.B(n_346),
.Y(n_375)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_297),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_312),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_349),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_306),
.B(n_256),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_350),
.B(n_352),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_317),
.B(n_218),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_305),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_315),
.A2(n_245),
.B1(n_44),
.B2(n_67),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_306),
.B(n_41),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_356),
.B(n_357),
.Y(n_377)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_303),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_310),
.B(n_327),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_348),
.A2(n_319),
.B(n_325),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_361),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_354),
.A2(n_321),
.B1(n_314),
.B2(n_300),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_362),
.A2(n_347),
.B1(n_338),
.B2(n_343),
.Y(n_391)
);

AO21x1_ASAP7_75t_L g401 ( 
.A1(n_363),
.A2(n_376),
.B(n_381),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_349),
.B(n_345),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_366),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_331),
.B(n_316),
.C(n_295),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_367),
.B(n_328),
.C(n_301),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_356),
.B(n_308),
.Y(n_369)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_369),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_344),
.B(n_308),
.Y(n_370)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_370),
.Y(n_403)
);

NAND2x1_ASAP7_75t_SL g376 ( 
.A(n_353),
.B(n_310),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_337),
.B(n_358),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_378),
.B(n_338),
.Y(n_398)
);

BUFx5_ASAP7_75t_L g380 ( 
.A(n_335),
.Y(n_380)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_380),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_348),
.A2(n_325),
.B(n_318),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_383),
.A2(n_313),
.B1(n_352),
.B2(n_341),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_339),
.B(n_304),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_384),
.B(n_339),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_337),
.B(n_299),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_385),
.B(n_367),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_383),
.A2(n_354),
.B1(n_346),
.B2(n_374),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_386),
.A2(n_405),
.B1(n_406),
.B2(n_364),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_SL g423 ( 
.A(n_388),
.B(n_375),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_389),
.B(n_407),
.Y(n_412)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_390),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_391),
.A2(n_400),
.B1(n_404),
.B2(n_408),
.Y(n_414)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_373),
.Y(n_395)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_395),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_378),
.B(n_328),
.C(n_336),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_396),
.B(n_379),
.C(n_377),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_365),
.B(n_326),
.Y(n_397)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_397),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_398),
.B(n_381),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_365),
.B(n_366),
.Y(n_399)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_399),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_L g400 ( 
.A1(n_380),
.A2(n_334),
.B1(n_355),
.B2(n_342),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_359),
.B(n_326),
.Y(n_402)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_402),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_362),
.A2(n_364),
.B1(n_361),
.B2(n_371),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_374),
.A2(n_334),
.B1(n_330),
.B2(n_350),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_385),
.B(n_307),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_364),
.A2(n_357),
.B1(n_352),
.B2(n_303),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_410),
.B(n_411),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_393),
.B(n_373),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_413),
.B(n_416),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_392),
.A2(n_371),
.B1(n_363),
.B2(n_376),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_417),
.B(n_421),
.C(n_422),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_394),
.A2(n_368),
.B1(n_375),
.B2(n_377),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_419),
.A2(n_426),
.B1(n_387),
.B2(n_294),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_388),
.B(n_379),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_392),
.A2(n_376),
.B(n_363),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_423),
.B(n_41),
.C(n_22),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_386),
.A2(n_382),
.B1(n_372),
.B2(n_360),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_424),
.Y(n_436)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_403),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_398),
.B(n_382),
.Y(n_427)
);

XOR2x2_ASAP7_75t_L g431 ( 
.A(n_427),
.B(n_405),
.Y(n_431)
);

OAI322xp33_ASAP7_75t_L g428 ( 
.A1(n_411),
.A2(n_396),
.A3(n_404),
.B1(n_401),
.B2(n_389),
.C1(n_407),
.C2(n_408),
.Y(n_428)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_428),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_416),
.A2(n_401),
.B(n_391),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_430),
.A2(n_438),
.B(n_414),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_431),
.B(n_439),
.Y(n_443)
);

A2O1A1O1Ixp25_ASAP7_75t_L g433 ( 
.A1(n_422),
.A2(n_395),
.B(n_372),
.C(n_387),
.D(n_360),
.Y(n_433)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_433),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_435),
.B(n_440),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_409),
.A2(n_294),
.B1(n_309),
.B2(n_2),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_437),
.A2(n_442),
.B1(n_0),
.B2(n_5),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_420),
.A2(n_41),
.B(n_22),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_412),
.B(n_41),
.C(n_1),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_412),
.B(n_0),
.C(n_2),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_441),
.B(n_418),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_425),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_430),
.A2(n_410),
.B(n_415),
.Y(n_445)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_445),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_446),
.B(n_447),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_434),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_436),
.A2(n_424),
.B1(n_414),
.B2(n_417),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_448),
.A2(n_454),
.B1(n_439),
.B2(n_8),
.Y(n_462)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_449),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_432),
.B(n_413),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_450),
.B(n_453),
.C(n_429),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_432),
.A2(n_427),
.B(n_423),
.Y(n_452)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_452),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_429),
.B(n_421),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_456),
.B(n_462),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_455),
.A2(n_436),
.B1(n_431),
.B2(n_433),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_457),
.B(n_460),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_440),
.C(n_441),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_453),
.B(n_6),
.C(n_8),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_463),
.A2(n_465),
.B(n_461),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_450),
.B(n_448),
.C(n_443),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_466),
.B(n_467),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_456),
.A2(n_452),
.B(n_451),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_459),
.A2(n_445),
.B1(n_443),
.B2(n_9),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_468),
.B(n_463),
.Y(n_473)
);

OAI21x1_ASAP7_75t_L g469 ( 
.A1(n_464),
.A2(n_6),
.B(n_8),
.Y(n_469)
);

AOI31xp67_ASAP7_75t_L g475 ( 
.A1(n_469),
.A2(n_9),
.A3(n_10),
.B(n_11),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_470),
.B(n_465),
.C(n_458),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_472),
.A2(n_474),
.B(n_470),
.Y(n_477)
);

AOI21x1_ASAP7_75t_L g476 ( 
.A1(n_473),
.A2(n_475),
.B(n_471),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_476),
.B(n_477),
.C(n_9),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_478),
.B(n_9),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g480 ( 
.A(n_479),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_480),
.A2(n_10),
.B(n_12),
.Y(n_481)
);

OR2x2_ASAP7_75t_L g482 ( 
.A(n_481),
.B(n_10),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_482),
.B(n_12),
.Y(n_483)
);


endmodule