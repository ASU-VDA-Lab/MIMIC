module fake_aes_10005_n_38 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_38);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NAND2xp5_ASAP7_75t_L g12 ( .A(n_1), .B(n_4), .Y(n_12) );
NOR2xp67_ASAP7_75t_L g13 ( .A(n_7), .B(n_5), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_8), .B(n_5), .Y(n_14) );
NAND2xp33_ASAP7_75t_L g15 ( .A(n_3), .B(n_8), .Y(n_15) );
OAI21x1_ASAP7_75t_L g16 ( .A1(n_4), .A2(n_7), .B(n_6), .Y(n_16) );
BUFx6f_ASAP7_75t_L g17 ( .A(n_10), .Y(n_17) );
NAND2xp5_ASAP7_75t_SL g18 ( .A(n_17), .B(n_0), .Y(n_18) );
BUFx2_ASAP7_75t_L g19 ( .A(n_14), .Y(n_19) );
NAND2xp5_ASAP7_75t_SL g20 ( .A(n_17), .B(n_0), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_18), .Y(n_21) );
AOI21xp5_ASAP7_75t_L g22 ( .A1(n_19), .A2(n_17), .B(n_12), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_21), .B(n_14), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_21), .B(n_16), .Y(n_24) );
BUFx2_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
INVx2_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g27 ( .A(n_25), .B(n_23), .Y(n_27) );
HB1xp67_ASAP7_75t_L g28 ( .A(n_26), .Y(n_28) );
AOI22xp5_ASAP7_75t_L g29 ( .A1(n_27), .A2(n_15), .B1(n_22), .B2(n_20), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
NOR2x1_ASAP7_75t_L g31 ( .A(n_27), .B(n_13), .Y(n_31) );
AOI21xp33_ASAP7_75t_SL g32 ( .A1(n_30), .A2(n_16), .B(n_2), .Y(n_32) );
NOR3xp33_ASAP7_75t_L g33 ( .A(n_31), .B(n_13), .C(n_2), .Y(n_33) );
AOI21xp5_ASAP7_75t_L g34 ( .A1(n_29), .A2(n_17), .B(n_9), .Y(n_34) );
AOI22x1_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_17), .B1(n_3), .B2(n_6), .Y(n_35) );
AND2x2_ASAP7_75t_L g36 ( .A(n_33), .B(n_17), .Y(n_36) );
OAI31xp33_ASAP7_75t_L g37 ( .A1(n_36), .A2(n_32), .A3(n_1), .B(n_11), .Y(n_37) );
AOI22xp5_ASAP7_75t_SL g38 ( .A1(n_37), .A2(n_35), .B1(n_36), .B2(n_30), .Y(n_38) );
endmodule