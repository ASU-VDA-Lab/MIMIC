module real_aes_6588_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_166;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g176 ( .A1(n_0), .A2(n_177), .B(n_180), .C(n_184), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_1), .B(n_168), .Y(n_187) );
INVx1_ASAP7_75t_L g110 ( .A(n_2), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_3), .B(n_178), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_4), .A2(n_137), .B(n_507), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_5), .A2(n_142), .B(n_145), .C(n_534), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_6), .A2(n_137), .B(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_7), .B(n_168), .Y(n_513) );
AO21x2_ASAP7_75t_L g244 ( .A1(n_8), .A2(n_170), .B(n_245), .Y(n_244) );
AND2x6_ASAP7_75t_L g142 ( .A(n_9), .B(n_143), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_10), .A2(n_142), .B(n_145), .C(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g547 ( .A(n_11), .Y(n_547) );
INVx1_ASAP7_75t_L g108 ( .A(n_12), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_12), .B(n_43), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_13), .B(n_183), .Y(n_536) );
INVx1_ASAP7_75t_L g163 ( .A(n_14), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_15), .B(n_178), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g566 ( .A1(n_16), .A2(n_179), .B(n_567), .C(n_569), .Y(n_566) );
XOR2xp5_ASAP7_75t_L g120 ( .A(n_17), .B(n_121), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_17), .B(n_168), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_18), .B(n_451), .Y(n_450) );
AOI222xp33_ASAP7_75t_SL g453 ( .A1(n_19), .A2(n_454), .B1(n_455), .B2(n_464), .C1(n_731), .C2(n_732), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_20), .B(n_157), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_L g144 ( .A1(n_21), .A2(n_145), .B(n_148), .C(n_156), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g554 ( .A1(n_22), .A2(n_182), .B(n_238), .C(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_23), .B(n_183), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_24), .A2(n_42), .B1(n_461), .B2(n_462), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_24), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_25), .B(n_183), .Y(n_521) );
CKINVDCx16_ASAP7_75t_R g481 ( .A(n_26), .Y(n_481) );
INVx1_ASAP7_75t_L g520 ( .A(n_27), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_28), .A2(n_145), .B(n_156), .C(n_248), .Y(n_247) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_29), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_30), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g124 ( .A1(n_31), .A2(n_80), .B1(n_125), .B2(n_126), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_31), .Y(n_126) );
INVx1_ASAP7_75t_L g498 ( .A(n_32), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_33), .A2(n_137), .B(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g140 ( .A(n_34), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g195 ( .A1(n_35), .A2(n_196), .B(n_197), .C(n_201), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_36), .Y(n_538) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_37), .A2(n_182), .B(n_510), .C(n_512), .Y(n_509) );
INVxp67_ASAP7_75t_L g499 ( .A(n_38), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_39), .B(n_250), .Y(n_249) );
CKINVDCx14_ASAP7_75t_R g508 ( .A(n_40), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_41), .A2(n_145), .B(n_156), .C(n_519), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_42), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_43), .B(n_108), .Y(n_107) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_44), .A2(n_184), .B(n_545), .C(n_546), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_45), .B(n_136), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g241 ( .A(n_46), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_47), .B(n_178), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_48), .B(n_137), .Y(n_246) );
OAI22xp5_ASAP7_75t_SL g455 ( .A1(n_49), .A2(n_456), .B1(n_457), .B2(n_463), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_49), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_50), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_51), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_52), .A2(n_196), .B(n_201), .C(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g181 ( .A(n_53), .Y(n_181) );
INVx1_ASAP7_75t_L g224 ( .A(n_54), .Y(n_224) );
INVx1_ASAP7_75t_L g553 ( .A(n_55), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_56), .B(n_137), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_57), .Y(n_165) );
CKINVDCx14_ASAP7_75t_R g543 ( .A(n_58), .Y(n_543) );
INVx1_ASAP7_75t_L g143 ( .A(n_59), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_60), .B(n_137), .Y(n_269) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_61), .A2(n_105), .B1(n_114), .B2(n_738), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_62), .B(n_168), .Y(n_215) );
A2O1A1Ixp33_ASAP7_75t_L g210 ( .A1(n_63), .A2(n_155), .B(n_211), .C(n_213), .Y(n_210) );
INVx1_ASAP7_75t_L g162 ( .A(n_64), .Y(n_162) );
INVx1_ASAP7_75t_SL g511 ( .A(n_65), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_66), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_67), .B(n_178), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_68), .B(n_168), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_69), .B(n_179), .Y(n_235) );
INVx1_ASAP7_75t_L g484 ( .A(n_70), .Y(n_484) );
CKINVDCx16_ASAP7_75t_R g174 ( .A(n_71), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_72), .B(n_150), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g263 ( .A1(n_73), .A2(n_145), .B(n_201), .C(n_264), .Y(n_263) );
CKINVDCx16_ASAP7_75t_R g209 ( .A(n_74), .Y(n_209) );
INVx1_ASAP7_75t_L g113 ( .A(n_75), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_76), .A2(n_137), .B(n_542), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_77), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_78), .A2(n_137), .B(n_564), .Y(n_563) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_79), .A2(n_123), .B1(n_124), .B2(n_127), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_79), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_80), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_81), .A2(n_136), .B(n_494), .Y(n_493) );
CKINVDCx16_ASAP7_75t_R g517 ( .A(n_82), .Y(n_517) );
INVx1_ASAP7_75t_L g565 ( .A(n_83), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_84), .B(n_153), .Y(n_152) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_85), .A2(n_458), .B1(n_459), .B2(n_460), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_85), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_86), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_87), .A2(n_137), .B(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g568 ( .A(n_88), .Y(n_568) );
INVx2_ASAP7_75t_L g160 ( .A(n_89), .Y(n_160) );
INVx1_ASAP7_75t_L g535 ( .A(n_90), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g271 ( .A(n_91), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_92), .B(n_183), .Y(n_236) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_93), .B(n_110), .C(n_111), .Y(n_109) );
OR2x2_ASAP7_75t_L g446 ( .A(n_93), .B(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g467 ( .A(n_93), .B(n_448), .Y(n_467) );
INVx2_ASAP7_75t_L g469 ( .A(n_93), .Y(n_469) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_94), .A2(n_145), .B(n_201), .C(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_95), .B(n_137), .Y(n_194) );
INVx1_ASAP7_75t_L g198 ( .A(n_96), .Y(n_198) );
INVxp67_ASAP7_75t_L g214 ( .A(n_97), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_98), .B(n_170), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_99), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g231 ( .A(n_100), .Y(n_231) );
INVx1_ASAP7_75t_L g265 ( .A(n_101), .Y(n_265) );
INVx2_ASAP7_75t_L g556 ( .A(n_102), .Y(n_556) );
AND2x2_ASAP7_75t_L g226 ( .A(n_103), .B(n_159), .Y(n_226) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
BUFx2_ASAP7_75t_L g738 ( .A(n_106), .Y(n_738) );
OR2x4_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
AND2x2_ASAP7_75t_L g448 ( .A(n_110), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
OA21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_119), .B(n_452), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g737 ( .A(n_118), .Y(n_737) );
OAI21xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_443), .B(n_450), .Y(n_119) );
AOI22xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_128), .B1(n_441), .B2(n_442), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_122), .Y(n_441) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g442 ( .A(n_128), .Y(n_442) );
OAI22xp5_ASAP7_75t_SL g732 ( .A1(n_128), .A2(n_733), .B1(n_734), .B2(n_735), .Y(n_732) );
AND2x2_ASAP7_75t_SL g128 ( .A(n_129), .B(n_377), .Y(n_128) );
NOR5xp2_ASAP7_75t_L g129 ( .A(n_130), .B(n_308), .C(n_337), .D(n_357), .E(n_364), .Y(n_129) );
OAI211xp5_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_188), .B(n_252), .C(n_295), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_132), .A2(n_380), .B1(n_382), .B2(n_383), .Y(n_379) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_167), .Y(n_132) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_133), .Y(n_255) );
AND2x4_ASAP7_75t_L g288 ( .A(n_133), .B(n_289), .Y(n_288) );
INVx5_ASAP7_75t_L g306 ( .A(n_133), .Y(n_306) );
AND2x2_ASAP7_75t_L g315 ( .A(n_133), .B(n_307), .Y(n_315) );
AND2x2_ASAP7_75t_L g327 ( .A(n_133), .B(n_192), .Y(n_327) );
AND2x2_ASAP7_75t_L g423 ( .A(n_133), .B(n_291), .Y(n_423) );
OR2x6_ASAP7_75t_L g133 ( .A(n_134), .B(n_164), .Y(n_133) );
AOI21xp5_ASAP7_75t_SL g134 ( .A1(n_135), .A2(n_144), .B(n_157), .Y(n_134) );
BUFx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_142), .Y(n_137) );
NAND2x1p5_ASAP7_75t_L g232 ( .A(n_138), .B(n_142), .Y(n_232) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_141), .Y(n_138) );
INVx1_ASAP7_75t_L g155 ( .A(n_139), .Y(n_155) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g146 ( .A(n_140), .Y(n_146) );
INVx1_ASAP7_75t_L g239 ( .A(n_140), .Y(n_239) );
INVx1_ASAP7_75t_L g147 ( .A(n_141), .Y(n_147) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_141), .Y(n_151) );
INVx3_ASAP7_75t_L g179 ( .A(n_141), .Y(n_179) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_141), .Y(n_183) );
INVx1_ASAP7_75t_L g250 ( .A(n_141), .Y(n_250) );
BUFx3_ASAP7_75t_L g156 ( .A(n_142), .Y(n_156) );
INVx4_ASAP7_75t_SL g186 ( .A(n_142), .Y(n_186) );
INVx5_ASAP7_75t_L g175 ( .A(n_145), .Y(n_175) );
AND2x6_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
BUFx3_ASAP7_75t_L g185 ( .A(n_146), .Y(n_185) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_146), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_152), .B(n_154), .Y(n_148) );
INVx2_ASAP7_75t_L g153 ( .A(n_150), .Y(n_153) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx4_ASAP7_75t_L g212 ( .A(n_151), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g197 ( .A1(n_153), .A2(n_198), .B(n_199), .C(n_200), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g223 ( .A1(n_153), .A2(n_200), .B(n_224), .C(n_225), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_L g483 ( .A1(n_153), .A2(n_484), .B(n_485), .C(n_486), .Y(n_483) );
O2A1O1Ixp5_ASAP7_75t_L g534 ( .A1(n_153), .A2(n_486), .B(n_535), .C(n_536), .Y(n_534) );
O2A1O1Ixp33_ASAP7_75t_L g519 ( .A1(n_154), .A2(n_178), .B(n_520), .C(n_521), .Y(n_519) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_155), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_158), .B(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g166 ( .A(n_159), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_159), .A2(n_194), .B(n_195), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_159), .A2(n_221), .B(n_222), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_L g516 ( .A1(n_159), .A2(n_232), .B(n_517), .C(n_518), .Y(n_516) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_159), .A2(n_541), .B(n_548), .Y(n_540) );
AND2x2_ASAP7_75t_SL g159 ( .A(n_160), .B(n_161), .Y(n_159) );
AND2x2_ASAP7_75t_L g171 ( .A(n_160), .B(n_161), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_162), .B(n_163), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_166), .A2(n_531), .B(n_537), .Y(n_530) );
INVx2_ASAP7_75t_L g289 ( .A(n_167), .Y(n_289) );
AND2x2_ASAP7_75t_L g307 ( .A(n_167), .B(n_261), .Y(n_307) );
AND2x2_ASAP7_75t_L g326 ( .A(n_167), .B(n_260), .Y(n_326) );
AND2x2_ASAP7_75t_L g366 ( .A(n_167), .B(n_306), .Y(n_366) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_172), .B(n_187), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_169), .B(n_203), .Y(n_202) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_169), .A2(n_230), .B(n_240), .Y(n_229) );
AO21x2_ASAP7_75t_L g261 ( .A1(n_169), .A2(n_262), .B(n_270), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_169), .B(n_271), .Y(n_270) );
AO21x2_ASAP7_75t_L g479 ( .A1(n_169), .A2(n_480), .B(n_487), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_169), .B(n_523), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_169), .B(n_538), .Y(n_537) );
INVx4_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_170), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_170), .A2(n_246), .B(n_247), .Y(n_245) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g242 ( .A(n_171), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_SL g173 ( .A1(n_174), .A2(n_175), .B(n_176), .C(n_186), .Y(n_173) );
INVx2_ASAP7_75t_L g196 ( .A(n_175), .Y(n_196) );
O2A1O1Ixp33_ASAP7_75t_L g208 ( .A1(n_175), .A2(n_186), .B(n_209), .C(n_210), .Y(n_208) );
O2A1O1Ixp33_ASAP7_75t_SL g494 ( .A1(n_175), .A2(n_186), .B(n_495), .C(n_496), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_L g507 ( .A1(n_175), .A2(n_186), .B(n_508), .C(n_509), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_SL g542 ( .A1(n_175), .A2(n_186), .B(n_543), .C(n_544), .Y(n_542) );
O2A1O1Ixp33_ASAP7_75t_SL g552 ( .A1(n_175), .A2(n_186), .B(n_553), .C(n_554), .Y(n_552) );
O2A1O1Ixp33_ASAP7_75t_SL g564 ( .A1(n_175), .A2(n_186), .B(n_565), .C(n_566), .Y(n_564) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_178), .B(n_214), .Y(n_213) );
OAI22xp33_ASAP7_75t_L g497 ( .A1(n_178), .A2(n_212), .B1(n_498), .B2(n_499), .Y(n_497) );
INVx5_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_179), .B(n_547), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_182), .B(n_511), .Y(n_510) );
INVx4_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g545 ( .A(n_183), .Y(n_545) );
INVx2_ASAP7_75t_L g486 ( .A(n_184), .Y(n_486) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_185), .Y(n_200) );
INVx1_ASAP7_75t_L g569 ( .A(n_185), .Y(n_569) );
INVx1_ASAP7_75t_L g201 ( .A(n_186), .Y(n_201) );
INVxp67_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_190), .B(n_216), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AOI322xp5_ASAP7_75t_L g425 ( .A1(n_191), .A2(n_227), .A3(n_280), .B1(n_288), .B2(n_342), .C1(n_426), .C2(n_429), .Y(n_425) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_204), .Y(n_191) );
INVx5_ASAP7_75t_L g257 ( .A(n_192), .Y(n_257) );
AND2x2_ASAP7_75t_L g274 ( .A(n_192), .B(n_259), .Y(n_274) );
BUFx2_ASAP7_75t_L g352 ( .A(n_192), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_192), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g429 ( .A(n_192), .B(n_336), .Y(n_429) );
OR2x6_ASAP7_75t_L g192 ( .A(n_193), .B(n_202), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_204), .B(n_218), .Y(n_283) );
INVx1_ASAP7_75t_L g310 ( .A(n_204), .Y(n_310) );
AND2x2_ASAP7_75t_L g323 ( .A(n_204), .B(n_243), .Y(n_323) );
AND2x2_ASAP7_75t_L g424 ( .A(n_204), .B(n_342), .Y(n_424) );
INVx3_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
OR2x2_ASAP7_75t_L g278 ( .A(n_205), .B(n_218), .Y(n_278) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_205), .Y(n_286) );
OR2x2_ASAP7_75t_L g293 ( .A(n_205), .B(n_243), .Y(n_293) );
AND2x2_ASAP7_75t_L g303 ( .A(n_205), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_205), .B(n_229), .Y(n_332) );
INVxp67_ASAP7_75t_L g356 ( .A(n_205), .Y(n_356) );
AND2x2_ASAP7_75t_L g363 ( .A(n_205), .B(n_227), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_205), .B(n_243), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_205), .B(n_228), .Y(n_389) );
OA21x2_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_215), .Y(n_205) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_206), .A2(n_506), .B(n_513), .Y(n_505) );
OA21x2_ASAP7_75t_L g550 ( .A1(n_206), .A2(n_551), .B(n_557), .Y(n_550) );
OA21x2_ASAP7_75t_L g562 ( .A1(n_206), .A2(n_563), .B(n_570), .Y(n_562) );
O2A1O1Ixp33_ASAP7_75t_L g264 ( .A1(n_211), .A2(n_265), .B(n_266), .C(n_267), .Y(n_264) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_212), .B(n_556), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_212), .B(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_227), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_218), .B(n_244), .Y(n_333) );
OR2x2_ASAP7_75t_L g355 ( .A(n_218), .B(n_228), .Y(n_355) );
AND2x2_ASAP7_75t_L g368 ( .A(n_218), .B(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_218), .B(n_323), .Y(n_374) );
OAI211xp5_ASAP7_75t_SL g378 ( .A1(n_218), .A2(n_379), .B(n_384), .C(n_393), .Y(n_378) );
AND2x2_ASAP7_75t_L g439 ( .A(n_218), .B(n_243), .Y(n_439) );
INVx5_ASAP7_75t_SL g218 ( .A(n_219), .Y(n_218) );
OR2x2_ASAP7_75t_L g292 ( .A(n_219), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_219), .B(n_298), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_219), .B(n_287), .Y(n_299) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_219), .Y(n_301) );
OR2x2_ASAP7_75t_L g312 ( .A(n_219), .B(n_228), .Y(n_312) );
AND2x2_ASAP7_75t_SL g317 ( .A(n_219), .B(n_303), .Y(n_317) );
AND2x2_ASAP7_75t_L g342 ( .A(n_219), .B(n_228), .Y(n_342) );
AND2x2_ASAP7_75t_L g362 ( .A(n_219), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g400 ( .A(n_219), .B(n_227), .Y(n_400) );
OR2x2_ASAP7_75t_L g403 ( .A(n_219), .B(n_389), .Y(n_403) );
OR2x6_ASAP7_75t_L g219 ( .A(n_220), .B(n_226), .Y(n_219) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_243), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g346 ( .A1(n_228), .A2(n_347), .B(n_350), .C(n_356), .Y(n_346) );
INVx5_ASAP7_75t_SL g228 ( .A(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_229), .B(n_243), .Y(n_277) );
AND2x2_ASAP7_75t_L g281 ( .A(n_229), .B(n_244), .Y(n_281) );
OR2x2_ASAP7_75t_L g287 ( .A(n_229), .B(n_243), .Y(n_287) );
OAI21xp5_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_233), .Y(n_230) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_232), .A2(n_481), .B(n_482), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_232), .A2(n_532), .B(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B(n_237), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_237), .A2(n_249), .B(n_251), .Y(n_248) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx3_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
INVx2_ASAP7_75t_L g491 ( .A(n_242), .Y(n_491) );
INVx1_ASAP7_75t_SL g304 ( .A(n_243), .Y(n_304) );
OR2x2_ASAP7_75t_L g432 ( .A(n_243), .B(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_272), .B(n_275), .C(n_284), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AOI31xp33_ASAP7_75t_L g357 ( .A1(n_254), .A2(n_358), .A3(n_360), .B(n_361), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_255), .B(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_256), .B(n_288), .Y(n_294) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_257), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g314 ( .A(n_257), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g319 ( .A(n_257), .B(n_289), .Y(n_319) );
AND2x2_ASAP7_75t_L g329 ( .A(n_257), .B(n_288), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_257), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g349 ( .A(n_257), .B(n_306), .Y(n_349) );
AND2x2_ASAP7_75t_L g354 ( .A(n_257), .B(n_326), .Y(n_354) );
OR2x2_ASAP7_75t_L g373 ( .A(n_257), .B(n_259), .Y(n_373) );
OR2x2_ASAP7_75t_L g375 ( .A(n_257), .B(n_376), .Y(n_375) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_257), .Y(n_422) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g322 ( .A(n_259), .B(n_289), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_259), .B(n_306), .Y(n_345) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
BUFx2_ASAP7_75t_L g291 ( .A(n_261), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_269), .Y(n_262) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx3_ASAP7_75t_L g512 ( .A(n_268), .Y(n_512) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g382 ( .A(n_274), .B(n_306), .Y(n_382) );
AOI322xp5_ASAP7_75t_L g384 ( .A1(n_274), .A2(n_288), .A3(n_326), .B1(n_385), .B2(n_386), .C1(n_387), .C2(n_390), .Y(n_384) );
INVx1_ASAP7_75t_L g392 ( .A(n_274), .Y(n_392) );
NAND2xp33_ASAP7_75t_L g275 ( .A(n_276), .B(n_279), .Y(n_275) );
INVx1_ASAP7_75t_SL g386 ( .A(n_276), .Y(n_386) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
OR2x2_ASAP7_75t_L g338 ( .A(n_277), .B(n_283), .Y(n_338) );
INVx1_ASAP7_75t_L g369 ( .A(n_277), .Y(n_369) );
INVx2_ASAP7_75t_SL g279 ( .A(n_280), .Y(n_279) );
AND2x4_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OAI32xp33_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_288), .A3(n_290), .B1(n_292), .B2(n_294), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
AOI21xp33_ASAP7_75t_SL g324 ( .A1(n_287), .A2(n_302), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_SL g339 ( .A(n_288), .Y(n_339) );
AND2x4_ASAP7_75t_L g336 ( .A(n_289), .B(n_306), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_289), .B(n_372), .Y(n_371) );
AOI322xp5_ASAP7_75t_L g401 ( .A1(n_290), .A2(n_317), .A3(n_336), .B1(n_369), .B2(n_402), .C1(n_404), .C2(n_405), .Y(n_401) );
OAI221xp5_ASAP7_75t_L g430 ( .A1(n_290), .A2(n_367), .B1(n_431), .B2(n_432), .C(n_434), .Y(n_430) );
AND2x2_ASAP7_75t_L g318 ( .A(n_291), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_SL g298 ( .A(n_293), .Y(n_298) );
OR2x2_ASAP7_75t_L g370 ( .A(n_293), .B(n_355), .Y(n_370) );
OAI31xp33_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_299), .A3(n_300), .B(n_305), .Y(n_295) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_296), .A2(n_329), .B1(n_330), .B2(n_334), .Y(n_328) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g341 ( .A(n_298), .B(n_342), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_300), .A2(n_341), .B1(n_394), .B2(n_397), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g383 ( .A(n_303), .B(n_352), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_303), .B(n_342), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_304), .B(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g417 ( .A(n_304), .B(n_355), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_305), .A2(n_400), .B1(n_413), .B2(n_416), .Y(n_412) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx2_ASAP7_75t_L g321 ( .A(n_306), .Y(n_321) );
AND2x2_ASAP7_75t_L g404 ( .A(n_306), .B(n_326), .Y(n_404) );
OR2x2_ASAP7_75t_L g406 ( .A(n_306), .B(n_373), .Y(n_406) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_306), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_307), .B(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_307), .B(n_352), .Y(n_360) );
OAI211xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_313), .B(n_316), .C(n_328), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AOI221xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_318), .B1(n_320), .B2(n_323), .C(n_324), .Y(n_316) );
INVxp67_ASAP7_75t_L g428 ( .A(n_319), .Y(n_428) );
INVx1_ASAP7_75t_L g395 ( .A(n_320), .Y(n_395) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
AND2x2_ASAP7_75t_L g359 ( .A(n_321), .B(n_326), .Y(n_359) );
INVx1_ASAP7_75t_L g376 ( .A(n_322), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_322), .B(n_349), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVx1_ASAP7_75t_L g391 ( .A(n_326), .Y(n_391) );
AND2x2_ASAP7_75t_L g397 ( .A(n_326), .B(n_352), .Y(n_397) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx1_ASAP7_75t_SL g385 ( .A(n_333), .Y(n_385) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_336), .B(n_372), .Y(n_396) );
OAI221xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_339), .B1(n_340), .B2(n_343), .C(n_346), .Y(n_337) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g433 ( .A(n_342), .Y(n_433) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g351 ( .A(n_345), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_349), .B(n_408), .Y(n_407) );
AOI21xp33_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_353), .B(n_355), .Y(n_350) );
OAI211xp5_ASAP7_75t_SL g398 ( .A1(n_353), .A2(n_399), .B(n_401), .C(n_407), .Y(n_398) );
INVx1_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g410 ( .A(n_355), .Y(n_410) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI222xp33_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_367), .B1(n_370), .B2(n_371), .C1(n_374), .C2(n_375), .Y(n_364) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g440 ( .A(n_371), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_372), .B(n_415), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_372), .A2(n_419), .B1(n_421), .B2(n_424), .Y(n_418) );
INVx2_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
NOR4xp25_ASAP7_75t_L g377 ( .A(n_378), .B(n_398), .C(n_411), .D(n_430), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_380), .B(n_410), .Y(n_420) );
INVx1_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g387 ( .A(n_385), .B(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_388), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NAND3xp33_ASAP7_75t_L g411 ( .A(n_412), .B(n_418), .C(n_425), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
INVx2_ASAP7_75t_L g427 ( .A(n_423), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
OAI21xp5_ASAP7_75t_SL g434 ( .A1(n_435), .A2(n_437), .B(n_440), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_442), .A2(n_465), .B1(n_468), .B2(n_470), .Y(n_464) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_SL g451 ( .A(n_446), .Y(n_451) );
NOR2x2_ASAP7_75t_L g731 ( .A(n_447), .B(n_469), .Y(n_731) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g468 ( .A(n_448), .B(n_469), .Y(n_468) );
NAND3xp33_ASAP7_75t_L g452 ( .A(n_450), .B(n_453), .C(n_737), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g733 ( .A(n_466), .Y(n_733) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g736 ( .A(n_468), .Y(n_736) );
INVx2_ASAP7_75t_L g734 ( .A(n_470), .Y(n_734) );
OR2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_665), .Y(n_470) );
NAND5xp2_ASAP7_75t_L g471 ( .A(n_472), .B(n_594), .C(n_624), .D(n_645), .E(n_651), .Y(n_471) );
AOI221xp5_ASAP7_75t_SL g472 ( .A1(n_473), .A2(n_527), .B1(n_558), .B2(n_560), .C(n_571), .Y(n_472) );
INVxp67_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_524), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_476), .B(n_502), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_SL g645 ( .A1(n_477), .A2(n_514), .B(n_646), .C(n_649), .Y(n_645) );
AND2x2_ASAP7_75t_L g715 ( .A(n_477), .B(n_515), .Y(n_715) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_489), .Y(n_477) );
AND2x2_ASAP7_75t_L g573 ( .A(n_478), .B(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g577 ( .A(n_478), .B(n_574), .Y(n_577) );
OR2x2_ASAP7_75t_L g603 ( .A(n_478), .B(n_515), .Y(n_603) );
AND2x2_ASAP7_75t_L g605 ( .A(n_478), .B(n_505), .Y(n_605) );
AND2x2_ASAP7_75t_L g623 ( .A(n_478), .B(n_504), .Y(n_623) );
INVx1_ASAP7_75t_L g656 ( .A(n_478), .Y(n_656) );
INVx2_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
BUFx2_ASAP7_75t_L g526 ( .A(n_479), .Y(n_526) );
AND2x2_ASAP7_75t_L g559 ( .A(n_479), .B(n_505), .Y(n_559) );
AND2x2_ASAP7_75t_L g712 ( .A(n_479), .B(n_515), .Y(n_712) );
AND2x2_ASAP7_75t_L g593 ( .A(n_489), .B(n_503), .Y(n_593) );
OR2x2_ASAP7_75t_L g597 ( .A(n_489), .B(n_515), .Y(n_597) );
AND2x2_ASAP7_75t_L g622 ( .A(n_489), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_SL g669 ( .A(n_489), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_489), .B(n_631), .Y(n_717) );
AO21x2_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_492), .B(n_500), .Y(n_489) );
INVx1_ASAP7_75t_L g575 ( .A(n_490), .Y(n_575) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OA21x2_ASAP7_75t_L g574 ( .A1(n_493), .A2(n_501), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
OAI322xp33_ASAP7_75t_L g718 ( .A1(n_502), .A2(n_654), .A3(n_677), .B1(n_698), .B2(n_719), .C1(n_721), .C2(n_722), .Y(n_718) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_503), .B(n_574), .Y(n_721) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_514), .Y(n_503) );
AND2x2_ASAP7_75t_L g525 ( .A(n_504), .B(n_526), .Y(n_525) );
AND2x4_ASAP7_75t_L g590 ( .A(n_504), .B(n_515), .Y(n_590) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g631 ( .A(n_505), .B(n_515), .Y(n_631) );
AND2x2_ASAP7_75t_L g675 ( .A(n_505), .B(n_514), .Y(n_675) );
AND2x2_ASAP7_75t_L g558 ( .A(n_514), .B(n_559), .Y(n_558) );
OR2x2_ASAP7_75t_L g576 ( .A(n_514), .B(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_514), .B(n_605), .Y(n_729) );
INVx3_ASAP7_75t_SL g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g524 ( .A(n_515), .B(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_515), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g643 ( .A(n_515), .B(n_574), .Y(n_643) );
AND2x2_ASAP7_75t_L g670 ( .A(n_515), .B(n_605), .Y(n_670) );
OR2x2_ASAP7_75t_L g726 ( .A(n_515), .B(n_577), .Y(n_726) );
OR2x6_ASAP7_75t_L g515 ( .A(n_516), .B(n_522), .Y(n_515) );
INVx1_ASAP7_75t_SL g612 ( .A(n_524), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_525), .B(n_643), .Y(n_644) );
AND2x2_ASAP7_75t_L g678 ( .A(n_525), .B(n_668), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_525), .B(n_601), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_525), .B(n_723), .Y(n_722) );
OAI31xp33_ASAP7_75t_L g696 ( .A1(n_527), .A2(n_558), .A3(n_697), .B(n_699), .Y(n_696) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_539), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_528), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g679 ( .A(n_528), .B(n_614), .Y(n_679) );
OR2x2_ASAP7_75t_L g686 ( .A(n_528), .B(n_687), .Y(n_686) );
OR2x2_ASAP7_75t_L g698 ( .A(n_528), .B(n_587), .Y(n_698) );
CKINVDCx16_ASAP7_75t_R g528 ( .A(n_529), .Y(n_528) );
OR2x2_ASAP7_75t_L g632 ( .A(n_529), .B(n_633), .Y(n_632) );
BUFx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g560 ( .A(n_530), .B(n_561), .Y(n_560) );
INVx4_ASAP7_75t_L g581 ( .A(n_530), .Y(n_581) );
AND2x2_ASAP7_75t_L g618 ( .A(n_530), .B(n_562), .Y(n_618) );
AND2x2_ASAP7_75t_L g617 ( .A(n_539), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_SL g687 ( .A(n_539), .Y(n_687) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_549), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_540), .B(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g587 ( .A(n_540), .B(n_550), .Y(n_587) );
INVx2_ASAP7_75t_L g607 ( .A(n_540), .Y(n_607) );
AND2x2_ASAP7_75t_L g621 ( .A(n_540), .B(n_550), .Y(n_621) );
AND2x2_ASAP7_75t_L g628 ( .A(n_540), .B(n_584), .Y(n_628) );
BUFx3_ASAP7_75t_L g638 ( .A(n_540), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_540), .B(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g583 ( .A(n_549), .Y(n_583) );
AND2x2_ASAP7_75t_L g591 ( .A(n_549), .B(n_581), .Y(n_591) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g561 ( .A(n_550), .B(n_562), .Y(n_561) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_550), .Y(n_615) );
INVx2_ASAP7_75t_SL g598 ( .A(n_559), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_559), .B(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_559), .B(n_668), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g691 ( .A(n_560), .B(n_638), .Y(n_691) );
INVx1_ASAP7_75t_SL g725 ( .A(n_560), .Y(n_725) );
INVx1_ASAP7_75t_SL g633 ( .A(n_561), .Y(n_633) );
INVx1_ASAP7_75t_SL g584 ( .A(n_562), .Y(n_584) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_562), .Y(n_595) );
OR2x2_ASAP7_75t_L g606 ( .A(n_562), .B(n_581), .Y(n_606) );
AND2x2_ASAP7_75t_L g620 ( .A(n_562), .B(n_581), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_562), .B(n_610), .Y(n_672) );
A2O1A1Ixp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_576), .B(n_578), .C(n_589), .Y(n_571) );
AOI31xp33_ASAP7_75t_L g688 ( .A1(n_572), .A2(n_689), .A3(n_690), .B(n_691), .Y(n_688) );
AND2x2_ASAP7_75t_L g661 ( .A(n_573), .B(n_590), .Y(n_661) );
BUFx3_ASAP7_75t_L g601 ( .A(n_574), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_574), .B(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g637 ( .A(n_574), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_574), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_SL g592 ( .A(n_577), .Y(n_592) );
OAI222xp33_ASAP7_75t_L g701 ( .A1(n_577), .A2(n_702), .B1(n_705), .B2(n_706), .C1(n_707), .C2(n_708), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_579), .B(n_585), .Y(n_578) );
INVx1_ASAP7_75t_L g707 ( .A(n_579), .Y(n_707) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_581), .B(n_584), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_581), .B(n_607), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_581), .B(n_582), .Y(n_677) );
INVx1_ASAP7_75t_L g728 ( .A(n_581), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g658 ( .A(n_582), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g730 ( .A(n_582), .Y(n_730) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx2_ASAP7_75t_L g610 ( .A(n_583), .Y(n_610) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_584), .Y(n_653) );
AOI32xp33_ASAP7_75t_L g589 ( .A1(n_585), .A2(n_590), .A3(n_591), .B1(n_592), .B2(n_593), .Y(n_589) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_587), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g664 ( .A(n_587), .Y(n_664) );
OR2x2_ASAP7_75t_L g705 ( .A(n_587), .B(n_606), .Y(n_705) );
INVx1_ASAP7_75t_L g641 ( .A(n_588), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_590), .B(n_601), .Y(n_626) );
INVx3_ASAP7_75t_L g635 ( .A(n_590), .Y(n_635) );
AOI322xp5_ASAP7_75t_L g651 ( .A1(n_590), .A2(n_635), .A3(n_652), .B1(n_654), .B2(n_657), .C1(n_661), .C2(n_662), .Y(n_651) );
AND2x2_ASAP7_75t_L g627 ( .A(n_591), .B(n_628), .Y(n_627) );
INVxp67_ASAP7_75t_L g704 ( .A(n_591), .Y(n_704) );
A2O1A1O1Ixp25_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B(n_599), .C(n_607), .D(n_608), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_595), .B(n_638), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
OAI221xp5_ASAP7_75t_L g608 ( .A1(n_597), .A2(n_609), .B1(n_612), .B2(n_613), .C(n_616), .Y(n_608) );
INVx1_ASAP7_75t_SL g723 ( .A(n_597), .Y(n_723) );
AOI21xp33_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_604), .B(n_606), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
NAND2xp5_ASAP7_75t_SL g711 ( .A(n_601), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OAI221xp5_ASAP7_75t_SL g693 ( .A1(n_603), .A2(n_687), .B1(n_694), .B2(n_695), .C(n_696), .Y(n_693) );
OAI222xp33_ASAP7_75t_L g724 ( .A1(n_604), .A2(n_725), .B1(n_726), .B2(n_727), .C1(n_729), .C2(n_730), .Y(n_724) );
AND2x2_ASAP7_75t_L g682 ( .A(n_605), .B(n_668), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g694 ( .A1(n_605), .A2(n_620), .B(n_667), .Y(n_694) );
INVx1_ASAP7_75t_L g708 ( .A(n_605), .Y(n_708) );
INVx2_ASAP7_75t_SL g611 ( .A(n_606), .Y(n_611) );
AND2x2_ASAP7_75t_L g614 ( .A(n_607), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx1_ASAP7_75t_SL g648 ( .A(n_610), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_610), .B(n_620), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_611), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_611), .B(n_621), .Y(n_650) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OAI21xp5_ASAP7_75t_SL g616 ( .A1(n_617), .A2(n_619), .B(n_622), .Y(n_616) );
INVx1_ASAP7_75t_SL g634 ( .A(n_618), .Y(n_634) );
AND2x2_ASAP7_75t_L g681 ( .A(n_618), .B(n_664), .Y(n_681) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
AND2x2_ASAP7_75t_L g720 ( .A(n_620), .B(n_638), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_621), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g706 ( .A(n_622), .Y(n_706) );
AOI221xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_627), .B1(n_629), .B2(n_636), .C(n_639), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_632), .B1(n_634), .B2(n_635), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OAI22xp33_ASAP7_75t_L g639 ( .A1(n_633), .A2(n_640), .B1(n_642), .B2(n_644), .Y(n_639) );
OR2x2_ASAP7_75t_L g710 ( .A(n_634), .B(n_638), .Y(n_710) );
OR2x2_ASAP7_75t_L g713 ( .A(n_634), .B(n_648), .Y(n_713) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OAI221xp5_ASAP7_75t_L g709 ( .A1(n_655), .A2(n_710), .B1(n_711), .B2(n_713), .C(n_714), .Y(n_709) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVxp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND3xp33_ASAP7_75t_SL g665 ( .A(n_666), .B(n_680), .C(n_692), .Y(n_665) );
AOI222xp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_671), .B1(n_673), .B2(n_676), .C1(n_678), .C2(n_679), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_670), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_668), .B(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g690 ( .A(n_670), .Y(n_690) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVxp67_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_682), .B1(n_683), .B2(n_685), .C(n_688), .Y(n_680) );
INVx1_ASAP7_75t_L g695 ( .A(n_681), .Y(n_695) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
OAI21xp33_ASAP7_75t_L g714 ( .A1(n_685), .A2(n_715), .B(n_716), .Y(n_714) );
INVx1_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
NOR5xp2_ASAP7_75t_L g692 ( .A(n_693), .B(n_701), .C(n_709), .D(n_718), .E(n_724), .Y(n_692) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
OR2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
INVxp67_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
endmodule