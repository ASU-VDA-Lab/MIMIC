module fake_jpeg_1006_n_345 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_16),
.B(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_43),
.B(n_50),
.Y(n_101)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_22),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_46),
.B(n_48),
.Y(n_80)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_22),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_22),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_53),
.B(n_66),
.Y(n_103)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_16),
.B(n_13),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_56),
.B(n_64),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_21),
.B(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_75),
.Y(n_92)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_32),
.B(n_14),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_21),
.B(n_14),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_27),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_71),
.Y(n_113)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_28),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_32),
.B(n_12),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_74),
.B(n_11),
.Y(n_124)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_21),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_33),
.B1(n_19),
.B2(n_31),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_77),
.A2(n_111),
.B1(n_116),
.B2(n_88),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_52),
.A2(n_39),
.B1(n_24),
.B2(n_29),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_78),
.A2(n_104),
.B1(n_109),
.B2(n_110),
.Y(n_128)
);

INVx4_ASAP7_75t_SL g155 ( 
.A(n_88),
.Y(n_155)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_46),
.A2(n_29),
.B1(n_40),
.B2(n_34),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_60),
.B(n_66),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_119),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_71),
.A2(n_41),
.B1(n_75),
.B2(n_45),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_108),
.A2(n_70),
.B1(n_69),
.B2(n_54),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_48),
.A2(n_29),
.B1(n_40),
.B2(n_34),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_50),
.A2(n_37),
.B1(n_26),
.B2(n_30),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_47),
.A2(n_31),
.B1(n_19),
.B2(n_15),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_53),
.A2(n_37),
.B1(n_30),
.B2(n_20),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_112),
.A2(n_118),
.B1(n_120),
.B2(n_57),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_63),
.A2(n_20),
.B1(n_36),
.B2(n_35),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_115),
.A2(n_117),
.B1(n_9),
.B2(n_80),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_49),
.A2(n_35),
.B1(n_33),
.B2(n_15),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_55),
.A2(n_36),
.B1(n_20),
.B2(n_38),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_76),
.A2(n_36),
.B1(n_2),
.B2(n_3),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_44),
.B(n_1),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_65),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_73),
.B(n_13),
.C(n_12),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_6),
.C(n_8),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_51),
.B(n_13),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_124),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_125),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_113),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_126),
.B(n_129),
.Y(n_170)
);

AND2x2_ASAP7_75t_SL g127 ( 
.A(n_92),
.B(n_62),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_127),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_107),
.B(n_61),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_119),
.A2(n_59),
.B1(n_58),
.B2(n_72),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_131),
.A2(n_149),
.B1(n_151),
.B2(n_96),
.Y(n_173)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_105),
.B(n_101),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_133),
.B(n_153),
.Y(n_195)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_135),
.A2(n_141),
.B1(n_98),
.B2(n_81),
.Y(n_180)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_137),
.A2(n_156),
.B1(n_81),
.B2(n_114),
.Y(n_185)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_138),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_92),
.A2(n_67),
.B1(n_11),
.B2(n_5),
.Y(n_141)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_143),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_1),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_144),
.B(n_147),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_145),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_90),
.B(n_4),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_162),
.Y(n_182)
);

OA22x2_ASAP7_75t_L g148 ( 
.A1(n_108),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_148),
.A2(n_114),
.B(n_93),
.C(n_97),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_90),
.A2(n_9),
.B1(n_6),
.B2(n_8),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

INVxp33_ASAP7_75t_L g188 ( 
.A(n_150),
.Y(n_188)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_82),
.B(n_83),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_154),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_117),
.A2(n_82),
.B1(n_83),
.B2(n_89),
.Y(n_156)
);

BUFx12_ASAP7_75t_L g157 ( 
.A(n_89),
.Y(n_157)
);

INVx13_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_84),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_158),
.Y(n_192)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_91),
.Y(n_159)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_99),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_85),
.B(n_95),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_99),
.B(n_79),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_163),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_87),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_164),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_114),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_79),
.B(n_122),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_167),
.Y(n_183)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_94),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_128),
.A2(n_114),
.B(n_94),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_168),
.A2(n_184),
.B(n_201),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_148),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_127),
.A2(n_96),
.B1(n_97),
.B2(n_93),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_175),
.A2(n_180),
.B1(n_190),
.B2(n_202),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_155),
.A2(n_87),
.B1(n_95),
.B2(n_122),
.Y(n_176)
);

INVxp33_ASAP7_75t_SL g218 ( 
.A(n_176),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_184),
.Y(n_208)
);

OAI22x1_ASAP7_75t_L g217 ( 
.A1(n_185),
.A2(n_201),
.B1(n_125),
.B2(n_157),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_135),
.A2(n_141),
.B1(n_155),
.B2(n_151),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_189),
.A2(n_193),
.B1(n_139),
.B2(n_159),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_130),
.A2(n_127),
.B1(n_146),
.B2(n_126),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_130),
.B(n_154),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_147),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_138),
.A2(n_143),
.B1(n_148),
.B2(n_134),
.Y(n_193)
);

OAI22x1_ASAP7_75t_L g201 ( 
.A1(n_160),
.A2(n_139),
.B1(n_125),
.B2(n_136),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_205),
.A2(n_210),
.B1(n_211),
.B2(n_217),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_164),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_206),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_183),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_207),
.B(n_226),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_191),
.B(n_140),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_212),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_192),
.A2(n_148),
.B1(n_161),
.B2(n_152),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_192),
.A2(n_142),
.B1(n_145),
.B2(n_167),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_132),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_214),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_181),
.A2(n_150),
.B1(n_125),
.B2(n_157),
.Y(n_215)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_187),
.Y(n_216)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_216),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_219),
.A2(n_221),
.B(n_222),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_182),
.B(n_198),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_222),
.C(n_209),
.Y(n_247)
);

AO21x1_ASAP7_75t_L g221 ( 
.A1(n_179),
.A2(n_189),
.B(n_193),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_181),
.A2(n_199),
.B(n_195),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_223),
.Y(n_256)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_224),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_180),
.A2(n_182),
.B1(n_168),
.B2(n_199),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_227),
.Y(n_246)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_174),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_200),
.A2(n_183),
.B1(n_197),
.B2(n_175),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_188),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_228),
.B(n_229),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_170),
.B(n_172),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_174),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_231),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_196),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_235),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_178),
.A2(n_172),
.B(n_202),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_233),
.A2(n_206),
.B(n_223),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_178),
.B(n_203),
.Y(n_234)
);

BUFx24_ASAP7_75t_SL g262 ( 
.A(n_234),
.Y(n_262)
);

AND2x6_ASAP7_75t_L g235 ( 
.A(n_186),
.B(n_194),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_186),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_236),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_219),
.A2(n_194),
.B(n_177),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_241),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_231),
.A2(n_204),
.B1(n_169),
.B2(n_171),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_244),
.A2(n_208),
.B1(n_232),
.B2(n_217),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_230),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_259),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_247),
.B(n_206),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_204),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_254),
.C(n_255),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_212),
.B(n_169),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_207),
.B(n_203),
.C(n_171),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_213),
.B(n_171),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_221),
.A2(n_177),
.B(n_196),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_261),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_221),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_246),
.Y(n_273)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_264),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_275),
.C(n_281),
.Y(n_289)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_268),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_237),
.B(n_224),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_273),
.Y(n_291)
);

INVx8_ASAP7_75t_L g270 ( 
.A(n_262),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_270),
.A2(n_278),
.B1(n_280),
.B2(n_248),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_237),
.B(n_225),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_284),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_216),
.C(n_214),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_277),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_228),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_246),
.A2(n_250),
.B1(n_205),
.B2(n_248),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_245),
.B(n_210),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_279),
.Y(n_300)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_252),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_254),
.B(n_233),
.C(n_211),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_263),
.A2(n_205),
.B1(n_208),
.B2(n_218),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_282),
.A2(n_260),
.B1(n_243),
.B2(n_258),
.Y(n_287)
);

OAI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_283),
.A2(n_250),
.B1(n_241),
.B2(n_279),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_247),
.B(n_226),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_283),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_287),
.B(n_292),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_288),
.A2(n_297),
.B1(n_266),
.B2(n_244),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_282),
.A2(n_260),
.B1(n_252),
.B2(n_239),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_251),
.C(n_255),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_296),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_273),
.A2(n_239),
.B1(n_243),
.B2(n_244),
.Y(n_295)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_295),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_251),
.C(n_255),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_280),
.A2(n_250),
.B1(n_253),
.B2(n_259),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_267),
.B(n_265),
.C(n_275),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_299),
.B(n_281),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_290),
.B(n_274),
.Y(n_301)
);

MAJx2_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_304),
.C(n_306),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_303),
.B(n_308),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_253),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_287),
.A2(n_272),
.B(n_271),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_305),
.A2(n_307),
.B(n_310),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_272),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_293),
.A2(n_261),
.B(n_271),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_289),
.B(n_242),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_312),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_292),
.A2(n_242),
.B(n_266),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_313),
.A2(n_291),
.B(n_295),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_296),
.C(n_294),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_314),
.B(n_316),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_305),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_286),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_290),
.C(n_300),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_319),
.A2(n_323),
.B1(n_312),
.B2(n_240),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_297),
.C(n_286),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_302),
.C(n_309),
.Y(n_324)
);

FAx1_ASAP7_75t_SL g323 ( 
.A(n_301),
.B(n_235),
.CI(n_240),
.CON(n_323),
.SN(n_323)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_324),
.B(n_327),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_326),
.A2(n_328),
.B1(n_315),
.B2(n_320),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_304),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_270),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_329),
.B(n_330),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_319),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_322),
.A2(n_298),
.B(n_238),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_331),
.A2(n_318),
.B1(n_264),
.B2(n_238),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_332),
.A2(n_318),
.B1(n_331),
.B2(n_323),
.Y(n_338)
);

AOI221xp5_ASAP7_75t_L g339 ( 
.A1(n_334),
.A2(n_328),
.B1(n_336),
.B2(n_323),
.C(n_257),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_324),
.B(n_314),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_335),
.A2(n_325),
.B(n_327),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_337),
.B(n_338),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_339),
.A2(n_256),
.B1(n_257),
.B2(n_335),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_341),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_340),
.C(n_333),
.Y(n_343)
);

NAND2xp33_ASAP7_75t_SL g344 ( 
.A(n_343),
.B(n_333),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_321),
.B1(n_341),
.B2(n_340),
.Y(n_345)
);


endmodule