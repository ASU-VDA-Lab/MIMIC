module real_jpeg_26124_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_89;

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_2),
.B(n_49),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_2),
.B(n_41),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_2),
.B(n_64),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_2),
.B(n_28),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_2),
.B(n_46),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx8_ASAP7_75t_SL g47 ( 
.A(n_4),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_5),
.B(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_5),
.B(n_64),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_5),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_5),
.B(n_49),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_5),
.B(n_54),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_5),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_5),
.B(n_28),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_6),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_6),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_6),
.B(n_64),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_6),
.B(n_49),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_6),
.B(n_54),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_6),
.B(n_28),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_6),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_6),
.B(n_41),
.Y(n_234)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_8),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_8),
.B(n_41),
.Y(n_69)
);

INVxp33_ASAP7_75t_L g103 ( 
.A(n_8),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_8),
.B(n_34),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_8),
.B(n_64),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_8),
.B(n_28),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_8),
.B(n_54),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_8),
.B(n_192),
.Y(n_191)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_10),
.B(n_28),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_10),
.B(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_10),
.B(n_49),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_10),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_10),
.B(n_17),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_11),
.B(n_54),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_11),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_11),
.B(n_41),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_11),
.B(n_28),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_11),
.B(n_180),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_12),
.B(n_28),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_12),
.B(n_54),
.Y(n_92)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_13),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_13),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_13),
.B(n_64),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_15),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_16),
.B(n_34),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_16),
.B(n_46),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_16),
.B(n_49),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_16),
.B(n_54),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_16),
.B(n_64),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_16),
.B(n_28),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_16),
.B(n_17),
.Y(n_205)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_17),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_148),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_125),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_70),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_51),
.C(n_57),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_22),
.B(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.C(n_44),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_23),
.B(n_264),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_24),
.B(n_52),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_24),
.B(n_53),
.C(n_56),
.Y(n_114)
);

FAx1_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_30),
.CI(n_33),
.CON(n_24),
.SN(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_27),
.B(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_36),
.A2(n_37),
.B(n_40),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_36),
.B(n_44),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_39),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_48),
.C(n_50),
.Y(n_44)
);

FAx1_ASAP7_75t_SL g129 ( 
.A(n_45),
.B(n_48),
.CI(n_50),
.CON(n_129),
.SN(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_46),
.Y(n_76)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_51),
.B(n_57),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_54),
.Y(n_211)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_66),
.C(n_68),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_58),
.B(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_62),
.C(n_63),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_59),
.B(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_60),
.B(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_62),
.B(n_63),
.Y(n_253)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_66),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_93),
.B2(n_124),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_84),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_80),
.B1(n_82),
.B2(n_83),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_78),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_79),
.B(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_80),
.A2(n_82),
.B1(n_86),
.B2(n_113),
.Y(n_112)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_81),
.Y(n_180)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_81),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_86),
.C(n_87),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_89),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_86),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_88),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx24_ASAP7_75t_SL g270 ( 
.A(n_89),
.Y(n_270)
);

FAx1_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_91),
.CI(n_92),
.CON(n_89),
.SN(n_89)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

BUFx24_ASAP7_75t_SL g275 ( 
.A(n_93),
.Y(n_275)
);

FAx1_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_114),
.CI(n_115),
.CON(n_93),
.SN(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_104),
.C(n_110),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_95),
.B(n_145),
.Y(n_144)
);

BUFx24_ASAP7_75t_SL g271 ( 
.A(n_95),
.Y(n_271)
);

FAx1_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_99),
.CI(n_102),
.CON(n_95),
.SN(n_95)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_99),
.C(n_102),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_100),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_110),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.C(n_108),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_105),
.A2(n_106),
.B1(n_108),
.B2(n_109),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_123),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_119),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_144),
.C(n_146),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_126),
.A2(n_127),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_140),
.C(n_142),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_128),
.B(n_260),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.C(n_136),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_129),
.B(n_246),
.Y(n_245)
);

BUFx24_ASAP7_75t_SL g273 ( 
.A(n_129),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_130),
.A2(n_131),
.B1(n_136),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_136),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.C(n_139),
.Y(n_136)
);

FAx1_ASAP7_75t_SL g227 ( 
.A(n_137),
.B(n_138),
.CI(n_139),
.CON(n_227),
.SN(n_227)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_140),
.B(n_142),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_144),
.B(n_146),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_266),
.C(n_267),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_256),
.C(n_257),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_239),
.C(n_240),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_221),
.C(n_222),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_182),
.C(n_194),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_167),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_162),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_155),
.B(n_162),
.C(n_167),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_160),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_156),
.A2(n_157),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_185)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_163),
.B(n_165),
.C(n_166),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_174),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_168),
.B(n_175),
.C(n_176),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_169),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_181),
.Y(n_176)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_177),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_178),
.B(n_181),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.C(n_193),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_186),
.A2(n_187),
.B1(n_193),
.B2(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_198)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_217),
.C(n_218),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_203),
.C(n_208),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_201),
.C(n_202),
.Y(n_217)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.C(n_212),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_228),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_229),
.C(n_238),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_226),
.C(n_227),
.Y(n_243)
);

BUFx24_ASAP7_75t_SL g272 ( 
.A(n_227),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_238),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_236),
.B2(n_237),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_232),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_235),
.C(n_237),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_236),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_248),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_244),
.C(n_248),
.Y(n_256)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_252),
.C(n_254),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_251),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_252),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_261),
.B2(n_265),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_262),
.C(n_263),
.Y(n_266)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_261),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_268),
.Y(n_269)
);


endmodule