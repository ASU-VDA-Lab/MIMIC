module fake_netlist_1_2161_n_660 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_660);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_660;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx2_ASAP7_75t_SL g78 ( .A(n_34), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_29), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_74), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_4), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_18), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_45), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_61), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_20), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_22), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_9), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_21), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_59), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_7), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_54), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_20), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_11), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_38), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_0), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_8), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_35), .Y(n_97) );
INVxp67_ASAP7_75t_SL g98 ( .A(n_77), .Y(n_98) );
NOR2xp67_ASAP7_75t_L g99 ( .A(n_73), .B(n_6), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_23), .Y(n_100) );
INVx1_ASAP7_75t_SL g101 ( .A(n_50), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_68), .Y(n_102) );
INVxp67_ASAP7_75t_SL g103 ( .A(n_7), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_40), .Y(n_104) );
INVxp67_ASAP7_75t_SL g105 ( .A(n_30), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_26), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_47), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_44), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_56), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_24), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_27), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_31), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_39), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_43), .Y(n_114) );
INVxp67_ASAP7_75t_SL g115 ( .A(n_64), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_41), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_12), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_52), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_71), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_65), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_48), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_46), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_53), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_13), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_33), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_84), .Y(n_126) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_81), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_83), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_88), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_118), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_83), .Y(n_131) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_81), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_86), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_86), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_88), .Y(n_135) );
BUFx2_ASAP7_75t_L g136 ( .A(n_90), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_89), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_119), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_89), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_91), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_94), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_122), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_94), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_90), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_91), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_97), .Y(n_146) );
CKINVDCx16_ASAP7_75t_R g147 ( .A(n_78), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_97), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_114), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_114), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g151 ( .A(n_110), .Y(n_151) );
OA21x2_ASAP7_75t_L g152 ( .A1(n_116), .A2(n_28), .B(n_75), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_116), .Y(n_153) );
INVxp67_ASAP7_75t_L g154 ( .A(n_82), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_121), .Y(n_155) );
AND2x2_ASAP7_75t_L g156 ( .A(n_82), .B(n_0), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_85), .B(n_1), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_121), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_123), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_123), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_79), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_80), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_100), .Y(n_163) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_85), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_102), .Y(n_165) );
OAI21x1_ASAP7_75t_L g166 ( .A1(n_104), .A2(n_25), .B(n_72), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_106), .B(n_1), .Y(n_167) );
NOR2xp67_ASAP7_75t_L g168 ( .A(n_107), .B(n_2), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_129), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_127), .B(n_87), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_136), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_129), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_136), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_156), .Y(n_174) );
BUFx3_ASAP7_75t_L g175 ( .A(n_162), .Y(n_175) );
INVx4_ASAP7_75t_SL g176 ( .A(n_156), .Y(n_176) );
INVx1_ASAP7_75t_SL g177 ( .A(n_151), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_154), .B(n_125), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_156), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_129), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_154), .B(n_92), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_147), .B(n_125), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_129), .Y(n_183) );
BUFx3_ASAP7_75t_L g184 ( .A(n_162), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_150), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_147), .B(n_112), .Y(n_186) );
BUFx10_ASAP7_75t_L g187 ( .A(n_126), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_127), .B(n_124), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_130), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_129), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_150), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_161), .B(n_110), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_161), .B(n_111), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_150), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_150), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_129), .Y(n_196) );
AND2x4_ASAP7_75t_L g197 ( .A(n_132), .B(n_124), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_132), .B(n_87), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_139), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_163), .B(n_113), .Y(n_200) );
INVx2_ASAP7_75t_SL g201 ( .A(n_164), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_164), .B(n_117), .Y(n_202) );
BUFx4f_ASAP7_75t_L g203 ( .A(n_128), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_129), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_163), .B(n_109), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_139), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g207 ( .A1(n_165), .A2(n_95), .B1(n_117), .B2(n_96), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_135), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_139), .B(n_108), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_139), .Y(n_210) );
OAI221xp5_ASAP7_75t_L g211 ( .A1(n_157), .A2(n_92), .B1(n_95), .B2(n_96), .C(n_103), .Y(n_211) );
BUFx3_ASAP7_75t_L g212 ( .A(n_162), .Y(n_212) );
INVx1_ASAP7_75t_SL g213 ( .A(n_138), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_139), .Y(n_214) );
OR2x2_ASAP7_75t_SL g215 ( .A(n_157), .B(n_93), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_135), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_153), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_153), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_135), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_153), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_159), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_159), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_165), .B(n_101), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_128), .B(n_120), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_159), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_135), .Y(n_226) );
AND2x6_ASAP7_75t_L g227 ( .A(n_131), .B(n_78), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_131), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_133), .B(n_115), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_133), .B(n_99), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_183), .Y(n_231) );
NOR3xp33_ASAP7_75t_SL g232 ( .A(n_211), .B(n_142), .C(n_167), .Y(n_232) );
INVxp67_ASAP7_75t_SL g233 ( .A(n_201), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_183), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_178), .B(n_146), .Y(n_235) );
AOI22xp33_ASAP7_75t_SL g236 ( .A1(n_201), .A2(n_146), .B1(n_134), .B2(n_145), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_171), .B(n_145), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_192), .B(n_148), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_227), .Y(n_239) );
INVxp67_ASAP7_75t_L g240 ( .A(n_177), .Y(n_240) );
BUFx4f_ASAP7_75t_L g241 ( .A(n_227), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_181), .B(n_148), .Y(n_242) );
INVx4_ASAP7_75t_L g243 ( .A(n_176), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_189), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_199), .Y(n_245) );
INVx6_ASAP7_75t_L g246 ( .A(n_176), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_176), .Y(n_247) );
INVx3_ASAP7_75t_L g248 ( .A(n_227), .Y(n_248) );
INVx4_ASAP7_75t_L g249 ( .A(n_227), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_170), .Y(n_250) );
BUFx2_ASAP7_75t_L g251 ( .A(n_170), .Y(n_251) );
AND2x4_ASAP7_75t_L g252 ( .A(n_170), .B(n_168), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_188), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_181), .B(n_160), .Y(n_254) );
INVx3_ASAP7_75t_L g255 ( .A(n_227), .Y(n_255) );
INVx2_ASAP7_75t_SL g256 ( .A(n_188), .Y(n_256) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_188), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_227), .Y(n_258) );
INVx3_ASAP7_75t_L g259 ( .A(n_217), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_206), .Y(n_260) );
O2A1O1Ixp5_ASAP7_75t_L g261 ( .A1(n_203), .A2(n_167), .B(n_155), .C(n_140), .Y(n_261) );
NOR2xp33_ASAP7_75t_R g262 ( .A(n_189), .B(n_134), .Y(n_262) );
INVx4_ASAP7_75t_L g263 ( .A(n_203), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_210), .Y(n_264) );
BUFx2_ASAP7_75t_L g265 ( .A(n_197), .Y(n_265) );
INVx5_ASAP7_75t_L g266 ( .A(n_183), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_203), .B(n_140), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_214), .Y(n_268) );
INVx1_ASAP7_75t_SL g269 ( .A(n_213), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_197), .B(n_149), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_197), .Y(n_271) );
NOR2xp33_ASAP7_75t_R g272 ( .A(n_187), .B(n_137), .Y(n_272) );
AND2x4_ASAP7_75t_L g273 ( .A(n_198), .B(n_168), .Y(n_273) );
AND2x2_ASAP7_75t_SL g274 ( .A(n_198), .B(n_152), .Y(n_274) );
OAI21xp5_ASAP7_75t_L g275 ( .A1(n_185), .A2(n_166), .B(n_152), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_218), .Y(n_276) );
INVx3_ASAP7_75t_L g277 ( .A(n_220), .Y(n_277) );
BUFx3_ASAP7_75t_L g278 ( .A(n_198), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_191), .Y(n_279) );
INVx5_ASAP7_75t_L g280 ( .A(n_183), .Y(n_280) );
O2A1O1Ixp33_ASAP7_75t_L g281 ( .A1(n_173), .A2(n_155), .B(n_137), .C(n_160), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_194), .Y(n_282) );
AND2x4_ASAP7_75t_L g283 ( .A(n_174), .B(n_158), .Y(n_283) );
BUFx6f_ASAP7_75t_L g284 ( .A(n_204), .Y(n_284) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_204), .Y(n_285) );
NOR3xp33_ASAP7_75t_SL g286 ( .A(n_186), .B(n_149), .C(n_158), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_186), .A2(n_179), .B1(n_202), .B2(n_182), .Y(n_287) );
AND2x4_ASAP7_75t_L g288 ( .A(n_224), .B(n_144), .Y(n_288) );
AOI211xp5_ASAP7_75t_L g289 ( .A1(n_224), .A2(n_144), .B(n_141), .C(n_143), .Y(n_289) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_223), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_195), .Y(n_291) );
INVx2_ASAP7_75t_SL g292 ( .A(n_228), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_229), .B(n_144), .Y(n_293) );
NOR2xp33_ASAP7_75t_R g294 ( .A(n_187), .B(n_144), .Y(n_294) );
NOR3xp33_ASAP7_75t_SL g295 ( .A(n_230), .B(n_98), .C(n_105), .Y(n_295) );
CKINVDCx16_ASAP7_75t_R g296 ( .A(n_187), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_296), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_259), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_292), .A2(n_209), .B(n_152), .Y(n_299) );
INVx3_ASAP7_75t_SL g300 ( .A(n_269), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_290), .B(n_229), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_272), .Y(n_302) );
AND2x4_ASAP7_75t_L g303 ( .A(n_278), .B(n_205), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_278), .B(n_205), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_257), .Y(n_305) );
INVx4_ASAP7_75t_L g306 ( .A(n_243), .Y(n_306) );
AND2x4_ASAP7_75t_L g307 ( .A(n_250), .B(n_200), .Y(n_307) );
INVx4_ASAP7_75t_L g308 ( .A(n_243), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_251), .Y(n_309) );
AOI221xp5_ASAP7_75t_L g310 ( .A1(n_237), .A2(n_200), .B1(n_193), .B2(n_207), .C(n_230), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_256), .B(n_193), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_259), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_251), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_262), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_243), .Y(n_315) );
INVx2_ASAP7_75t_SL g316 ( .A(n_294), .Y(n_316) );
INVx4_ASAP7_75t_L g317 ( .A(n_246), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_292), .A2(n_209), .B(n_152), .Y(n_318) );
INVx8_ASAP7_75t_L g319 ( .A(n_283), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_265), .B(n_222), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_256), .B(n_221), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_270), .B(n_225), .Y(n_322) );
BUFx3_ASAP7_75t_L g323 ( .A(n_246), .Y(n_323) );
AOI22xp5_ASAP7_75t_L g324 ( .A1(n_265), .A2(n_215), .B1(n_141), .B2(n_143), .Y(n_324) );
INVx5_ASAP7_75t_L g325 ( .A(n_246), .Y(n_325) );
OAI21xp33_ASAP7_75t_L g326 ( .A1(n_236), .A2(n_184), .B(n_212), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_253), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_259), .Y(n_328) );
NOR2x1_ASAP7_75t_SL g329 ( .A(n_249), .B(n_141), .Y(n_329) );
INVx3_ASAP7_75t_L g330 ( .A(n_246), .Y(n_330) );
INVxp67_ASAP7_75t_SL g331 ( .A(n_240), .Y(n_331) );
AND2x4_ASAP7_75t_L g332 ( .A(n_271), .B(n_166), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_249), .Y(n_333) );
CKINVDCx11_ASAP7_75t_R g334 ( .A(n_252), .Y(n_334) );
INVx2_ASAP7_75t_SL g335 ( .A(n_276), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_242), .B(n_143), .Y(n_336) );
CKINVDCx6p67_ASAP7_75t_R g337 ( .A(n_252), .Y(n_337) );
OR2x6_ASAP7_75t_L g338 ( .A(n_252), .B(n_166), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_244), .B(n_2), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_254), .B(n_162), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_287), .B(n_3), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_276), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_273), .B(n_162), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_233), .B(n_162), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_283), .B(n_162), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_283), .Y(n_346) );
OAI21xp33_ASAP7_75t_SL g347 ( .A1(n_235), .A2(n_190), .B(n_169), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_319), .A2(n_273), .B1(n_288), .B2(n_293), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_319), .A2(n_276), .B1(n_277), .B2(n_286), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_327), .Y(n_350) );
CKINVDCx16_ASAP7_75t_R g351 ( .A(n_300), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_319), .B(n_273), .Y(n_352) );
OAI211xp5_ASAP7_75t_L g353 ( .A1(n_310), .A2(n_232), .B(n_289), .C(n_281), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_319), .A2(n_288), .B1(n_293), .B2(n_267), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_300), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_322), .A2(n_277), .B1(n_263), .B2(n_238), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_341), .B(n_277), .Y(n_357) );
OAI22xp33_ASAP7_75t_L g358 ( .A1(n_314), .A2(n_244), .B1(n_249), .B2(n_241), .Y(n_358) );
OAI22xp5_ASAP7_75t_SL g359 ( .A1(n_314), .A2(n_274), .B1(n_288), .B2(n_247), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_301), .B(n_295), .Y(n_360) );
INVx4_ASAP7_75t_SL g361 ( .A(n_333), .Y(n_361) );
OAI22xp33_ASAP7_75t_L g362 ( .A1(n_302), .A2(n_241), .B1(n_263), .B2(n_258), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_298), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_346), .B(n_282), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_305), .Y(n_365) );
OR2x4_ASAP7_75t_L g366 ( .A(n_339), .B(n_258), .Y(n_366) );
AOI221xp5_ASAP7_75t_L g367 ( .A1(n_307), .A2(n_279), .B1(n_261), .B2(n_267), .C(n_291), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_309), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_313), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_331), .B(n_282), .Y(n_370) );
INVx4_ASAP7_75t_L g371 ( .A(n_306), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_297), .Y(n_372) );
AOI21xp33_ASAP7_75t_SL g373 ( .A1(n_297), .A2(n_3), .B(n_4), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_298), .Y(n_374) );
NAND2x1_ASAP7_75t_L g375 ( .A(n_335), .B(n_239), .Y(n_375) );
AND2x4_ASAP7_75t_SL g376 ( .A(n_337), .B(n_263), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_336), .Y(n_377) );
AOI32xp33_ASAP7_75t_L g378 ( .A1(n_302), .A2(n_291), .A3(n_268), .B1(n_264), .B2(n_260), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_312), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_357), .A2(n_334), .B1(n_307), .B2(n_303), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_377), .B(n_320), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_350), .Y(n_382) );
OAI222xp33_ASAP7_75t_L g383 ( .A1(n_378), .A2(n_338), .B1(n_324), .B2(n_316), .C1(n_311), .C2(n_335), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_357), .B(n_312), .Y(n_384) );
BUFx2_ASAP7_75t_L g385 ( .A(n_355), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_370), .B(n_328), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_350), .B(n_307), .Y(n_387) );
AOI221xp5_ASAP7_75t_L g388 ( .A1(n_353), .A2(n_303), .B1(n_304), .B2(n_343), .C(n_340), .Y(n_388) );
AO31x2_ASAP7_75t_L g389 ( .A1(n_349), .A2(n_343), .A3(n_299), .B(n_318), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_370), .B(n_328), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_364), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_364), .B(n_303), .Y(n_392) );
AOI211xp5_ASAP7_75t_L g393 ( .A1(n_373), .A2(n_326), .B(n_304), .C(n_347), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g394 ( .A(n_351), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_363), .Y(n_395) );
BUFx3_ASAP7_75t_L g396 ( .A(n_371), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_366), .A2(n_337), .B1(n_338), .B2(n_321), .Y(n_397) );
BUFx2_ASAP7_75t_L g398 ( .A(n_355), .Y(n_398) );
BUFx12f_ASAP7_75t_L g399 ( .A(n_372), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_359), .A2(n_334), .B1(n_304), .B2(n_345), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_363), .B(n_342), .Y(n_401) );
INVx4_ASAP7_75t_L g402 ( .A(n_361), .Y(n_402) );
OAI211xp5_ASAP7_75t_L g403 ( .A1(n_348), .A2(n_344), .B(n_342), .C(n_306), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_368), .A2(n_274), .B1(n_338), .B2(n_332), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_374), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_360), .B(n_306), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_374), .Y(n_407) );
OAI211xp5_ASAP7_75t_SL g408 ( .A1(n_380), .A2(n_365), .B(n_369), .C(n_352), .Y(n_408) );
OAI222xp33_ASAP7_75t_L g409 ( .A1(n_400), .A2(n_371), .B1(n_372), .B2(n_358), .C1(n_356), .C2(n_366), .Y(n_409) );
OAI22xp33_ASAP7_75t_L g410 ( .A1(n_385), .A2(n_366), .B1(n_371), .B2(n_379), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_381), .B(n_354), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_395), .Y(n_412) );
BUFx2_ASAP7_75t_L g413 ( .A(n_385), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_385), .B(n_379), .Y(n_414) );
BUFx2_ASAP7_75t_L g415 ( .A(n_398), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_381), .B(n_376), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_394), .Y(n_417) );
AOI22xp33_ASAP7_75t_SL g418 ( .A1(n_398), .A2(n_376), .B1(n_329), .B2(n_308), .Y(n_418) );
CKINVDCx20_ASAP7_75t_R g419 ( .A(n_394), .Y(n_419) );
OAI221xp5_ASAP7_75t_L g420 ( .A1(n_380), .A2(n_367), .B1(n_315), .B2(n_375), .C(n_275), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_381), .B(n_332), .Y(n_421) );
OAI211xp5_ASAP7_75t_L g422 ( .A1(n_400), .A2(n_152), .B(n_135), .C(n_375), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_398), .B(n_332), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_382), .Y(n_424) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_402), .Y(n_425) );
OAI211xp5_ASAP7_75t_SL g426 ( .A1(n_393), .A2(n_169), .B(n_219), .C(n_208), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_382), .B(n_308), .Y(n_427) );
OAI211xp5_ASAP7_75t_SL g428 ( .A1(n_393), .A2(n_180), .B(n_172), .C(n_190), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_386), .B(n_390), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_395), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_386), .B(n_361), .Y(n_431) );
AOI221xp5_ASAP7_75t_L g432 ( .A1(n_387), .A2(n_135), .B1(n_264), .B2(n_268), .C(n_260), .Y(n_432) );
INVx3_ASAP7_75t_L g433 ( .A(n_402), .Y(n_433) );
NAND2xp33_ASAP7_75t_R g434 ( .A(n_406), .B(n_5), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_399), .B(n_308), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_386), .Y(n_436) );
A2O1A1Ixp33_ASAP7_75t_L g437 ( .A1(n_388), .A2(n_241), .B(n_315), .C(n_239), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_395), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_388), .A2(n_315), .B1(n_362), .B2(n_333), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_390), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_390), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_429), .B(n_405), .Y(n_442) );
OAI31xp33_ASAP7_75t_L g443 ( .A1(n_408), .A2(n_383), .A3(n_397), .B(n_406), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_429), .B(n_405), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_424), .Y(n_445) );
OAI22xp5_ASAP7_75t_SL g446 ( .A1(n_419), .A2(n_399), .B1(n_396), .B2(n_402), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_436), .B(n_391), .Y(n_447) );
AND2x4_ASAP7_75t_L g448 ( .A(n_433), .B(n_402), .Y(n_448) );
INVx2_ASAP7_75t_SL g449 ( .A(n_414), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_412), .Y(n_450) );
INVx2_ASAP7_75t_SL g451 ( .A(n_414), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_440), .B(n_405), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_441), .B(n_392), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_434), .A2(n_387), .B1(n_392), .B2(n_403), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_413), .Y(n_455) );
AND2x4_ASAP7_75t_L g456 ( .A(n_433), .B(n_402), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_412), .Y(n_457) );
AOI221xp5_ASAP7_75t_L g458 ( .A1(n_411), .A2(n_383), .B1(n_391), .B2(n_384), .C(n_404), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_427), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_430), .B(n_407), .Y(n_460) );
OAI33xp33_ASAP7_75t_L g461 ( .A1(n_417), .A2(n_5), .A3(n_6), .B1(n_8), .B2(n_9), .B3(n_10), .Y(n_461) );
INVx4_ASAP7_75t_L g462 ( .A(n_433), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_413), .B(n_407), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_421), .B(n_384), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_427), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_430), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_415), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_415), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_438), .B(n_407), .Y(n_469) );
AOI221xp5_ASAP7_75t_L g470 ( .A1(n_409), .A2(n_384), .B1(n_404), .B2(n_135), .C(n_403), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_425), .Y(n_471) );
NOR2xp33_ASAP7_75t_SL g472 ( .A(n_417), .B(n_399), .Y(n_472) );
OAI33xp33_ASAP7_75t_L g473 ( .A1(n_410), .A2(n_10), .A3(n_11), .B1(n_12), .B2(n_13), .B3(n_14), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_431), .B(n_423), .Y(n_474) );
NOR3xp33_ASAP7_75t_L g475 ( .A(n_426), .B(n_396), .C(n_330), .Y(n_475) );
AOI222xp33_ASAP7_75t_L g476 ( .A1(n_416), .A2(n_419), .B1(n_435), .B2(n_431), .C1(n_396), .C2(n_439), .Y(n_476) );
INVx1_ASAP7_75t_SL g477 ( .A(n_423), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_418), .Y(n_478) );
INVx3_ASAP7_75t_L g479 ( .A(n_425), .Y(n_479) );
NOR3xp33_ASAP7_75t_L g480 ( .A(n_428), .B(n_330), .C(n_401), .Y(n_480) );
INVx2_ASAP7_75t_SL g481 ( .A(n_425), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_420), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_437), .B(n_401), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_425), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_432), .B(n_389), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_425), .B(n_389), .Y(n_486) );
AOI211xp5_ASAP7_75t_L g487 ( .A1(n_422), .A2(n_226), .B(n_204), .C(n_216), .Y(n_487) );
OAI31xp33_ASAP7_75t_L g488 ( .A1(n_408), .A2(n_255), .A3(n_248), .B(n_239), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_486), .B(n_389), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_442), .B(n_389), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_445), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_486), .B(n_389), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_442), .B(n_389), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_444), .B(n_389), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_444), .B(n_389), .Y(n_495) );
INVxp67_ASAP7_75t_L g496 ( .A(n_472), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_474), .B(n_14), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_449), .B(n_15), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_459), .Y(n_499) );
NOR3xp33_ASAP7_75t_L g500 ( .A(n_461), .B(n_196), .C(n_330), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_478), .B(n_15), .Y(n_501) );
NOR3xp33_ASAP7_75t_L g502 ( .A(n_473), .B(n_317), .C(n_248), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_446), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_465), .B(n_449), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_451), .B(n_16), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_467), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_451), .B(n_16), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_468), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_477), .B(n_17), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_474), .B(n_450), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_455), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_452), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_450), .B(n_457), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_463), .B(n_17), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_452), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_463), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_457), .B(n_18), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_466), .B(n_19), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_466), .B(n_19), .Y(n_519) );
INVx1_ASAP7_75t_SL g520 ( .A(n_460), .Y(n_520) );
NOR2xp33_ASAP7_75t_SL g521 ( .A(n_462), .B(n_317), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_460), .B(n_361), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_447), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_469), .B(n_361), .Y(n_524) );
INVx2_ASAP7_75t_SL g525 ( .A(n_462), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_469), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_471), .B(n_204), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_453), .B(n_245), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_462), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_471), .B(n_216), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_464), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_481), .B(n_32), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_484), .Y(n_533) );
CKINVDCx16_ASAP7_75t_R g534 ( .A(n_448), .Y(n_534) );
AND2x2_ASAP7_75t_SL g535 ( .A(n_448), .B(n_333), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_476), .A2(n_245), .B1(n_226), .B2(n_216), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_448), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_482), .B(n_216), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_481), .B(n_36), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_458), .B(n_226), .Y(n_540) );
NOR2x1_ASAP7_75t_L g541 ( .A(n_456), .B(n_317), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_479), .B(n_37), .Y(n_542) );
O2A1O1Ixp33_ASAP7_75t_SL g543 ( .A1(n_496), .A2(n_470), .B(n_454), .C(n_487), .Y(n_543) );
O2A1O1Ixp33_ASAP7_75t_SL g544 ( .A1(n_525), .A2(n_485), .B(n_483), .C(n_443), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_531), .B(n_456), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_536), .A2(n_475), .B1(n_480), .B2(n_456), .Y(n_546) );
AOI21xp33_ASAP7_75t_SL g547 ( .A1(n_503), .A2(n_488), .B(n_479), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_536), .A2(n_479), .B1(n_325), .B2(n_323), .Y(n_548) );
OAI22xp33_ASAP7_75t_L g549 ( .A1(n_534), .A2(n_503), .B1(n_525), .B2(n_521), .Y(n_549) );
INVx3_ASAP7_75t_SL g550 ( .A(n_535), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_510), .B(n_226), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_501), .A2(n_255), .B1(n_248), .B2(n_323), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_491), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_497), .A2(n_325), .B1(n_333), .B2(n_258), .Y(n_554) );
OAI22xp33_ASAP7_75t_L g555 ( .A1(n_498), .A2(n_325), .B1(n_258), .B2(n_255), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_523), .B(n_42), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_501), .B(n_49), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_499), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_511), .Y(n_559) );
OAI221xp5_ASAP7_75t_SL g560 ( .A1(n_497), .A2(n_212), .B1(n_184), .B2(n_175), .C(n_58), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_506), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_520), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_510), .B(n_51), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_508), .Y(n_564) );
NAND3xp33_ASAP7_75t_L g565 ( .A(n_509), .B(n_175), .C(n_325), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_513), .Y(n_566) );
AOI222xp33_ASAP7_75t_L g567 ( .A1(n_494), .A2(n_55), .B1(n_57), .B2(n_60), .C1(n_62), .C2(n_63), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_504), .Y(n_568) );
AOI221xp5_ASAP7_75t_L g569 ( .A1(n_505), .A2(n_231), .B1(n_234), .B2(n_285), .C(n_284), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_507), .B(n_66), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_537), .B(n_67), .Y(n_571) );
OAI221xp5_ASAP7_75t_L g572 ( .A1(n_514), .A2(n_280), .B1(n_266), .B2(n_285), .C(n_231), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_526), .B(n_69), .Y(n_573) );
OAI21xp5_ASAP7_75t_L g574 ( .A1(n_517), .A2(n_266), .B(n_280), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_489), .A2(n_285), .B1(n_231), .B2(n_234), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_512), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_535), .A2(n_266), .B1(n_280), .B2(n_70), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_529), .A2(n_266), .B1(n_280), .B2(n_76), .Y(n_578) );
OAI211xp5_ASAP7_75t_L g579 ( .A1(n_490), .A2(n_266), .B(n_280), .C(n_231), .Y(n_579) );
AOI21xp33_ASAP7_75t_SL g580 ( .A1(n_517), .A2(n_231), .B(n_234), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_522), .A2(n_234), .B1(n_285), .B2(n_284), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_528), .A2(n_234), .B1(n_285), .B2(n_284), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_515), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_533), .Y(n_584) );
OAI22xp33_ASAP7_75t_SL g585 ( .A1(n_519), .A2(n_284), .B1(n_516), .B2(n_542), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_493), .B(n_495), .Y(n_586) );
AOI33xp33_ASAP7_75t_L g587 ( .A1(n_489), .A2(n_492), .A3(n_494), .B1(n_518), .B2(n_513), .B3(n_524), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_492), .B(n_518), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_538), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_553), .Y(n_590) );
BUFx2_ASAP7_75t_SL g591 ( .A(n_571), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_566), .B(n_527), .Y(n_592) );
OAI21xp33_ASAP7_75t_SL g593 ( .A1(n_587), .A2(n_541), .B(n_532), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_586), .B(n_527), .Y(n_594) );
INVx3_ASAP7_75t_L g595 ( .A(n_550), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_584), .Y(n_596) );
OAI211xp5_ASAP7_75t_SL g597 ( .A1(n_567), .A2(n_540), .B(n_500), .C(n_539), .Y(n_597) );
OAI21xp5_ASAP7_75t_L g598 ( .A1(n_567), .A2(n_502), .B(n_530), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_561), .Y(n_599) );
NOR3xp33_ASAP7_75t_L g600 ( .A(n_565), .B(n_549), .C(n_547), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_564), .Y(n_601) );
OAI21xp33_ASAP7_75t_L g602 ( .A1(n_568), .A2(n_588), .B(n_562), .Y(n_602) );
AOI321xp33_ASAP7_75t_R g603 ( .A1(n_544), .A2(n_559), .A3(n_583), .B1(n_576), .B2(n_558), .C(n_545), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_589), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_551), .B(n_554), .Y(n_605) );
INVxp67_ASAP7_75t_L g606 ( .A(n_563), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_585), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_571), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_579), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_574), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_546), .B(n_574), .Y(n_611) );
INVx1_ASAP7_75t_SL g612 ( .A(n_573), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_556), .Y(n_613) );
BUFx3_ASAP7_75t_L g614 ( .A(n_581), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_580), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_554), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_582), .Y(n_617) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_565), .B(n_548), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_575), .B(n_569), .Y(n_619) );
INVxp67_ASAP7_75t_L g620 ( .A(n_570), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_543), .B(n_555), .Y(n_621) );
NOR3x1_ASAP7_75t_L g622 ( .A(n_603), .B(n_577), .C(n_572), .Y(n_622) );
XNOR2xp5_ASAP7_75t_L g623 ( .A(n_595), .B(n_552), .Y(n_623) );
INVx2_ASAP7_75t_SL g624 ( .A(n_595), .Y(n_624) );
XNOR2xp5_ASAP7_75t_L g625 ( .A(n_595), .B(n_578), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_611), .B(n_557), .Y(n_626) );
XNOR2xp5_ASAP7_75t_L g627 ( .A(n_594), .B(n_560), .Y(n_627) );
OAI22xp33_ASAP7_75t_SL g628 ( .A1(n_607), .A2(n_609), .B1(n_618), .B2(n_621), .Y(n_628) );
INVxp67_ASAP7_75t_L g629 ( .A(n_614), .Y(n_629) );
CKINVDCx20_ASAP7_75t_R g630 ( .A(n_606), .Y(n_630) );
OAI21xp5_ASAP7_75t_L g631 ( .A1(n_593), .A2(n_600), .B(n_609), .Y(n_631) );
NAND4xp25_ASAP7_75t_L g632 ( .A(n_598), .B(n_597), .C(n_614), .D(n_618), .Y(n_632) );
INVx3_ASAP7_75t_L g633 ( .A(n_608), .Y(n_633) );
AOI21xp33_ASAP7_75t_L g634 ( .A1(n_615), .A2(n_610), .B(n_620), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_602), .B(n_604), .Y(n_635) );
OAI21xp5_ASAP7_75t_SL g636 ( .A1(n_619), .A2(n_612), .B(n_616), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_596), .Y(n_637) );
INVx1_ASAP7_75t_SL g638 ( .A(n_624), .Y(n_638) );
INVx1_ASAP7_75t_SL g639 ( .A(n_630), .Y(n_639) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_629), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_632), .A2(n_590), .B1(n_601), .B2(n_599), .C(n_613), .Y(n_641) );
AOI221xp5_ASAP7_75t_L g642 ( .A1(n_628), .A2(n_619), .B1(n_617), .B2(n_591), .C(n_592), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_626), .A2(n_605), .B1(n_627), .B2(n_634), .Y(n_643) );
OAI211xp5_ASAP7_75t_SL g644 ( .A1(n_636), .A2(n_605), .B(n_626), .C(n_635), .Y(n_644) );
NAND3xp33_ASAP7_75t_L g645 ( .A(n_635), .B(n_625), .C(n_623), .Y(n_645) );
NAND3xp33_ASAP7_75t_SL g646 ( .A(n_630), .B(n_622), .C(n_637), .Y(n_646) );
OAI211xp5_ASAP7_75t_SL g647 ( .A1(n_633), .A2(n_631), .B(n_629), .C(n_636), .Y(n_647) );
A2O1A1Ixp33_ASAP7_75t_L g648 ( .A1(n_631), .A2(n_632), .B(n_636), .C(n_603), .Y(n_648) );
NOR2x1_ASAP7_75t_L g649 ( .A(n_632), .B(n_631), .Y(n_649) );
CKINVDCx5p33_ASAP7_75t_R g650 ( .A(n_639), .Y(n_650) );
BUFx2_ASAP7_75t_L g651 ( .A(n_640), .Y(n_651) );
OAI21x1_ASAP7_75t_SL g652 ( .A1(n_642), .A2(n_649), .B(n_641), .Y(n_652) );
NAND3xp33_ASAP7_75t_L g653 ( .A(n_651), .B(n_648), .C(n_647), .Y(n_653) );
OR3x1_ASAP7_75t_L g654 ( .A(n_652), .B(n_646), .C(n_644), .Y(n_654) );
OAI21xp5_ASAP7_75t_L g655 ( .A1(n_651), .A2(n_643), .B(n_645), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_655), .B(n_650), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_653), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_656), .Y(n_658) );
AOI22xp5_ASAP7_75t_SL g659 ( .A1(n_658), .A2(n_650), .B1(n_657), .B2(n_654), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_659), .A2(n_643), .B(n_638), .Y(n_660) );
endmodule