module real_jpeg_17553_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_525;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVxp33_ASAP7_75t_L g529 ( 
.A(n_0),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_1),
.A2(n_19),
.B(n_528),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_1),
.B(n_529),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_2),
.B(n_40),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_2),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_2),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_2),
.B(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_2),
.B(n_155),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_2),
.B(n_195),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_2),
.B(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_3),
.Y(n_82)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_3),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_3),
.Y(n_299)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_4),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_4),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_4),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_4),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_5),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_5),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_5),
.B(n_265),
.Y(n_264)
);

AND2x2_ASAP7_75t_SL g277 ( 
.A(n_5),
.B(n_278),
.Y(n_277)
);

AND2x2_ASAP7_75t_SL g300 ( 
.A(n_5),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_5),
.B(n_432),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_5),
.B(n_437),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_5),
.B(n_295),
.Y(n_459)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_6),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_6),
.B(n_231),
.Y(n_230)
);

AND2x2_ASAP7_75t_SL g298 ( 
.A(n_6),
.B(n_299),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_6),
.A2(n_11),
.B1(n_313),
.B2(n_315),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_6),
.B(n_451),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_6),
.B(n_462),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_6),
.B(n_493),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_7),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_7),
.B(n_341),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_7),
.B(n_385),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_7),
.B(n_446),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_7),
.B(n_455),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_7),
.B(n_502),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_7),
.B(n_507),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_8),
.B(n_28),
.Y(n_27)
);

NAND2x1p5_ASAP7_75t_L g35 ( 
.A(n_8),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_8),
.B(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_8),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_8),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_8),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_8),
.B(n_169),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_8),
.B(n_66),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_9),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g248 ( 
.A(n_9),
.Y(n_248)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_9),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_9),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_10),
.Y(n_130)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_10),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_10),
.Y(n_205)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_10),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_10),
.Y(n_383)
);

NAND2x1_ASAP7_75t_SL g54 ( 
.A(n_11),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_11),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_11),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_11),
.B(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_11),
.B(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_11),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_11),
.B(n_101),
.Y(n_250)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_11),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_12),
.Y(n_88)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_12),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_12),
.Y(n_289)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_13),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_13),
.B(n_127),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_13),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_13),
.B(n_268),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_13),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_13),
.B(n_294),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_14),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_15),
.B(n_66),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_15),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_15),
.B(n_338),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_15),
.B(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_15),
.B(n_454),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_15),
.B(n_155),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_15),
.B(n_489),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_15),
.B(n_493),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_16),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g197 ( 
.A(n_16),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_17),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_109),
.Y(n_19)
);

NAND2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_108),
.Y(n_20)
);

INVxp33_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_67),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_23),
.B(n_67),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_50),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_38),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_31),
.C(n_34),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_26),
.A2(n_27),
.B1(n_34),
.B2(n_35),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_26),
.A2(n_27),
.B1(n_57),
.B2(n_58),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_26),
.B(n_159),
.C(n_230),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_26),
.A2(n_27),
.B1(n_230),
.B2(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_27),
.B(n_57),
.C(n_61),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_30),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_SL g51 ( 
.A(n_31),
.B(n_52),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_31),
.B(n_123),
.C(n_128),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_31),
.B(n_158),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_35),
.B1(n_44),
.B2(n_47),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_34),
.B(n_241),
.C(n_249),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_34),
.A2(n_35),
.B1(n_249),
.B2(n_250),
.Y(n_358)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_37),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_43),
.B1(n_48),
.B2(n_49),
.Y(n_38)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_74),
.C(n_80),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_39),
.A2(n_48),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_44),
.B(n_133),
.C(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_44),
.B(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_53),
.C(n_56),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g69 ( 
.A(n_51),
.B(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_57),
.A2(n_58),
.B1(n_99),
.B2(n_100),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_57),
.A2(n_58),
.B1(n_153),
.B2(n_154),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_99),
.C(n_102),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_58),
.B(n_154),
.C(n_273),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_63),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_63),
.B(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_66),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_72),
.C(n_93),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_68),
.A2(n_69),
.B1(n_72),
.B2(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_83),
.C(n_89),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_73),
.B(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_74),
.A2(n_75),
.B1(n_80),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g265 ( 
.A(n_79),
.Y(n_265)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_79),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_79),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_79),
.Y(n_387)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_80),
.Y(n_163)
);

MAJx2_ASAP7_75t_L g201 ( 
.A(n_80),
.B(n_202),
.C(n_206),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_80),
.B(n_206),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_82),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_89),
.B1(n_90),
.B2(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

MAJx2_ASAP7_75t_L g200 ( 
.A(n_89),
.B(n_201),
.C(n_208),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_89),
.A2(n_90),
.B1(n_208),
.B2(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_90),
.B(n_165),
.C(n_170),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_90),
.B(n_171),
.Y(n_213)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_98),
.C(n_106),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_94),
.A2(n_95),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_106),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_99),
.A2(n_100),
.B1(n_132),
.B2(n_133),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_99),
.A2(n_100),
.B1(n_298),
.B2(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_132),
.C(n_137),
.Y(n_131)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_100),
.B(n_298),
.C(n_300),
.Y(n_297)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_101),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_101),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_121),
.Y(n_120)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_105),
.Y(n_207)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_105),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_172),
.B(n_526),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_115),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_112),
.B(n_115),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_119),
.C(n_141),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_116),
.B(n_119),
.Y(n_178)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.C(n_131),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_120),
.B(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_122),
.B(n_131),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_123),
.A2(n_124),
.B1(n_128),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_128),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_128),
.A2(n_159),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_132),
.A2(n_133),
.B1(n_167),
.B2(n_168),
.Y(n_188)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_133),
.B(n_247),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_133),
.B(n_308),
.Y(n_429)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_136),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_137),
.B(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_160),
.C(n_164),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.C(n_157),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_143),
.B(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_145),
.B(n_157),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_151),
.C(n_153),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_146),
.A2(n_147),
.B1(n_151),
.B2(n_152),
.Y(n_199)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_154),
.B(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_164),
.Y(n_181)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

AO22x1_ASAP7_75t_SL g212 ( 
.A1(n_165),
.A2(n_166),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_190),
.C(n_193),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_167),
.A2(n_168),
.B1(n_193),
.B2(n_194),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_167),
.B(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_168),
.B(n_436),
.Y(n_465)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_169),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_251),
.B(n_523),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_215),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_176),
.A2(n_524),
.B(n_525),
.Y(n_523)
);

NOR2xp67_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_177),
.B(n_179),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.C(n_184),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_182),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_217),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_200),
.C(n_212),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_185),
.A2(n_186),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.C(n_198),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_187),
.B(n_404),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_189),
.B(n_198),
.Y(n_404)
);

XNOR2x1_ASAP7_75t_L g233 ( 
.A(n_190),
.B(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_191),
.B(n_325),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_191),
.B(n_382),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_193),
.A2(n_194),
.B1(n_292),
.B2(n_293),
.Y(n_375)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_194),
.B(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_197),
.Y(n_196)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_197),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_197),
.Y(n_437)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_197),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_200),
.B(n_212),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_210),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_213),
.Y(n_214)
);

OR2x6_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_216),
.B(n_218),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_222),
.C(n_224),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_219),
.B(n_222),
.Y(n_412)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_220),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_224),
.B(n_412),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_235),
.C(n_239),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_225),
.A2(n_226),
.B1(n_401),
.B2(n_402),
.Y(n_400)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.C(n_232),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_227),
.B(n_350),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_229),
.A2(n_232),
.B1(n_233),
.B2(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_229),
.Y(n_351)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_235),
.A2(n_236),
.B1(n_239),
.B2(n_240),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_241),
.A2(n_242),
.B1(n_357),
.B2(n_358),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_242),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_246),
.C(n_247),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_243),
.A2(n_247),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_243),
.Y(n_307)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_245),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_246),
.B(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_247),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_250),
.Y(n_249)
);

NAND2x1_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_414),
.Y(n_251)
);

A2O1A1O1Ixp25_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_391),
.B(n_407),
.C(n_408),
.D(n_413),
.Y(n_252)
);

OAI21x1_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_363),
.B(n_390),
.Y(n_253)
);

NOR2x1_ASAP7_75t_L g415 ( 
.A(n_254),
.B(n_416),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_343),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g390 ( 
.A(n_255),
.B(n_343),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_304),
.C(n_320),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_256),
.B(n_389),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_275),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_262),
.Y(n_257)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_258),
.Y(n_345)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_262),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_272),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_266),
.B1(n_267),
.B2(n_271),
.Y(n_263)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_264),
.Y(n_271)
);

A2O1A1Ixp33_ASAP7_75t_L g359 ( 
.A1(n_264),
.A2(n_267),
.B(n_272),
.C(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_266),
.B(n_271),
.Y(n_360)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_273),
.B(n_322),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_275),
.B(n_345),
.C(n_346),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_290),
.C(n_297),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_276),
.B(n_369),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_282),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_277),
.B(n_283),
.C(n_286),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_286),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_285),
.Y(n_491)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_289),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_290),
.A2(n_291),
.B1(n_297),
.B2(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_296),
.Y(n_495)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_297),
.Y(n_370)
);

CKINVDCx14_ASAP7_75t_R g374 ( 
.A(n_298),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_300),
.B(n_373),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_303),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_304),
.B(n_320),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_309),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_305),
.B(n_311),
.C(n_319),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_312),
.B2(n_319),
.Y(n_309)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_310),
.Y(n_319)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_312),
.A2(n_324),
.B(n_329),
.Y(n_323)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_317),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_323),
.C(n_334),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_321),
.B(n_323),
.Y(n_366)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_334),
.B(n_366),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.C(n_339),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_335),
.B(n_427),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_336),
.A2(n_337),
.B1(n_339),
.B2(n_340),
.Y(n_427)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_347),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_344),
.B(n_352),
.C(n_393),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_348),
.A2(n_349),
.B1(n_352),
.B2(n_353),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_349),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_353),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_354),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_356),
.A2(n_359),
.B1(n_361),
.B2(n_362),
.Y(n_355)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_356),
.Y(n_361)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_359),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_359),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_361),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_388),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_364),
.B(n_388),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_367),
.C(n_371),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_365),
.B(n_420),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_367),
.A2(n_368),
.B1(n_371),
.B2(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_371),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_375),
.C(n_376),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_372),
.B(n_425),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_375),
.B(n_376),
.Y(n_425)
);

MAJx2_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_381),
.C(n_384),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_377),
.B(n_384),
.Y(n_470)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_381),
.B(n_470),
.Y(n_469)
);

INVx5_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

NAND4xp25_ASAP7_75t_SL g414 ( 
.A(n_391),
.B(n_408),
.C(n_415),
.D(n_417),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_394),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_392),
.B(n_394),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_399),
.Y(n_394)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_395),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.C(n_398),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_400),
.A2(n_403),
.B1(n_405),
.B2(n_406),
.Y(n_399)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_400),
.Y(n_405)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_401),
.Y(n_402)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_403),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_403),
.B(n_405),
.C(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_411),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_409),
.B(n_411),
.Y(n_413)
);

OAI21x1_ASAP7_75t_SL g417 ( 
.A1(n_418),
.A2(n_438),
.B(n_522),
.Y(n_417)
);

NOR2xp67_ASAP7_75t_SL g418 ( 
.A(n_419),
.B(n_422),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_419),
.B(n_422),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_426),
.C(n_428),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_423),
.A2(n_424),
.B1(n_519),
.B2(n_520),
.Y(n_518)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_SL g520 ( 
.A(n_426),
.B(n_428),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.C(n_435),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_429),
.A2(n_430),
.B1(n_431),
.B2(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_429),
.Y(n_473)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx6_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_435),
.B(n_472),
.Y(n_471)
);

AOI21x1_ASAP7_75t_SL g438 ( 
.A1(n_439),
.A2(n_516),
.B(n_521),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_440),
.A2(n_474),
.B(n_515),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_466),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_441),
.B(n_466),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_457),
.C(n_464),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_SL g481 ( 
.A1(n_442),
.A2(n_443),
.B1(n_482),
.B2(n_484),
.Y(n_481)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_453),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_450),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_445),
.B(n_450),
.C(n_453),
.Y(n_468)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_457),
.A2(n_464),
.B1(n_465),
.B2(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_457),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_460),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_458),
.A2(n_459),
.B1(n_460),
.B2(n_461),
.Y(n_477)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_471),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_469),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_468),
.B(n_469),
.C(n_471),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_475),
.A2(n_485),
.B(n_514),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_481),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_476),
.B(n_481),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_478),
.C(n_480),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_477),
.B(n_497),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_478),
.A2(n_479),
.B1(n_480),
.B2(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_480),
.Y(n_498)
);

INVxp67_ASAP7_75t_SL g484 ( 
.A(n_482),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_486),
.A2(n_499),
.B(n_513),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_496),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_487),
.B(n_496),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_492),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_488),
.B(n_492),
.Y(n_504)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_500),
.A2(n_505),
.B(n_512),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_504),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_501),
.B(n_504),
.Y(n_512)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_511),
.Y(n_505)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_518),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_517),
.B(n_518),
.Y(n_521)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);


endmodule