module fake_jpeg_11277_n_512 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_512);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_512;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVxp33_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_10),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_60),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_61),
.B(n_67),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_62),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_15),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_63),
.B(n_75),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_64),
.Y(n_175)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_33),
.B(n_0),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_66),
.B(n_71),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_33),
.B(n_55),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_68),
.Y(n_183)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_70),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_20),
.B(n_14),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_72),
.Y(n_182)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_57),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_78),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_30),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_79),
.B(n_90),
.Y(n_142)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_81),
.Y(n_159)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_82),
.Y(n_192)
);

BUFx8_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx6_ASAP7_75t_SL g134 ( 
.A(n_83),
.Y(n_134)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_84),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_85),
.Y(n_195)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx11_ASAP7_75t_L g189 ( 
.A(n_86),
.Y(n_189)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_87),
.Y(n_169)
);

INVx6_ASAP7_75t_SL g88 ( 
.A(n_30),
.Y(n_88)
);

BUFx16f_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_89),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_30),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_91),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_20),
.B(n_14),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_96),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

INVx6_ASAP7_75t_SL g95 ( 
.A(n_30),
.Y(n_95)
);

BUFx12_ASAP7_75t_L g177 ( 
.A(n_95),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_27),
.B(n_14),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_99),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_100),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_27),
.B(n_0),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_103),
.Y(n_131)
);

INVx5_ASAP7_75t_SL g102 ( 
.A(n_47),
.Y(n_102)
);

INVx2_ASAP7_75t_R g156 ( 
.A(n_102),
.Y(n_156)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_104),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_108),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

NAND2xp33_ASAP7_75t_SL g174 ( 
.A(n_106),
.B(n_107),
.Y(n_174)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_41),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_111),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_34),
.B(n_0),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_113),
.Y(n_126)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_112),
.B(n_114),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_34),
.B(n_0),
.Y(n_113)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_115),
.B(n_116),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_117),
.B(n_118),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_50),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_119),
.B(n_120),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_55),
.B(n_1),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_121),
.B(n_1),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_80),
.A2(n_39),
.B1(n_21),
.B2(n_51),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_127),
.A2(n_130),
.B1(n_194),
.B2(n_13),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_114),
.A2(n_39),
.B1(n_21),
.B2(n_51),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_102),
.A2(n_21),
.B1(n_40),
.B2(n_52),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_135),
.A2(n_145),
.B1(n_146),
.B2(n_158),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_75),
.A2(n_39),
.B1(n_51),
.B2(n_40),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_141),
.A2(n_154),
.B1(n_165),
.B2(n_170),
.Y(n_211)
);

OA22x2_ASAP7_75t_SL g143 ( 
.A1(n_104),
.A2(n_21),
.B1(n_24),
.B2(n_40),
.Y(n_143)
);

NAND2xp67_ASAP7_75t_SL g234 ( 
.A(n_143),
.B(n_134),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_70),
.A2(n_52),
.B1(n_24),
.B2(n_39),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_107),
.A2(n_52),
.B1(n_24),
.B2(n_54),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_26),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_152),
.B(n_172),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_61),
.A2(n_120),
.B1(n_118),
.B2(n_106),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_60),
.A2(n_59),
.B1(n_43),
.B2(n_37),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_L g201 ( 
.A1(n_155),
.A2(n_168),
.B1(n_181),
.B2(n_11),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_63),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_180),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_117),
.A2(n_24),
.B1(n_54),
.B2(n_48),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_64),
.A2(n_24),
.B1(n_43),
.B2(n_37),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_68),
.A2(n_59),
.B1(n_23),
.B2(n_26),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_72),
.A2(n_22),
.B1(n_44),
.B2(n_42),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_74),
.B(n_22),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_85),
.A2(n_48),
.B1(n_44),
.B2(n_42),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_173),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_105),
.A2(n_38),
.B1(n_31),
.B2(n_29),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_176),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_178),
.B(n_6),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_77),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_81),
.A2(n_38),
.B1(n_31),
.B2(n_29),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_89),
.A2(n_28),
.B1(n_23),
.B2(n_5),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_184),
.A2(n_165),
.B1(n_141),
.B2(n_131),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_91),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_148),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_105),
.A2(n_28),
.B1(n_99),
.B2(n_93),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_186),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_100),
.B(n_2),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_188),
.B(n_194),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_83),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_191),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_108),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_125),
.Y(n_197)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_197),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_198),
.B(n_203),
.Y(n_264)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_125),
.Y(n_199)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_199),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_200),
.A2(n_207),
.B1(n_231),
.B2(n_232),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_201),
.B(n_229),
.Y(n_308)
);

O2A1O1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_156),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_L g268 ( 
.A1(n_202),
.A2(n_247),
.B(n_259),
.C(n_261),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_142),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_129),
.B(n_12),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_204),
.B(n_226),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_206),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_L g207 ( 
.A1(n_127),
.A2(n_130),
.B1(n_143),
.B2(n_172),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_124),
.Y(n_208)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_208),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_140),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_209),
.Y(n_263)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_136),
.Y(n_210)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_210),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_212),
.A2(n_216),
.B1(n_244),
.B2(n_254),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_139),
.B(n_138),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_214),
.Y(n_286)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_136),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_184),
.A2(n_131),
.B1(n_129),
.B2(n_143),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_148),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_217),
.Y(n_305)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_148),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_219),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_152),
.B(n_126),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_220),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_221),
.B(n_243),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_126),
.B(n_129),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_222),
.Y(n_296)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_192),
.Y(n_224)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_224),
.Y(n_307)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_124),
.Y(n_225)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_225),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_131),
.B(n_156),
.Y(n_226)
);

INVx11_ASAP7_75t_L g227 ( 
.A(n_134),
.Y(n_227)
);

INVx3_ASAP7_75t_SL g297 ( 
.A(n_227),
.Y(n_297)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_164),
.Y(n_228)
);

INVxp67_ASAP7_75t_SL g301 ( 
.A(n_228),
.Y(n_301)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_164),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_188),
.B(n_123),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_230),
.B(n_257),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_161),
.A2(n_163),
.B1(n_171),
.B2(n_123),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_174),
.A2(n_122),
.B1(n_151),
.B2(n_159),
.Y(n_232)
);

OA22x2_ASAP7_75t_L g262 ( 
.A1(n_234),
.A2(n_261),
.B1(n_227),
.B2(n_212),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_144),
.A2(n_183),
.B1(n_128),
.B2(n_175),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_235),
.A2(n_241),
.B1(n_252),
.B2(n_251),
.Y(n_294)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_193),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_236),
.B(n_240),
.Y(n_283)
);

AND2x2_ASAP7_75t_SL g237 ( 
.A(n_160),
.B(n_195),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_237),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_160),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_239),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_150),
.B(n_132),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_128),
.A2(n_183),
.B1(n_175),
.B2(n_193),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_147),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_242),
.B(n_245),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_149),
.B(n_169),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_122),
.A2(n_151),
.B1(n_159),
.B2(n_187),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_169),
.B(n_149),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_147),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_246),
.B(n_249),
.Y(n_292)
);

O2A1O1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_174),
.A2(n_162),
.B(n_189),
.C(n_177),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_177),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_133),
.B(n_137),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_256),
.Y(n_269)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_187),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_251),
.B(n_255),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_190),
.A2(n_153),
.B1(n_182),
.B2(n_133),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_153),
.B(n_137),
.C(n_195),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_253),
.B(n_237),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_190),
.A2(n_189),
.B1(n_182),
.B2(n_167),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_167),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_179),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_179),
.B(n_177),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_179),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_260),
.Y(n_270)
);

AOI32xp33_ASAP7_75t_L g259 ( 
.A1(n_157),
.A2(n_172),
.A3(n_188),
.B1(n_126),
.B2(n_152),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_134),
.Y(n_260)
);

O2A1O1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_156),
.A2(n_102),
.B(n_143),
.C(n_131),
.Y(n_261)
);

OR2x2_ASAP7_75t_SL g343 ( 
.A(n_262),
.B(n_291),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_211),
.A2(n_221),
.B1(n_207),
.B2(n_223),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_265),
.A2(n_295),
.B1(n_304),
.B2(n_311),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_196),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_272),
.B(n_275),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_243),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_233),
.A2(n_248),
.B1(n_205),
.B2(n_252),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_276),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_233),
.A2(n_248),
.B(n_247),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_278),
.A2(n_256),
.B(n_249),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_281),
.B(n_215),
.C(n_217),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_243),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_288),
.B(n_299),
.Y(n_338)
);

BUFx24_ASAP7_75t_SL g290 ( 
.A(n_203),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_290),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_213),
.B(n_230),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_293),
.B(n_218),
.Y(n_325)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_294),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_211),
.A2(n_213),
.B1(n_238),
.B2(n_259),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_257),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_202),
.A2(n_237),
.B(n_234),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_300),
.A2(n_278),
.B(n_275),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_231),
.B(n_197),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_303),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_199),
.B(n_253),
.Y(n_303)
);

OAI22x1_ASAP7_75t_L g304 ( 
.A1(n_200),
.A2(n_255),
.B1(n_201),
.B2(n_210),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_235),
.A2(n_228),
.B1(n_208),
.B2(n_229),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_241),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_225),
.A2(n_236),
.B1(n_198),
.B2(n_246),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_300),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_313),
.B(n_314),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_270),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_315),
.B(n_327),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_274),
.A2(n_242),
.B1(n_224),
.B2(n_219),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_316),
.A2(n_326),
.B1(n_279),
.B2(n_308),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_317),
.Y(n_372)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_287),
.Y(n_319)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_319),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_320),
.B(n_291),
.C(n_262),
.Y(n_356)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_287),
.Y(n_321)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_321),
.Y(n_355)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_309),
.Y(n_322)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_322),
.Y(n_353)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_309),
.Y(n_323)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_323),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_298),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_324),
.B(n_344),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_325),
.B(n_285),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_274),
.A2(n_302),
.B1(n_265),
.B2(n_273),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_293),
.B(n_273),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_301),
.Y(n_328)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_328),
.Y(n_375)
);

A2O1A1O1Ixp25_ASAP7_75t_L g330 ( 
.A1(n_277),
.A2(n_281),
.B(n_268),
.C(n_296),
.D(n_303),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_330),
.A2(n_337),
.B(n_342),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_295),
.B(n_277),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_332),
.B(n_335),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_305),
.Y(n_333)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_333),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_299),
.B(n_268),
.Y(n_335)
);

INVx13_ASAP7_75t_L g336 ( 
.A(n_297),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_336),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_289),
.B(n_283),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_339),
.B(n_341),
.Y(n_354)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_266),
.Y(n_340)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_340),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_283),
.B(n_272),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_262),
.A2(n_308),
.B(n_292),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_343),
.B(n_349),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_298),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_271),
.B(n_264),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_345),
.B(n_346),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_264),
.B(n_311),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_292),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_347),
.B(n_350),
.Y(n_383)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_266),
.Y(n_349)
);

INVx5_ASAP7_75t_L g350 ( 
.A(n_305),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_284),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_351),
.B(n_305),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_356),
.B(n_363),
.C(n_324),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_357),
.B(n_344),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_334),
.A2(n_294),
.B1(n_304),
.B2(n_262),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_358),
.A2(n_360),
.B1(n_313),
.B2(n_337),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_318),
.A2(n_304),
.B1(n_262),
.B2(n_279),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_362),
.A2(n_365),
.B1(n_374),
.B2(n_379),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_327),
.B(n_282),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_364),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_326),
.A2(n_308),
.B1(n_288),
.B2(n_263),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_335),
.B(n_282),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_368),
.B(n_332),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_345),
.B(n_286),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_373),
.B(n_382),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_318),
.A2(n_280),
.B1(n_297),
.B2(n_267),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_316),
.A2(n_280),
.B1(n_297),
.B2(n_267),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_312),
.A2(n_285),
.B1(n_306),
.B2(n_307),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_381),
.A2(n_323),
.B1(n_349),
.B2(n_340),
.Y(n_409)
);

AND2x6_ASAP7_75t_L g382 ( 
.A(n_330),
.B(n_269),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_376),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_384),
.B(n_391),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_386),
.A2(n_397),
.B(n_370),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_388),
.B(n_405),
.Y(n_429)
);

OAI32xp33_ASAP7_75t_L g389 ( 
.A1(n_371),
.A2(n_312),
.A3(n_346),
.B1(n_338),
.B2(n_331),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_389),
.B(n_393),
.Y(n_411)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_352),
.Y(n_390)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_390),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_383),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_377),
.B(n_320),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_392),
.B(n_398),
.C(n_408),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_361),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_381),
.Y(n_394)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_394),
.Y(n_424)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_353),
.Y(n_396)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_396),
.Y(n_427)
);

OAI22x1_ASAP7_75t_L g397 ( 
.A1(n_365),
.A2(n_343),
.B1(n_342),
.B2(n_317),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_368),
.B(n_330),
.Y(n_398)
);

XNOR2x2_ASAP7_75t_SL g399 ( 
.A(n_377),
.B(n_338),
.Y(n_399)
);

OAI21xp33_ASAP7_75t_L g417 ( 
.A1(n_399),
.A2(n_359),
.B(n_382),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_358),
.A2(n_347),
.B1(n_329),
.B2(n_315),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_400),
.B(n_403),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_373),
.B(n_339),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_401),
.B(n_402),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_367),
.B(n_341),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_359),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_361),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_404),
.B(n_357),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_372),
.A2(n_331),
.B(n_325),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_406),
.A2(n_354),
.B(n_369),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_367),
.B(n_314),
.Y(n_407)
);

CKINVDCx14_ASAP7_75t_R g419 ( 
.A(n_407),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_409),
.A2(n_352),
.B1(n_369),
.B2(n_355),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_371),
.B(n_321),
.Y(n_410)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_410),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_408),
.B(n_356),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_413),
.B(n_428),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_403),
.A2(n_372),
.B(n_386),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_414),
.A2(n_417),
.B(n_418),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_395),
.A2(n_360),
.B1(n_359),
.B2(n_354),
.Y(n_418)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_420),
.Y(n_448)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_421),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_422),
.B(n_397),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_393),
.A2(n_404),
.B1(n_410),
.B2(n_406),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_425),
.A2(n_379),
.B1(n_380),
.B2(n_396),
.Y(n_452)
);

NAND2x1_ASAP7_75t_SL g436 ( 
.A(n_426),
.B(n_399),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_392),
.B(n_363),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_398),
.B(n_362),
.C(n_375),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_431),
.B(n_432),
.C(n_405),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_388),
.B(n_375),
.C(n_355),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_419),
.B(n_384),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_434),
.B(n_442),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_430),
.B(n_348),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_435),
.B(n_443),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_436),
.A2(n_438),
.B(n_412),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_428),
.B(n_399),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_437),
.B(n_439),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_425),
.B(n_387),
.Y(n_440)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_440),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_419),
.B(n_391),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_413),
.B(n_400),
.C(n_385),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_415),
.B(n_390),
.C(n_387),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_444),
.B(n_446),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_415),
.B(n_380),
.C(n_319),
.Y(n_446)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_430),
.Y(n_449)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_449),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_433),
.B(n_389),
.Y(n_450)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_450),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_432),
.B(n_374),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_451),
.B(n_418),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_452),
.B(n_412),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_431),
.B(n_429),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_453),
.B(n_429),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_452),
.B(n_414),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_454),
.A2(n_467),
.B(n_438),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_440),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_455),
.B(n_465),
.Y(n_471)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_460),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_463),
.B(n_464),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_437),
.B(n_429),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_444),
.B(n_446),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_468),
.B(n_469),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_439),
.B(n_422),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_456),
.B(n_416),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_470),
.B(n_476),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_462),
.B(n_441),
.C(n_453),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_472),
.B(n_474),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_466),
.A2(n_450),
.B1(n_411),
.B2(n_416),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_475),
.B(n_426),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_461),
.B(n_441),
.C(n_451),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_461),
.B(n_443),
.C(n_445),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_477),
.B(n_480),
.C(n_463),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_469),
.A2(n_447),
.B(n_411),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_478),
.A2(n_436),
.B(n_457),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_464),
.B(n_445),
.C(n_448),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_476),
.B(n_458),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_482),
.B(n_485),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_474),
.A2(n_467),
.B(n_454),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_484),
.A2(n_487),
.B(n_490),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_472),
.B(n_417),
.Y(n_486)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_486),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_477),
.B(n_459),
.Y(n_487)
);

AO21x1_ASAP7_75t_L g495 ( 
.A1(n_489),
.A2(n_471),
.B(n_454),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_481),
.B(n_447),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_491),
.A2(n_424),
.B1(n_433),
.B2(n_420),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_488),
.B(n_480),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_493),
.B(n_497),
.Y(n_500)
);

AOI31xp67_ASAP7_75t_L g502 ( 
.A1(n_495),
.A2(n_465),
.A3(n_421),
.B(n_423),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_483),
.B(n_479),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_498),
.A2(n_427),
.B1(n_353),
.B2(n_322),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_484),
.A2(n_424),
.B(n_473),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_499),
.A2(n_491),
.B(n_473),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_501),
.A2(n_502),
.B(n_504),
.Y(n_505)
);

OAI21x1_ASAP7_75t_L g503 ( 
.A1(n_494),
.A2(n_423),
.B(n_427),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_503),
.A2(n_495),
.B(n_496),
.Y(n_506)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_506),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_500),
.A2(n_492),
.B(n_493),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_507),
.A2(n_498),
.B1(n_378),
.B2(n_333),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_509),
.Y(n_510)
);

OAI321xp33_ASAP7_75t_L g511 ( 
.A1(n_510),
.A2(n_508),
.A3(n_505),
.B1(n_378),
.B2(n_328),
.C(n_366),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_511),
.A2(n_350),
.B(n_351),
.Y(n_512)
);


endmodule