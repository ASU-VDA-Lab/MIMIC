module fake_netlist_1_761_n_669 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_669);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_669;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_581;
wire n_458;
wire n_504;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_32), .Y(n_77) );
INVx2_ASAP7_75t_L g78 ( .A(n_59), .Y(n_78) );
INVxp67_ASAP7_75t_SL g79 ( .A(n_38), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_54), .Y(n_80) );
INVx1_ASAP7_75t_SL g81 ( .A(n_12), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_20), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_43), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_51), .Y(n_84) );
BUFx3_ASAP7_75t_L g85 ( .A(n_19), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_57), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_53), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_4), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_30), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_61), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_0), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_0), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_68), .Y(n_93) );
CKINVDCx16_ASAP7_75t_R g94 ( .A(n_56), .Y(n_94) );
BUFx2_ASAP7_75t_L g95 ( .A(n_15), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_10), .Y(n_96) );
BUFx5_ASAP7_75t_L g97 ( .A(n_13), .Y(n_97) );
INVxp67_ASAP7_75t_L g98 ( .A(n_10), .Y(n_98) );
CKINVDCx16_ASAP7_75t_R g99 ( .A(n_33), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_25), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_48), .Y(n_101) );
INVxp67_ASAP7_75t_L g102 ( .A(n_47), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_13), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_22), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_17), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_72), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_24), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_73), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_42), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_44), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_71), .Y(n_111) );
INVxp67_ASAP7_75t_L g112 ( .A(n_6), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_35), .Y(n_113) );
HB1xp67_ASAP7_75t_L g114 ( .A(n_26), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_15), .Y(n_115) );
INVxp67_ASAP7_75t_SL g116 ( .A(n_39), .Y(n_116) );
INVxp67_ASAP7_75t_L g117 ( .A(n_16), .Y(n_117) );
INVxp33_ASAP7_75t_SL g118 ( .A(n_19), .Y(n_118) );
INVxp33_ASAP7_75t_SL g119 ( .A(n_40), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_27), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_37), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_62), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_74), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_78), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_80), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_97), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_78), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_105), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_111), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_97), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_95), .B(n_1), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_95), .B(n_1), .Y(n_132) );
XNOR2xp5_ASAP7_75t_L g133 ( .A(n_118), .B(n_2), .Y(n_133) );
NOR2xp33_ASAP7_75t_R g134 ( .A(n_94), .B(n_34), .Y(n_134) );
CKINVDCx16_ASAP7_75t_R g135 ( .A(n_99), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_109), .Y(n_136) );
INVxp67_ASAP7_75t_L g137 ( .A(n_85), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_109), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_104), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_96), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_96), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_119), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_97), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_97), .Y(n_144) );
NOR2xp67_ASAP7_75t_L g145 ( .A(n_114), .B(n_2), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_97), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_97), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_97), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_97), .Y(n_149) );
NAND3xp33_ASAP7_75t_L g150 ( .A(n_115), .B(n_36), .C(n_75), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_85), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_83), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_104), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_83), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_77), .B(n_3), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_102), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_81), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_84), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_108), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_98), .B(n_3), .Y(n_160) );
BUFx2_ASAP7_75t_L g161 ( .A(n_112), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_117), .Y(n_162) );
BUFx2_ASAP7_75t_L g163 ( .A(n_91), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_101), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_108), .Y(n_165) );
AND2x2_ASAP7_75t_SL g166 ( .A(n_131), .B(n_123), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_124), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_131), .B(n_82), .Y(n_168) );
BUFx3_ASAP7_75t_L g169 ( .A(n_151), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_124), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_163), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_163), .Y(n_172) );
OR2x2_ASAP7_75t_L g173 ( .A(n_135), .B(n_92), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_162), .A2(n_82), .B1(n_88), .B2(n_92), .Y(n_174) );
AND2x4_ASAP7_75t_L g175 ( .A(n_137), .B(n_88), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_124), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_126), .Y(n_177) );
AND2x4_ASAP7_75t_L g178 ( .A(n_145), .B(n_103), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_126), .Y(n_179) );
AND2x4_ASAP7_75t_L g180 ( .A(n_145), .B(n_103), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_156), .B(n_107), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_135), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_124), .Y(n_183) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_124), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_126), .Y(n_185) );
INVxp67_ASAP7_75t_L g186 ( .A(n_140), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_126), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_142), .B(n_113), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_136), .B(n_110), .Y(n_189) );
NOR2xp33_ASAP7_75t_SL g190 ( .A(n_138), .B(n_79), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_152), .A2(n_91), .B1(n_122), .B2(n_121), .Y(n_191) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_124), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_127), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_161), .B(n_123), .Y(n_194) );
NOR2xp33_ASAP7_75t_SL g195 ( .A(n_141), .B(n_116), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_164), .B(n_122), .Y(n_196) );
INVx2_ASAP7_75t_SL g197 ( .A(n_144), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_161), .B(n_121), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_144), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_127), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_144), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_144), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_146), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_146), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_127), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_152), .B(n_110), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_146), .Y(n_207) );
NOR2xp33_ASAP7_75t_SL g208 ( .A(n_157), .B(n_120), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_151), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_146), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_147), .Y(n_211) );
INVx1_ASAP7_75t_SL g212 ( .A(n_125), .Y(n_212) );
BUFx3_ASAP7_75t_L g213 ( .A(n_151), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_147), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_154), .B(n_120), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_149), .Y(n_216) );
AND2x6_ASAP7_75t_L g217 ( .A(n_154), .B(n_89), .Y(n_217) );
NOR3xp33_ASAP7_75t_L g218 ( .A(n_132), .B(n_89), .C(n_100), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_149), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_158), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_158), .B(n_106), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_151), .B(n_106), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_153), .Y(n_223) );
OR2x2_ASAP7_75t_SL g224 ( .A(n_160), .B(n_100), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_153), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_153), .B(n_93), .Y(n_226) );
INVx5_ASAP7_75t_L g227 ( .A(n_217), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g228 ( .A1(n_166), .A2(n_155), .B1(n_129), .B2(n_133), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_182), .Y(n_229) );
INVx4_ASAP7_75t_L g230 ( .A(n_217), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_220), .B(n_130), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_175), .B(n_130), .Y(n_232) );
NOR2xp33_ASAP7_75t_R g233 ( .A(n_182), .B(n_128), .Y(n_233) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_212), .Y(n_234) );
INVx3_ASAP7_75t_SL g235 ( .A(n_166), .Y(n_235) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_217), .Y(n_236) );
OR2x6_ASAP7_75t_L g237 ( .A(n_173), .B(n_133), .Y(n_237) );
NOR2xp67_ASAP7_75t_L g238 ( .A(n_186), .B(n_165), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_217), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_209), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_209), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_168), .B(n_175), .Y(n_242) );
BUFx3_ASAP7_75t_L g243 ( .A(n_225), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_175), .B(n_130), .Y(n_244) );
INVx5_ASAP7_75t_L g245 ( .A(n_217), .Y(n_245) );
NOR3xp33_ASAP7_75t_SL g246 ( .A(n_181), .B(n_150), .C(n_86), .Y(n_246) );
INVx5_ASAP7_75t_L g247 ( .A(n_217), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_L g248 ( .A1(n_171), .A2(n_165), .B(n_143), .C(n_148), .Y(n_248) );
INVx2_ASAP7_75t_SL g249 ( .A(n_168), .Y(n_249) );
INVx4_ASAP7_75t_L g250 ( .A(n_169), .Y(n_250) );
NOR2x1p5_ASAP7_75t_L g251 ( .A(n_173), .B(n_84), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_174), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_168), .B(n_134), .Y(n_253) );
XNOR2xp5_ASAP7_75t_L g254 ( .A(n_224), .B(n_4), .Y(n_254) );
BUFx2_ASAP7_75t_L g255 ( .A(n_194), .Y(n_255) );
CKINVDCx6p67_ASAP7_75t_R g256 ( .A(n_196), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_221), .B(n_143), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_208), .B(n_86), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_172), .B(n_87), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_206), .A2(n_165), .B(n_143), .C(n_148), .Y(n_260) );
OR2x6_ASAP7_75t_L g261 ( .A(n_178), .B(n_93), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_218), .B(n_148), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_209), .Y(n_263) );
INVx3_ASAP7_75t_L g264 ( .A(n_225), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_178), .B(n_90), .Y(n_265) );
OR2x6_ASAP7_75t_SL g266 ( .A(n_195), .B(n_87), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_178), .A2(n_159), .B1(n_139), .B2(n_127), .Y(n_267) );
INVxp33_ASAP7_75t_L g268 ( .A(n_194), .Y(n_268) );
CKINVDCx16_ASAP7_75t_R g269 ( .A(n_190), .Y(n_269) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_198), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_221), .B(n_90), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_225), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_223), .Y(n_273) );
BUFx3_ASAP7_75t_L g274 ( .A(n_169), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g275 ( .A1(n_198), .A2(n_159), .B1(n_139), .B2(n_127), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_188), .Y(n_276) );
A2O1A1Ixp33_ASAP7_75t_L g277 ( .A1(n_215), .A2(n_139), .B(n_127), .C(n_159), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_180), .B(n_159), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_180), .B(n_159), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_180), .B(n_159), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_226), .Y(n_281) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_213), .Y(n_282) );
NOR3xp33_ASAP7_75t_SL g283 ( .A(n_189), .B(n_5), .C(n_6), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_191), .B(n_139), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_211), .B(n_139), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_222), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_211), .B(n_139), .Y(n_287) );
INVx5_ASAP7_75t_L g288 ( .A(n_183), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_213), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_167), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_167), .Y(n_291) );
CKINVDCx20_ASAP7_75t_R g292 ( .A(n_234), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_230), .B(n_177), .Y(n_293) );
INVx3_ASAP7_75t_L g294 ( .A(n_230), .Y(n_294) );
INVx1_ASAP7_75t_SL g295 ( .A(n_236), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_285), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_285), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_287), .Y(n_298) );
CKINVDCx20_ASAP7_75t_R g299 ( .A(n_229), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_287), .Y(n_300) );
BUFx2_ASAP7_75t_SL g301 ( .A(n_236), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_273), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_257), .Y(n_303) );
AOI21x1_ASAP7_75t_L g304 ( .A1(n_231), .A2(n_170), .B(n_193), .Y(n_304) );
BUFx3_ASAP7_75t_L g305 ( .A(n_236), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_235), .B(n_214), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_286), .B(n_202), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_240), .Y(n_308) );
AOI222xp33_ASAP7_75t_L g309 ( .A1(n_252), .A2(n_255), .B1(n_270), .B2(n_268), .C1(n_254), .C2(n_242), .Y(n_309) );
BUFx12f_ASAP7_75t_L g310 ( .A(n_239), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_257), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_241), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_239), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_281), .B(n_214), .Y(n_314) );
AND2x4_ASAP7_75t_SL g315 ( .A(n_239), .B(n_201), .Y(n_315) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_251), .A2(n_216), .B1(n_219), .B2(n_203), .Y(n_316) );
INVx3_ASAP7_75t_L g317 ( .A(n_282), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_263), .Y(n_318) );
AO31x2_ASAP7_75t_L g319 ( .A1(n_260), .A2(n_170), .A3(n_193), .B(n_176), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_249), .B(n_216), .Y(n_320) );
AOI21xp33_ASAP7_75t_L g321 ( .A1(n_253), .A2(n_276), .B(n_261), .Y(n_321) );
INVxp67_ASAP7_75t_L g322 ( .A(n_266), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_232), .A2(n_197), .B(n_187), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_261), .A2(n_219), .B1(n_203), .B2(n_202), .Y(n_324) );
INVxp67_ASAP7_75t_SL g325 ( .A(n_282), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_232), .A2(n_197), .B(n_201), .Y(n_326) );
AND2x4_ASAP7_75t_L g327 ( .A(n_238), .B(n_177), .Y(n_327) );
CKINVDCx16_ASAP7_75t_R g328 ( .A(n_233), .Y(n_328) );
A2O1A1Ixp33_ASAP7_75t_L g329 ( .A1(n_248), .A2(n_187), .B(n_179), .C(n_207), .Y(n_329) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_227), .Y(n_330) );
BUFx3_ASAP7_75t_L g331 ( .A(n_282), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_272), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_261), .A2(n_179), .B1(n_210), .B2(n_204), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_271), .A2(n_224), .B1(n_185), .B2(n_199), .Y(n_334) );
BUFx4_ASAP7_75t_SL g335 ( .A(n_237), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_271), .B(n_5), .Y(n_336) );
CKINVDCx8_ASAP7_75t_R g337 ( .A(n_269), .Y(n_337) );
NAND3xp33_ASAP7_75t_L g338 ( .A(n_283), .B(n_205), .C(n_200), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_250), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_231), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_244), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_296), .Y(n_342) );
A2O1A1Ixp33_ASAP7_75t_L g343 ( .A1(n_340), .A2(n_259), .B(n_262), .C(n_244), .Y(n_343) );
NAND2xp33_ASAP7_75t_R g344 ( .A(n_335), .B(n_237), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_321), .B(n_237), .Y(n_345) );
CKINVDCx6p67_ASAP7_75t_R g346 ( .A(n_292), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_303), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_303), .B(n_228), .Y(n_348) );
INVx1_ASAP7_75t_SL g349 ( .A(n_299), .Y(n_349) );
AOI21x1_ASAP7_75t_L g350 ( .A1(n_304), .A2(n_258), .B(n_278), .Y(n_350) );
INVx3_ASAP7_75t_L g351 ( .A(n_310), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_328), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_311), .Y(n_353) );
BUFx3_ASAP7_75t_L g354 ( .A(n_310), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_311), .Y(n_355) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_306), .Y(n_356) );
AND2x4_ASAP7_75t_L g357 ( .A(n_306), .B(n_227), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_340), .B(n_256), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_314), .Y(n_359) );
AND2x6_ASAP7_75t_L g360 ( .A(n_294), .B(n_284), .Y(n_360) );
AO31x2_ASAP7_75t_L g361 ( .A1(n_334), .A2(n_277), .A3(n_280), .B(n_279), .Y(n_361) );
OAI21x1_ASAP7_75t_SL g362 ( .A1(n_302), .A2(n_278), .B(n_279), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_341), .A2(n_243), .B1(n_280), .B2(n_250), .Y(n_363) );
OAI21x1_ASAP7_75t_L g364 ( .A1(n_304), .A2(n_275), .B(n_267), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_314), .B(n_265), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_336), .Y(n_366) );
NAND2xp33_ASAP7_75t_R g367 ( .A(n_317), .B(n_246), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_341), .Y(n_368) );
AOI221xp5_ASAP7_75t_L g369 ( .A1(n_322), .A2(n_264), .B1(n_289), .B2(n_274), .C(n_291), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_302), .Y(n_370) );
OAI22xp5_ASAP7_75t_L g371 ( .A1(n_316), .A2(n_302), .B1(n_307), .B2(n_324), .Y(n_371) );
INVx3_ASAP7_75t_L g372 ( .A(n_310), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_345), .A2(n_309), .B1(n_338), .B2(n_328), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_347), .B(n_296), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_356), .Y(n_375) );
AOI221xp5_ASAP7_75t_L g376 ( .A1(n_359), .A2(n_334), .B1(n_316), .B2(n_338), .C(n_320), .Y(n_376) );
BUFx4f_ASAP7_75t_SL g377 ( .A(n_346), .Y(n_377) );
BUFx4f_ASAP7_75t_SL g378 ( .A(n_346), .Y(n_378) );
OAI22xp5_ASAP7_75t_SL g379 ( .A1(n_352), .A2(n_337), .B1(n_309), .B2(n_333), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_370), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_348), .A2(n_327), .B1(n_320), .B2(n_308), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g382 ( .A1(n_343), .A2(n_300), .B1(n_298), .B2(n_297), .Y(n_382) );
INVxp67_ASAP7_75t_L g383 ( .A(n_358), .Y(n_383) );
BUFx3_ASAP7_75t_L g384 ( .A(n_354), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_353), .B(n_296), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_348), .A2(n_366), .B1(n_371), .B2(n_358), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_354), .Y(n_387) );
NAND2xp33_ASAP7_75t_SL g388 ( .A(n_351), .B(n_313), .Y(n_388) );
OAI21x1_ASAP7_75t_L g389 ( .A1(n_350), .A2(n_323), .B(n_326), .Y(n_389) );
AO31x2_ASAP7_75t_L g390 ( .A1(n_343), .A2(n_329), .A3(n_300), .B(n_297), .Y(n_390) );
INVx2_ASAP7_75t_SL g391 ( .A(n_351), .Y(n_391) );
AOI22xp33_ASAP7_75t_SL g392 ( .A1(n_355), .A2(n_337), .B1(n_327), .B2(n_300), .Y(n_392) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_368), .A2(n_327), .B1(n_297), .B2(n_298), .C(n_332), .Y(n_393) );
NAND3xp33_ASAP7_75t_L g394 ( .A(n_363), .B(n_308), .C(n_312), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_342), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_342), .A2(n_298), .B(n_318), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_362), .Y(n_397) );
OAI22xp33_ASAP7_75t_L g398 ( .A1(n_344), .A2(n_294), .B1(n_308), .B2(n_312), .Y(n_398) );
INVx2_ASAP7_75t_SL g399 ( .A(n_351), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_364), .Y(n_400) );
OAI321xp33_ASAP7_75t_L g401 ( .A1(n_373), .A2(n_365), .A3(n_369), .B1(n_332), .B2(n_318), .C(n_312), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_395), .Y(n_402) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_392), .B(n_372), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_380), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_380), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_386), .A2(n_372), .B1(n_332), .B2(n_357), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_395), .B(n_361), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_395), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_400), .Y(n_409) );
AOI211xp5_ASAP7_75t_L g410 ( .A1(n_379), .A2(n_398), .B(n_383), .C(n_387), .Y(n_410) );
NOR2xp33_ASAP7_75t_R g411 ( .A(n_377), .B(n_352), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_374), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_374), .B(n_361), .Y(n_413) );
AOI211xp5_ASAP7_75t_L g414 ( .A1(n_379), .A2(n_349), .B(n_372), .C(n_357), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_397), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_400), .Y(n_416) );
OAI211xp5_ASAP7_75t_L g417 ( .A1(n_392), .A2(n_375), .B(n_381), .C(n_384), .Y(n_417) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_397), .Y(n_418) );
INVxp67_ASAP7_75t_L g419 ( .A(n_385), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_384), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_385), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_390), .B(n_361), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_400), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g424 ( .A1(n_382), .A2(n_327), .B1(n_357), .B2(n_318), .C(n_264), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_390), .B(n_361), .Y(n_425) );
CKINVDCx5p33_ASAP7_75t_R g426 ( .A(n_378), .Y(n_426) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_384), .Y(n_427) );
AOI221xp5_ASAP7_75t_L g428 ( .A1(n_382), .A2(n_339), .B1(n_293), .B2(n_325), .C(n_317), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_390), .B(n_361), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_390), .Y(n_430) );
INVx2_ASAP7_75t_SL g431 ( .A(n_391), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_390), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_390), .Y(n_433) );
AOI21xp33_ASAP7_75t_SL g434 ( .A1(n_391), .A2(n_367), .B(n_8), .Y(n_434) );
AO21x2_ASAP7_75t_L g435 ( .A1(n_394), .A2(n_364), .B(n_176), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_415), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_402), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_402), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_420), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_421), .B(n_393), .Y(n_440) );
AOI221xp5_ASAP7_75t_L g441 ( .A1(n_410), .A2(n_376), .B1(n_393), .B2(n_399), .C(n_394), .Y(n_441) );
INVx2_ASAP7_75t_SL g442 ( .A(n_427), .Y(n_442) );
NAND4xp25_ASAP7_75t_L g443 ( .A(n_410), .B(n_376), .C(n_396), .D(n_9), .Y(n_443) );
INVx3_ASAP7_75t_L g444 ( .A(n_402), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_419), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_426), .B(n_399), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_407), .B(n_396), .Y(n_447) );
INVx1_ASAP7_75t_SL g448 ( .A(n_411), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_414), .A2(n_339), .B1(n_331), .B2(n_317), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_415), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_408), .Y(n_451) );
NAND3xp33_ASAP7_75t_L g452 ( .A(n_414), .B(n_388), .C(n_183), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_413), .B(n_319), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_406), .A2(n_360), .B1(n_339), .B2(n_331), .Y(n_454) );
NOR3xp33_ASAP7_75t_SL g455 ( .A(n_417), .B(n_7), .C(n_8), .Y(n_455) );
OAI31xp33_ASAP7_75t_L g456 ( .A1(n_417), .A2(n_339), .A3(n_315), .B(n_293), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_407), .B(n_319), .Y(n_457) );
OAI31xp33_ASAP7_75t_L g458 ( .A1(n_406), .A2(n_315), .A3(n_293), .B(n_331), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_404), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_424), .A2(n_360), .B1(n_389), .B2(n_317), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_407), .B(n_319), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_404), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_413), .B(n_419), .Y(n_463) );
AOI221xp5_ASAP7_75t_L g464 ( .A1(n_434), .A2(n_183), .B1(n_184), .B2(n_192), .C(n_200), .Y(n_464) );
NAND3xp33_ASAP7_75t_L g465 ( .A(n_434), .B(n_183), .C(n_184), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_421), .B(n_319), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_422), .B(n_319), .Y(n_467) );
OAI31xp33_ASAP7_75t_SL g468 ( .A1(n_403), .A2(n_389), .A3(n_295), .B(n_360), .Y(n_468) );
INVxp67_ASAP7_75t_SL g469 ( .A(n_408), .Y(n_469) );
NAND3xp33_ASAP7_75t_SL g470 ( .A(n_424), .B(n_295), .C(n_9), .Y(n_470) );
INVx4_ASAP7_75t_L g471 ( .A(n_431), .Y(n_471) );
NOR2x1p5_ASAP7_75t_L g472 ( .A(n_412), .B(n_408), .Y(n_472) );
AND2x4_ASAP7_75t_SL g473 ( .A(n_412), .B(n_313), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_409), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_405), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_405), .Y(n_476) );
OAI31xp33_ASAP7_75t_L g477 ( .A1(n_418), .A2(n_315), .A3(n_293), .B(n_294), .Y(n_477) );
INVx2_ASAP7_75t_SL g478 ( .A(n_431), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_422), .B(n_319), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_409), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_418), .Y(n_481) );
INVxp67_ASAP7_75t_L g482 ( .A(n_431), .Y(n_482) );
BUFx3_ASAP7_75t_L g483 ( .A(n_409), .Y(n_483) );
AOI221xp5_ASAP7_75t_L g484 ( .A1(n_401), .A2(n_430), .B1(n_432), .B2(n_422), .C(n_429), .Y(n_484) );
OAI221xp5_ASAP7_75t_L g485 ( .A1(n_428), .A2(n_294), .B1(n_184), .B2(n_192), .C(n_200), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_472), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_463), .B(n_429), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_439), .B(n_425), .Y(n_488) );
NOR2xp33_ASAP7_75t_R g489 ( .A(n_470), .B(n_360), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_455), .A2(n_428), .B1(n_430), .B2(n_432), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_463), .B(n_429), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_452), .B(n_401), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_445), .B(n_469), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_459), .B(n_425), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_459), .B(n_425), .Y(n_495) );
INVx4_ASAP7_75t_L g496 ( .A(n_471), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_462), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_462), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_443), .A2(n_433), .B1(n_360), .B2(n_423), .Y(n_499) );
NOR2xp33_ASAP7_75t_R g500 ( .A(n_448), .B(n_442), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_444), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_447), .B(n_423), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_467), .B(n_7), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_444), .B(n_423), .Y(n_504) );
INVx4_ASAP7_75t_L g505 ( .A(n_471), .Y(n_505) );
NAND3xp33_ASAP7_75t_L g506 ( .A(n_443), .B(n_183), .C(n_184), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_444), .B(n_416), .Y(n_507) );
INVx1_ASAP7_75t_SL g508 ( .A(n_442), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_478), .B(n_416), .Y(n_509) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_483), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_475), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_452), .B(n_416), .Y(n_512) );
NAND2x1p5_ASAP7_75t_L g513 ( .A(n_471), .B(n_313), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_475), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_474), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_478), .B(n_435), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_476), .B(n_435), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_446), .Y(n_518) );
OAI211xp5_ASAP7_75t_SL g519 ( .A1(n_456), .A2(n_11), .B(n_12), .C(n_14), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_481), .B(n_435), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_474), .Y(n_521) );
BUFx2_ASAP7_75t_L g522 ( .A(n_471), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_476), .B(n_440), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_436), .Y(n_524) );
INVx1_ASAP7_75t_SL g525 ( .A(n_473), .Y(n_525) );
BUFx2_ASAP7_75t_L g526 ( .A(n_482), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_467), .B(n_11), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_437), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_436), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_450), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_450), .B(n_14), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_456), .B(n_468), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_481), .Y(n_533) );
NAND2xp33_ASAP7_75t_SL g534 ( .A(n_454), .B(n_435), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_437), .B(n_16), .Y(n_535) );
INVx1_ASAP7_75t_SL g536 ( .A(n_473), .Y(n_536) );
OAI31xp33_ASAP7_75t_L g537 ( .A1(n_465), .A2(n_17), .A3(n_18), .B(n_20), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_483), .Y(n_538) );
AOI31xp33_ASAP7_75t_L g539 ( .A1(n_465), .A2(n_18), .A3(n_21), .B(n_360), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_479), .B(n_21), .Y(n_540) );
AND2x4_ASAP7_75t_L g541 ( .A(n_479), .B(n_389), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_533), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_523), .B(n_484), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_488), .B(n_461), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_497), .Y(n_545) );
INVx1_ASAP7_75t_SL g546 ( .A(n_500), .Y(n_546) );
AOI21xp5_ASAP7_75t_SL g547 ( .A1(n_532), .A2(n_441), .B(n_464), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_498), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_493), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_539), .A2(n_460), .B1(n_453), .B2(n_485), .Y(n_550) );
OAI21xp33_ASAP7_75t_L g551 ( .A1(n_532), .A2(n_466), .B(n_453), .Y(n_551) );
INVx2_ASAP7_75t_SL g552 ( .A(n_500), .Y(n_552) );
INVx1_ASAP7_75t_SL g553 ( .A(n_518), .Y(n_553) );
O2A1O1Ixp33_ASAP7_75t_L g554 ( .A1(n_519), .A2(n_477), .B(n_458), .C(n_449), .Y(n_554) );
OAI21xp33_ASAP7_75t_L g555 ( .A1(n_492), .A2(n_461), .B(n_457), .Y(n_555) );
O2A1O1Ixp33_ASAP7_75t_L g556 ( .A1(n_519), .A2(n_477), .B(n_458), .C(n_451), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_511), .Y(n_557) );
NAND2xp33_ASAP7_75t_SL g558 ( .A(n_496), .B(n_451), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_508), .B(n_457), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_499), .A2(n_438), .B1(n_480), .B2(n_305), .Y(n_560) );
XNOR2x1_ASAP7_75t_L g561 ( .A(n_503), .B(n_438), .Y(n_561) );
AOI32xp33_ASAP7_75t_L g562 ( .A1(n_531), .A2(n_480), .A3(n_305), .B1(n_29), .B2(n_31), .Y(n_562) );
OAI21xp5_ASAP7_75t_L g563 ( .A1(n_506), .A2(n_247), .B(n_245), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_514), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_526), .B(n_23), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_524), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_512), .A2(n_313), .B(n_305), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_489), .A2(n_184), .B1(n_192), .B2(n_200), .Y(n_568) );
OAI221xp5_ASAP7_75t_SL g569 ( .A1(n_537), .A2(n_28), .B1(n_41), .B2(n_45), .C(n_46), .Y(n_569) );
OAI221xp5_ASAP7_75t_L g570 ( .A1(n_531), .A2(n_192), .B1(n_200), .B2(n_205), .C(n_301), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_529), .Y(n_571) );
AO211x2_ASAP7_75t_L g572 ( .A1(n_540), .A2(n_49), .B(n_50), .C(n_52), .Y(n_572) );
AOI22xp33_ASAP7_75t_SL g573 ( .A1(n_496), .A2(n_301), .B1(n_313), .B2(n_330), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_530), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_523), .B(n_205), .Y(n_575) );
XOR2x2_ASAP7_75t_L g576 ( .A(n_527), .B(n_55), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_492), .A2(n_192), .B1(n_205), .B2(n_313), .Y(n_577) );
OAI22xp33_ASAP7_75t_L g578 ( .A1(n_505), .A2(n_330), .B1(n_247), .B2(n_245), .Y(n_578) );
INVxp67_ASAP7_75t_L g579 ( .A(n_522), .Y(n_579) );
AOI321xp33_ASAP7_75t_L g580 ( .A1(n_490), .A2(n_58), .A3(n_60), .B1(n_63), .B2(n_64), .C(n_65), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_494), .B(n_205), .Y(n_581) );
AOI22xp33_ASAP7_75t_SL g582 ( .A1(n_505), .A2(n_330), .B1(n_227), .B2(n_245), .Y(n_582) );
AOI21xp33_ASAP7_75t_L g583 ( .A1(n_535), .A2(n_66), .B(n_67), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_487), .B(n_69), .Y(n_584) );
NAND4xp25_ASAP7_75t_L g585 ( .A(n_534), .B(n_290), .C(n_70), .D(n_76), .Y(n_585) );
OAI221xp5_ASAP7_75t_L g586 ( .A1(n_534), .A2(n_330), .B1(n_288), .B2(n_247), .C(n_245), .Y(n_586) );
OAI22xp33_ASAP7_75t_L g587 ( .A1(n_525), .A2(n_330), .B1(n_247), .B2(n_227), .Y(n_587) );
INVx1_ASAP7_75t_SL g588 ( .A(n_536), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_541), .A2(n_288), .B1(n_330), .B2(n_486), .Y(n_589) );
OAI211xp5_ASAP7_75t_L g590 ( .A1(n_489), .A2(n_288), .B(n_512), .C(n_538), .Y(n_590) );
O2A1O1Ixp33_ASAP7_75t_L g591 ( .A1(n_510), .A2(n_288), .B(n_538), .C(n_520), .Y(n_591) );
NOR4xp25_ASAP7_75t_SL g592 ( .A(n_558), .B(n_513), .C(n_516), .D(n_509), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_545), .Y(n_593) );
AOI211xp5_ASAP7_75t_SL g594 ( .A1(n_590), .A2(n_541), .B(n_495), .C(n_491), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_548), .Y(n_595) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_581), .Y(n_596) );
INVx1_ASAP7_75t_SL g597 ( .A(n_546), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_557), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_543), .B(n_502), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_564), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_549), .B(n_517), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_566), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_544), .B(n_501), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_571), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_551), .B(n_515), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_542), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_574), .Y(n_607) );
NOR4xp25_ASAP7_75t_SL g608 ( .A(n_586), .B(n_513), .C(n_507), .D(n_504), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_591), .Y(n_609) );
INVx3_ASAP7_75t_SL g610 ( .A(n_552), .Y(n_610) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_579), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_588), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_591), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_575), .Y(n_614) );
NOR3xp33_ASAP7_75t_SL g615 ( .A(n_590), .B(n_515), .C(n_521), .Y(n_615) );
XNOR2x1_ASAP7_75t_L g616 ( .A(n_576), .B(n_528), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_559), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_555), .B(n_521), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_589), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_561), .B(n_553), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_560), .B(n_550), .Y(n_621) );
INVxp33_ASAP7_75t_L g622 ( .A(n_584), .Y(n_622) );
INVxp67_ASAP7_75t_L g623 ( .A(n_565), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_547), .B(n_556), .Y(n_624) );
NAND3xp33_ASAP7_75t_L g625 ( .A(n_580), .B(n_562), .C(n_585), .Y(n_625) );
OAI322xp33_ASAP7_75t_L g626 ( .A1(n_624), .A2(n_554), .A3(n_556), .B1(n_570), .B2(n_577), .C1(n_587), .C2(n_578), .Y(n_626) );
NAND2x1_ASAP7_75t_L g627 ( .A(n_615), .B(n_568), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g628 ( .A1(n_594), .A2(n_554), .B(n_563), .Y(n_628) );
AND2x4_ASAP7_75t_L g629 ( .A(n_613), .B(n_567), .Y(n_629) );
NAND3xp33_ASAP7_75t_L g630 ( .A(n_624), .B(n_569), .C(n_583), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_599), .B(n_567), .Y(n_631) );
OR2x2_ASAP7_75t_L g632 ( .A(n_601), .B(n_573), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_610), .Y(n_633) );
AND2x4_ASAP7_75t_L g634 ( .A(n_609), .B(n_572), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_617), .B(n_582), .Y(n_635) );
AOI322xp5_ASAP7_75t_L g636 ( .A1(n_621), .A2(n_620), .A3(n_597), .B1(n_617), .B2(n_609), .C1(n_612), .C2(n_611), .Y(n_636) );
BUFx3_ASAP7_75t_L g637 ( .A(n_610), .Y(n_637) );
XNOR2xp5_ASAP7_75t_L g638 ( .A(n_616), .B(n_621), .Y(n_638) );
AOI211xp5_ASAP7_75t_L g639 ( .A1(n_625), .A2(n_622), .B(n_623), .C(n_619), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_619), .A2(n_616), .B1(n_614), .B2(n_596), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_595), .Y(n_641) );
NOR3x1_ASAP7_75t_L g642 ( .A(n_605), .B(n_601), .C(n_606), .Y(n_642) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_592), .A2(n_608), .B(n_618), .Y(n_643) );
AND2x4_ASAP7_75t_L g644 ( .A(n_642), .B(n_614), .Y(n_644) );
AOI21xp33_ASAP7_75t_SL g645 ( .A1(n_638), .A2(n_618), .B(n_607), .Y(n_645) );
AOI221xp5_ASAP7_75t_SL g646 ( .A1(n_639), .A2(n_593), .B1(n_604), .B2(n_598), .C(n_602), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g647 ( .A1(n_640), .A2(n_598), .B1(n_600), .B2(n_602), .C(n_604), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_631), .B(n_600), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_637), .Y(n_649) );
OAI211xp5_ASAP7_75t_SL g650 ( .A1(n_636), .A2(n_596), .B(n_603), .C(n_640), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_630), .A2(n_596), .B1(n_635), .B2(n_628), .Y(n_651) );
NAND4xp25_ASAP7_75t_L g652 ( .A(n_643), .B(n_633), .C(n_634), .D(n_629), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_634), .A2(n_632), .B1(n_627), .B2(n_629), .Y(n_653) );
OAI221xp5_ASAP7_75t_L g654 ( .A1(n_641), .A2(n_640), .B1(n_638), .B2(n_636), .C(n_639), .Y(n_654) );
A2O1A1Ixp33_ASAP7_75t_L g655 ( .A1(n_634), .A2(n_637), .B(n_636), .C(n_633), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_626), .A2(n_624), .B1(n_621), .B2(n_634), .Y(n_656) );
XOR2x1_ASAP7_75t_L g657 ( .A(n_644), .B(n_649), .Y(n_657) );
NAND3xp33_ASAP7_75t_L g658 ( .A(n_655), .B(n_651), .C(n_652), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_648), .Y(n_659) );
XOR2xp5_ASAP7_75t_L g660 ( .A(n_656), .B(n_653), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_659), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_657), .Y(n_662) );
OAI221xp5_ASAP7_75t_L g663 ( .A1(n_658), .A2(n_654), .B1(n_650), .B2(n_646), .C(n_647), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_661), .B(n_660), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_662), .Y(n_665) );
INVxp67_ASAP7_75t_SL g666 ( .A(n_665), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_664), .Y(n_667) );
BUFx2_ASAP7_75t_L g668 ( .A(n_666), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_668), .A2(n_663), .B1(n_667), .B2(n_645), .C(n_646), .Y(n_669) );
endmodule