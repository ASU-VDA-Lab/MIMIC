module fake_jpeg_31974_n_186 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_186);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_49),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_19),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_39),
.A2(n_33),
.B1(n_16),
.B2(n_24),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_50),
.B(n_33),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_25),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_18),
.B1(n_21),
.B2(n_25),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_54),
.A2(n_55),
.B1(n_65),
.B2(n_67),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_25),
.B1(n_31),
.B2(n_19),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_49),
.B(n_17),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_71),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_34),
.B(n_30),
.C(n_29),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_32),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_16),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_62),
.B(n_27),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_25),
.B1(n_31),
.B2(n_34),
.Y(n_65)
);

O2A1O1Ixp33_ASAP7_75t_SL g68 ( 
.A1(n_41),
.A2(n_17),
.B(n_32),
.C(n_24),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_68),
.A2(n_59),
.B1(n_52),
.B2(n_71),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_14),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_44),
.B(n_1),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_68),
.A2(n_47),
.B1(n_30),
.B2(n_22),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_76),
.A2(n_78),
.B1(n_97),
.B2(n_98),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_29),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_83),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_53),
.A2(n_22),
.B1(n_45),
.B2(n_51),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_80),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_67),
.A2(n_27),
.B1(n_32),
.B2(n_4),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_82),
.A2(n_89),
.B1(n_90),
.B2(n_56),
.Y(n_110)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_32),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_87),
.B(n_88),
.Y(n_108)
);

AO22x1_ASAP7_75t_L g90 ( 
.A1(n_60),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_5),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_92),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_93),
.Y(n_114)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_99),
.Y(n_112)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_82),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_53),
.B1(n_73),
.B2(n_75),
.Y(n_111)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_112),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_125),
.Y(n_136)
);

NOR3xp33_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_90),
.C(n_88),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_117),
.B(n_118),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_108),
.B(n_103),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

A2O1A1O1Ixp25_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_77),
.B(n_90),
.C(n_89),
.D(n_81),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_121),
.A2(n_124),
.B(n_102),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_122),
.A2(n_110),
.B1(n_83),
.B2(n_111),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_106),
.A2(n_85),
.B(n_92),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_123),
.A2(n_63),
.B(n_113),
.Y(n_134)
);

NOR2x1_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_85),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_81),
.C(n_83),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_101),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_126),
.B(n_127),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_99),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_128),
.A2(n_96),
.B1(n_113),
.B2(n_109),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_130),
.B(n_125),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_124),
.A2(n_100),
.B(n_105),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_134),
.B(n_123),
.Y(n_144)
);

AO22x2_ASAP7_75t_L g132 ( 
.A1(n_119),
.A2(n_115),
.B1(n_116),
.B2(n_122),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_132),
.B(n_115),
.Y(n_147)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_138),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_144),
.Y(n_151)
);

NAND4xp25_ASAP7_75t_SL g145 ( 
.A(n_132),
.B(n_59),
.C(n_64),
.D(n_98),
.Y(n_145)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_118),
.B(n_124),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_146),
.A2(n_131),
.B(n_130),
.C(n_136),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_148),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_121),
.B1(n_100),
.B2(n_109),
.Y(n_148)
);

AOI322xp5_ASAP7_75t_L g154 ( 
.A1(n_149),
.A2(n_132),
.A3(n_139),
.B1(n_128),
.B2(n_134),
.C1(n_75),
.C2(n_73),
.Y(n_154)
);

XNOR2x2_ASAP7_75t_SL g161 ( 
.A(n_150),
.B(n_158),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_157),
.Y(n_165)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

NOR3xp33_ASAP7_75t_SL g157 ( 
.A(n_146),
.B(n_132),
.C(n_114),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_132),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_143),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_160),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_141),
.C(n_104),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_105),
.C(n_104),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_156),
.Y(n_168)
);

AOI21xp33_ASAP7_75t_SL g163 ( 
.A1(n_157),
.A2(n_138),
.B(n_135),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_163),
.A2(n_80),
.B1(n_79),
.B2(n_56),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_158),
.A2(n_133),
.B(n_113),
.Y(n_164)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_164),
.Y(n_170)
);

AOI22x1_ASAP7_75t_L g167 ( 
.A1(n_161),
.A2(n_153),
.B1(n_156),
.B2(n_63),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_167),
.A2(n_169),
.B(n_165),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_171),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_64),
.B1(n_14),
.B2(n_13),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_168),
.B(n_166),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_175),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_160),
.Y(n_175)
);

NAND4xp25_ASAP7_75t_SL g176 ( 
.A(n_171),
.B(n_5),
.C(n_6),
.D(n_8),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_9),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_177),
.A2(n_174),
.B1(n_176),
.B2(n_167),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_179),
.C(n_172),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_181),
.A2(n_182),
.B(n_13),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_159),
.C(n_12),
.Y(n_182)
);

MAJx2_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_11),
.C(n_9),
.Y(n_184)
);

BUFx24_ASAP7_75t_SL g185 ( 
.A(n_184),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_185),
.B(n_10),
.Y(n_186)
);


endmodule