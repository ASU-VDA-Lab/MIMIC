module fake_jpeg_12807_n_73 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_73);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_73;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_51;
wire n_47;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_23),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_0),
.Y(n_35)
);

NOR3xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_13),
.C(n_24),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_30),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_28),
.B(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_39),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_43)
);

NOR2x1_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_17),
.Y(n_56)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_33),
.B1(n_25),
.B2(n_27),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_27),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_51),
.C(n_54),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_48),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_58),
.B1(n_20),
.B2(n_21),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_3),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_56),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_4),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_43),
.B(n_6),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_7),
.C(n_9),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_47),
.B(n_7),
.Y(n_58)
);

AO22x1_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_47),
.B1(n_48),
.B2(n_11),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_61),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_12),
.Y(n_63)
);

OAI22x1_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_64),
.B1(n_65),
.B2(n_22),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_50),
.A2(n_14),
.B1(n_16),
.B2(n_19),
.Y(n_64)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

AOI21x1_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_62),
.B(n_66),
.Y(n_69)
);

AOI31xp33_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_59),
.A3(n_63),
.B(n_62),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_60),
.C(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_72),
.Y(n_73)
);


endmodule