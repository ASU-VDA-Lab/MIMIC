module fake_netlist_1_7957_n_1272 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_1272);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1272;
wire n_963;
wire n_1034;
wire n_949;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_613;
wire n_648;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_619;
wire n_268;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_271;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_265;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_409;
wire n_315;
wire n_295;
wire n_677;
wire n_1242;
wire n_283;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_272;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_281;
wire n_451;
wire n_487;
wire n_748;
wire n_258;
wire n_253;
wire n_266;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_280;
wire n_395;
wire n_257;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_252;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_275;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_267;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_287;
wire n_606;
wire n_332;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_366;
wire n_596;
wire n_1215;
wire n_286;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_282;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_427;
wire n_703;
wire n_415;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_270;
wire n_1178;
wire n_259;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_254;
wire n_549;
wire n_832;
wire n_996;
wire n_285;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_260;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_956;
wire n_264;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_385;
wire n_1127;
wire n_269;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_288;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1204;
wire n_1094;
wire n_392;
wire n_1169;
wire n_975;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_255;
wire n_844;
wire n_1160;
wire n_274;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_256;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_262;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_276;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_948;
wire n_717;
wire n_861;
wire n_654;
wire n_263;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_335;
wire n_700;
wire n_534;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1219;
wire n_1120;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_261;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
INVx1_ASAP7_75t_L g252 ( .A(n_230), .Y(n_252) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_222), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_113), .Y(n_254) );
CKINVDCx16_ASAP7_75t_R g255 ( .A(n_101), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_6), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_199), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_99), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_185), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_160), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_141), .Y(n_261) );
CKINVDCx16_ASAP7_75t_R g262 ( .A(n_154), .Y(n_262) );
INVxp33_ASAP7_75t_SL g263 ( .A(n_2), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_66), .Y(n_264) );
CKINVDCx16_ASAP7_75t_R g265 ( .A(n_228), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_202), .Y(n_266) );
CKINVDCx16_ASAP7_75t_R g267 ( .A(n_55), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_117), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_26), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_81), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_22), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_84), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_153), .Y(n_273) );
INVxp67_ASAP7_75t_L g274 ( .A(n_59), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_197), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_167), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_48), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_234), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_208), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_24), .Y(n_280) );
BUFx10_ASAP7_75t_L g281 ( .A(n_90), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_238), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_150), .Y(n_283) );
BUFx2_ASAP7_75t_L g284 ( .A(n_170), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_2), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_107), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_30), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_53), .Y(n_288) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_184), .Y(n_289) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_82), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_158), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_112), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_98), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_147), .Y(n_294) );
CKINVDCx20_ASAP7_75t_R g295 ( .A(n_249), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_250), .Y(n_296) );
INVxp33_ASAP7_75t_L g297 ( .A(n_166), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_63), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_244), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_31), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_40), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_155), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_129), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_236), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_28), .Y(n_305) );
CKINVDCx20_ASAP7_75t_R g306 ( .A(n_119), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_135), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_188), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_189), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_140), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_39), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_191), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_67), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_148), .Y(n_314) );
BUFx3_ASAP7_75t_L g315 ( .A(n_181), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_88), .Y(n_316) );
INVxp33_ASAP7_75t_L g317 ( .A(n_137), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_221), .Y(n_318) );
BUFx2_ASAP7_75t_L g319 ( .A(n_10), .Y(n_319) );
INVxp33_ASAP7_75t_SL g320 ( .A(n_33), .Y(n_320) );
CKINVDCx20_ASAP7_75t_R g321 ( .A(n_65), .Y(n_321) );
CKINVDCx20_ASAP7_75t_R g322 ( .A(n_97), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_116), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_165), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_173), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_237), .Y(n_326) );
BUFx3_ASAP7_75t_L g327 ( .A(n_59), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_47), .Y(n_328) );
CKINVDCx14_ASAP7_75t_R g329 ( .A(n_20), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_161), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_78), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_27), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_164), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_89), .Y(n_334) );
INVxp67_ASAP7_75t_L g335 ( .A(n_19), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_218), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_1), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_245), .Y(n_338) );
BUFx2_ASAP7_75t_L g339 ( .A(n_247), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_178), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_136), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_111), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_13), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_235), .Y(n_344) );
CKINVDCx20_ASAP7_75t_R g345 ( .A(n_24), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_23), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_152), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_196), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_239), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_5), .Y(n_350) );
BUFx2_ASAP7_75t_L g351 ( .A(n_193), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_157), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_120), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_231), .Y(n_354) );
CKINVDCx20_ASAP7_75t_R g355 ( .A(n_69), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_87), .Y(n_356) );
CKINVDCx20_ASAP7_75t_R g357 ( .A(n_131), .Y(n_357) );
CKINVDCx14_ASAP7_75t_R g358 ( .A(n_83), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_175), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_35), .Y(n_360) );
INVx2_ASAP7_75t_SL g361 ( .A(n_91), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_134), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_226), .Y(n_363) );
INVxp67_ASAP7_75t_SL g364 ( .A(n_10), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_40), .Y(n_365) );
BUFx5_ASAP7_75t_L g366 ( .A(n_162), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_8), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_106), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_174), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_182), .B(n_33), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_95), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_118), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_64), .Y(n_373) );
CKINVDCx16_ASAP7_75t_R g374 ( .A(n_151), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_172), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_47), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_104), .B(n_121), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_69), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_215), .Y(n_379) );
INVx1_ASAP7_75t_SL g380 ( .A(n_192), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_103), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_177), .Y(n_382) );
INVx2_ASAP7_75t_SL g383 ( .A(n_194), .Y(n_383) );
CKINVDCx14_ASAP7_75t_R g384 ( .A(n_31), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_28), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_219), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_183), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_43), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_214), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_138), .Y(n_390) );
CKINVDCx14_ASAP7_75t_R g391 ( .A(n_251), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_280), .Y(n_392) );
OAI21x1_ASAP7_75t_L g393 ( .A1(n_273), .A2(n_80), .B(n_79), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_366), .Y(n_394) );
INVx3_ASAP7_75t_L g395 ( .A(n_281), .Y(n_395) );
INVx4_ASAP7_75t_L g396 ( .A(n_327), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_366), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_297), .B(n_0), .Y(n_398) );
AND2x6_ASAP7_75t_L g399 ( .A(n_315), .B(n_85), .Y(n_399) );
INVx3_ASAP7_75t_L g400 ( .A(n_281), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_284), .B(n_0), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_366), .Y(n_402) );
BUFx3_ASAP7_75t_L g403 ( .A(n_315), .Y(n_403) );
BUFx2_ASAP7_75t_L g404 ( .A(n_329), .Y(n_404) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_276), .Y(n_405) );
NAND2x1p5_ASAP7_75t_L g406 ( .A(n_377), .B(n_339), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_329), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_280), .Y(n_408) );
NOR2xp33_ASAP7_75t_R g409 ( .A(n_358), .B(n_86), .Y(n_409) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_276), .Y(n_410) );
AND2x4_ASAP7_75t_L g411 ( .A(n_351), .B(n_1), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_297), .B(n_3), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_317), .B(n_3), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_317), .B(n_4), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_319), .B(n_4), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_361), .B(n_383), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_366), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_328), .Y(n_418) );
INVx3_ASAP7_75t_L g419 ( .A(n_281), .Y(n_419) );
INVx3_ASAP7_75t_L g420 ( .A(n_327), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_384), .B(n_5), .Y(n_421) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_276), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_328), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_388), .Y(n_424) );
AND2x4_ASAP7_75t_L g425 ( .A(n_388), .B(n_6), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_366), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_273), .B(n_7), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_394), .Y(n_428) );
NAND2xp33_ASAP7_75t_SL g429 ( .A(n_404), .B(n_407), .Y(n_429) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_405), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_394), .Y(n_431) );
NOR2xp33_ASAP7_75t_SL g432 ( .A(n_399), .B(n_255), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_404), .Y(n_433) );
NAND3xp33_ASAP7_75t_L g434 ( .A(n_427), .B(n_258), .C(n_252), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_394), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_394), .Y(n_436) );
NAND2x1p5_ASAP7_75t_L g437 ( .A(n_427), .B(n_259), .Y(n_437) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_405), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_397), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_395), .B(n_253), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_397), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_397), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_397), .Y(n_443) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_405), .Y(n_444) );
INVx5_ASAP7_75t_L g445 ( .A(n_399), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_402), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_395), .B(n_290), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_402), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_402), .Y(n_449) );
INVx2_ASAP7_75t_SL g450 ( .A(n_404), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_427), .A2(n_384), .B1(n_264), .B2(n_271), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_407), .B(n_358), .Y(n_452) );
AND2x6_ASAP7_75t_L g453 ( .A(n_427), .B(n_260), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_395), .B(n_262), .Y(n_454) );
OAI22xp33_ASAP7_75t_L g455 ( .A1(n_406), .A2(n_267), .B1(n_300), .B2(n_365), .Y(n_455) );
BUFx3_ASAP7_75t_L g456 ( .A(n_403), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_395), .B(n_265), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_427), .Y(n_458) );
INVx4_ASAP7_75t_L g459 ( .A(n_399), .Y(n_459) );
INVx4_ASAP7_75t_L g460 ( .A(n_399), .Y(n_460) );
AND2x6_ASAP7_75t_L g461 ( .A(n_427), .B(n_261), .Y(n_461) );
INVx3_ASAP7_75t_L g462 ( .A(n_425), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_402), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_395), .B(n_269), .Y(n_464) );
INVx3_ASAP7_75t_L g465 ( .A(n_425), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_425), .A2(n_277), .B1(n_287), .B2(n_285), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_400), .B(n_374), .Y(n_467) );
BUFx10_ASAP7_75t_L g468 ( .A(n_411), .Y(n_468) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_405), .Y(n_469) );
INVx3_ASAP7_75t_L g470 ( .A(n_425), .Y(n_470) );
AND2x4_ASAP7_75t_L g471 ( .A(n_400), .B(n_298), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_398), .B(n_391), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_400), .B(n_312), .Y(n_473) );
INVx1_ASAP7_75t_SL g474 ( .A(n_421), .Y(n_474) );
INVx3_ASAP7_75t_L g475 ( .A(n_425), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_417), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_440), .A2(n_416), .B(n_393), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_464), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_472), .B(n_400), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_464), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_464), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_472), .B(n_419), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_440), .B(n_419), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g484 ( .A1(n_434), .A2(n_393), .B(n_417), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_453), .A2(n_411), .B1(n_412), .B2(n_398), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_428), .Y(n_486) );
INVxp67_ASAP7_75t_L g487 ( .A(n_433), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_447), .B(n_419), .Y(n_488) );
INVx4_ASAP7_75t_L g489 ( .A(n_468), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_432), .B(n_459), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_447), .B(n_419), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_452), .B(n_419), .Y(n_492) );
NAND2x1p5_ASAP7_75t_L g493 ( .A(n_474), .B(n_421), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_432), .B(n_411), .Y(n_494) );
AND2x6_ASAP7_75t_SL g495 ( .A(n_464), .B(n_415), .Y(n_495) );
NAND2xp33_ASAP7_75t_L g496 ( .A(n_453), .B(n_399), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_452), .B(n_406), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_471), .Y(n_498) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_474), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_450), .B(n_406), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_471), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_459), .B(n_411), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_459), .B(n_411), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_454), .B(n_406), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_471), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_450), .B(n_406), .Y(n_506) );
INVx3_ASAP7_75t_L g507 ( .A(n_462), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_428), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_451), .A2(n_295), .B1(n_322), .B2(n_306), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_462), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_428), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_459), .B(n_411), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_462), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_453), .B(n_398), .Y(n_514) );
NOR2xp67_ASAP7_75t_L g515 ( .A(n_434), .B(n_421), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_457), .B(n_416), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_468), .B(n_415), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_453), .B(n_412), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_429), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_467), .B(n_401), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_473), .A2(n_393), .B(n_417), .Y(n_521) );
NAND2x1_ASAP7_75t_L g522 ( .A(n_453), .B(n_399), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_460), .B(n_413), .Y(n_523) );
BUFx2_ASAP7_75t_L g524 ( .A(n_455), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_453), .B(n_413), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_461), .A2(n_414), .B1(n_425), .B2(n_320), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_461), .B(n_414), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_465), .Y(n_528) );
CKINVDCx14_ASAP7_75t_R g529 ( .A(n_461), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_460), .B(n_417), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_461), .B(n_403), .Y(n_531) );
INVx2_ASAP7_75t_SL g532 ( .A(n_437), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_473), .A2(n_393), .B(n_426), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_465), .Y(n_534) );
HB1xp67_ASAP7_75t_SL g535 ( .A(n_461), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_461), .A2(n_320), .B1(n_263), .B2(n_420), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_465), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_470), .B(n_396), .Y(n_538) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_437), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_470), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_431), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_461), .B(n_403), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_437), .B(n_396), .Y(n_543) );
NAND2x1p5_ASAP7_75t_L g544 ( .A(n_470), .B(n_301), .Y(n_544) );
AOI22x1_ASAP7_75t_L g545 ( .A1(n_460), .A2(n_426), .B1(n_396), .B2(n_420), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_466), .B(n_396), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_458), .B(n_396), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_470), .A2(n_263), .B1(n_420), .B2(n_396), .Y(n_548) );
AOI22xp33_ASAP7_75t_SL g549 ( .A1(n_475), .A2(n_345), .B1(n_355), .B2(n_321), .Y(n_549) );
OAI22xp33_ASAP7_75t_L g550 ( .A1(n_475), .A2(n_345), .B1(n_355), .B2(n_321), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_445), .B(n_426), .Y(n_551) );
INVxp67_ASAP7_75t_SL g552 ( .A(n_476), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_475), .A2(n_420), .B1(n_399), .B2(n_391), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_475), .A2(n_295), .B1(n_322), .B2(n_306), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_458), .B(n_409), .Y(n_555) );
NOR2xp67_ASAP7_75t_L g556 ( .A(n_458), .B(n_392), .Y(n_556) );
BUFx2_ASAP7_75t_L g557 ( .A(n_456), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_435), .A2(n_399), .B1(n_311), .B2(n_313), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_435), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_456), .B(n_254), .Y(n_560) );
OR2x6_ASAP7_75t_L g561 ( .A(n_476), .B(n_274), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_436), .A2(n_352), .B1(n_357), .B2(n_300), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_436), .B(n_254), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_439), .A2(n_318), .B(n_312), .Y(n_564) );
AND2x6_ASAP7_75t_SL g565 ( .A(n_439), .B(n_305), .Y(n_565) );
NOR2xp33_ASAP7_75t_SL g566 ( .A(n_489), .B(n_445), .Y(n_566) );
O2A1O1Ixp33_ASAP7_75t_L g567 ( .A1(n_499), .A2(n_335), .B(n_442), .C(n_441), .Y(n_567) );
O2A1O1Ixp33_ASAP7_75t_L g568 ( .A1(n_497), .A2(n_441), .B(n_443), .C(n_442), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_502), .A2(n_446), .B(n_443), .Y(n_569) );
OAI21x1_ASAP7_75t_L g570 ( .A1(n_521), .A2(n_449), .B(n_448), .Y(n_570) );
O2A1O1Ixp5_ASAP7_75t_L g571 ( .A1(n_490), .A2(n_449), .B(n_448), .C(n_446), .Y(n_571) );
AOI21x1_ASAP7_75t_L g572 ( .A1(n_522), .A2(n_463), .B(n_449), .Y(n_572) );
A2O1A1Ixp33_ASAP7_75t_L g573 ( .A1(n_477), .A2(n_448), .B(n_337), .C(n_346), .Y(n_573) );
NAND3xp33_ASAP7_75t_L g574 ( .A(n_548), .B(n_445), .C(n_350), .Y(n_574) );
O2A1O1Ixp33_ASAP7_75t_L g575 ( .A1(n_524), .A2(n_364), .B(n_360), .C(n_332), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_507), .Y(n_576) );
O2A1O1Ixp5_ASAP7_75t_L g577 ( .A1(n_490), .A2(n_370), .B(n_344), .C(n_349), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_504), .A2(n_357), .B1(n_352), .B2(n_256), .Y(n_578) );
O2A1O1Ixp33_ASAP7_75t_L g579 ( .A1(n_500), .A2(n_373), .B(n_376), .C(n_367), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_517), .B(n_288), .Y(n_580) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_561), .Y(n_581) );
OAI21x1_ASAP7_75t_L g582 ( .A1(n_533), .A2(n_344), .B(n_318), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_478), .Y(n_583) );
AOI21x1_ASAP7_75t_L g584 ( .A1(n_494), .A2(n_268), .B(n_266), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_485), .A2(n_385), .B1(n_408), .B2(n_392), .Y(n_585) );
NOR2xp33_ASAP7_75t_R g586 ( .A(n_529), .B(n_385), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_487), .B(n_343), .Y(n_587) );
OR2x6_ASAP7_75t_L g588 ( .A(n_554), .B(n_378), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_503), .A2(n_275), .B(n_272), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g590 ( .A1(n_503), .A2(n_282), .B(n_279), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_535), .A2(n_408), .B1(n_418), .B2(n_392), .Y(n_591) );
AND2x2_ASAP7_75t_SL g592 ( .A(n_562), .B(n_283), .Y(n_592) );
BUFx2_ASAP7_75t_SL g593 ( .A(n_539), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_480), .Y(n_594) );
AOI21xp5_ASAP7_75t_L g595 ( .A1(n_512), .A2(n_292), .B(n_286), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_481), .Y(n_596) );
NOR2xp33_ASAP7_75t_R g597 ( .A(n_529), .B(n_270), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_512), .A2(n_296), .B(n_294), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_483), .B(n_270), .Y(n_599) );
AOI33xp33_ASAP7_75t_L g600 ( .A1(n_549), .A2(n_424), .A3(n_423), .B1(n_418), .B2(n_408), .B3(n_310), .Y(n_600) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_530), .A2(n_303), .B(n_299), .Y(n_601) );
NAND2xp5_ASAP7_75t_SL g602 ( .A(n_514), .B(n_278), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_518), .B(n_278), .Y(n_603) );
BUFx4f_ASAP7_75t_L g604 ( .A(n_561), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_507), .Y(n_605) );
CKINVDCx8_ASAP7_75t_R g606 ( .A(n_495), .Y(n_606) );
A2O1A1Ixp33_ASAP7_75t_SL g607 ( .A1(n_520), .A2(n_423), .B(n_424), .C(n_418), .Y(n_607) );
INVx6_ASAP7_75t_L g608 ( .A(n_565), .Y(n_608) );
NOR3xp33_ASAP7_75t_L g609 ( .A(n_509), .B(n_424), .C(n_423), .Y(n_609) );
OAI22xp33_ASAP7_75t_L g610 ( .A1(n_550), .A2(n_356), .B1(n_362), .B2(n_302), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_488), .B(n_302), .Y(n_611) );
INVx8_ASAP7_75t_L g612 ( .A(n_561), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_493), .B(n_356), .Y(n_613) );
O2A1O1Ixp33_ASAP7_75t_L g614 ( .A1(n_506), .A2(n_308), .B(n_314), .C(n_307), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_491), .B(n_362), .Y(n_615) );
O2A1O1Ixp33_ASAP7_75t_SL g616 ( .A1(n_494), .A2(n_326), .B(n_330), .C(n_323), .Y(n_616) );
NOR2xp33_ASAP7_75t_R g617 ( .A(n_519), .B(n_368), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_498), .Y(n_618) );
NOR3xp33_ASAP7_75t_SL g619 ( .A(n_520), .B(n_369), .C(n_368), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_493), .A2(n_333), .B1(n_334), .B2(n_331), .Y(n_620) );
AO32x1_ASAP7_75t_L g621 ( .A1(n_501), .A2(n_372), .A3(n_336), .B1(n_338), .B2(n_340), .Y(n_621) );
INVx3_ASAP7_75t_L g622 ( .A(n_544), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_516), .B(n_371), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_547), .A2(n_342), .B(n_341), .Y(n_624) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_544), .Y(n_625) );
AO32x1_ASAP7_75t_L g626 ( .A1(n_505), .A2(n_382), .A3(n_347), .B1(n_348), .B2(n_354), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_525), .B(n_399), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_526), .A2(n_363), .B1(n_375), .B2(n_353), .Y(n_628) );
OAI21xp33_ASAP7_75t_SL g629 ( .A1(n_552), .A2(n_387), .B(n_386), .Y(n_629) );
NOR2xp33_ASAP7_75t_SL g630 ( .A(n_496), .B(n_399), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_492), .B(n_257), .Y(n_631) );
NOR2xp33_ASAP7_75t_R g632 ( .A(n_519), .B(n_291), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_536), .B(n_7), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_486), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_515), .A2(n_390), .B1(n_389), .B2(n_304), .Y(n_635) );
A2O1A1Ixp33_ASAP7_75t_SL g636 ( .A1(n_484), .A2(n_359), .B(n_381), .C(n_349), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_527), .A2(n_309), .B1(n_316), .B2(n_293), .Y(n_637) );
CKINVDCx6p67_ASAP7_75t_R g638 ( .A(n_479), .Y(n_638) );
INVx3_ASAP7_75t_L g639 ( .A(n_559), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_556), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_482), .B(n_324), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_563), .B(n_523), .Y(n_642) );
OR2x2_ASAP7_75t_SL g643 ( .A(n_543), .B(n_359), .Y(n_643) );
AOI21xp5_ASAP7_75t_L g644 ( .A1(n_523), .A2(n_381), .B(n_380), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_486), .B(n_8), .Y(n_645) );
NOR2x1_ASAP7_75t_SL g646 ( .A(n_531), .B(n_276), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_508), .B(n_325), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_555), .B(n_379), .Y(n_648) );
INVx2_ASAP7_75t_SL g649 ( .A(n_560), .Y(n_649) );
INVx2_ASAP7_75t_SL g650 ( .A(n_511), .Y(n_650) );
OAI21x1_ASAP7_75t_L g651 ( .A1(n_545), .A2(n_366), .B(n_430), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g652 ( .A1(n_538), .A2(n_438), .B(n_430), .Y(n_652) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_557), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_510), .Y(n_654) );
AO21x1_ASAP7_75t_L g655 ( .A1(n_496), .A2(n_410), .B(n_405), .Y(n_655) );
O2A1O1Ixp33_ASAP7_75t_L g656 ( .A1(n_546), .A2(n_9), .B(n_11), .C(n_12), .Y(n_656) );
A2O1A1Ixp33_ASAP7_75t_SL g657 ( .A1(n_553), .A2(n_422), .B(n_405), .C(n_410), .Y(n_657) );
BUFx3_ASAP7_75t_L g658 ( .A(n_541), .Y(n_658) );
A2O1A1Ixp33_ASAP7_75t_L g659 ( .A1(n_513), .A2(n_289), .B(n_422), .C(n_410), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_528), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_534), .Y(n_661) );
INVxp67_ASAP7_75t_L g662 ( .A(n_542), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_537), .B(n_12), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_540), .B(n_13), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_564), .B(n_14), .Y(n_665) );
INVx3_ASAP7_75t_L g666 ( .A(n_558), .Y(n_666) );
NOR2x1_ASAP7_75t_SL g667 ( .A(n_551), .B(n_289), .Y(n_667) );
INVx5_ASAP7_75t_L g668 ( .A(n_561), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_554), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_507), .Y(n_670) );
BUFx6f_ASAP7_75t_L g671 ( .A(n_532), .Y(n_671) );
BUFx12f_ASAP7_75t_L g672 ( .A(n_565), .Y(n_672) );
BUFx8_ASAP7_75t_L g673 ( .A(n_524), .Y(n_673) );
NAND3xp33_ASAP7_75t_L g674 ( .A(n_477), .B(n_410), .C(n_405), .Y(n_674) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_532), .Y(n_675) );
OAI22x1_ASAP7_75t_L g676 ( .A1(n_562), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_504), .A2(n_422), .B1(n_410), .B2(n_438), .Y(n_677) );
A2O1A1Ixp33_ASAP7_75t_L g678 ( .A1(n_477), .A2(n_422), .B(n_410), .C(n_469), .Y(n_678) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_499), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_507), .Y(n_680) );
BUFx2_ASAP7_75t_L g681 ( .A(n_499), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_487), .B(n_15), .Y(n_682) );
NAND3xp33_ASAP7_75t_SL g683 ( .A(n_519), .B(n_16), .C(n_17), .Y(n_683) );
A2O1A1Ixp33_ASAP7_75t_L g684 ( .A1(n_477), .A2(n_422), .B(n_410), .C(n_469), .Y(n_684) );
NAND3xp33_ASAP7_75t_SL g685 ( .A(n_519), .B(n_17), .C(n_18), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_487), .B(n_18), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_478), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_478), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_478), .Y(n_689) );
NOR2xp33_ASAP7_75t_SL g690 ( .A(n_604), .B(n_19), .Y(n_690) );
NOR2xp33_ASAP7_75t_SL g691 ( .A(n_604), .B(n_20), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_679), .Y(n_692) );
AO31x2_ASAP7_75t_L g693 ( .A1(n_573), .A2(n_410), .A3(n_422), .B(n_25), .Y(n_693) );
BUFx3_ASAP7_75t_L g694 ( .A(n_612), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_592), .A2(n_422), .B1(n_410), .B2(n_469), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_585), .A2(n_422), .B1(n_22), .B2(n_25), .Y(n_696) );
OAI22x1_ASAP7_75t_L g697 ( .A1(n_578), .A2(n_21), .B1(n_26), .B2(n_27), .Y(n_697) );
NAND3x1_ASAP7_75t_L g698 ( .A(n_600), .B(n_21), .C(n_29), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_663), .Y(n_699) );
A2O1A1Ixp33_ASAP7_75t_L g700 ( .A1(n_665), .A2(n_444), .B(n_30), .C(n_32), .Y(n_700) );
BUFx6f_ASAP7_75t_L g701 ( .A(n_671), .Y(n_701) );
OR2x2_ASAP7_75t_L g702 ( .A(n_681), .B(n_29), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_581), .B(n_32), .Y(n_703) );
AOI21xp33_ASAP7_75t_L g704 ( .A1(n_567), .A2(n_34), .B(n_35), .Y(n_704) );
AO32x2_ASAP7_75t_L g705 ( .A1(n_620), .A2(n_34), .A3(n_36), .B1(n_37), .B2(n_38), .Y(n_705) );
A2O1A1Ixp33_ASAP7_75t_L g706 ( .A1(n_614), .A2(n_444), .B(n_37), .C(n_38), .Y(n_706) );
O2A1O1Ixp33_ASAP7_75t_L g707 ( .A1(n_579), .A2(n_36), .B(n_39), .C(n_41), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_575), .A2(n_444), .B1(n_42), .B2(n_43), .C(n_44), .Y(n_708) );
BUFx8_ASAP7_75t_L g709 ( .A(n_672), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_583), .Y(n_710) );
AOI21xp5_ASAP7_75t_SL g711 ( .A1(n_591), .A2(n_93), .B(n_92), .Y(n_711) );
A2O1A1Ixp33_ASAP7_75t_L g712 ( .A1(n_629), .A2(n_41), .B(n_42), .C(n_44), .Y(n_712) );
NAND2xp5_ASAP7_75t_SL g713 ( .A(n_668), .B(n_671), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_594), .Y(n_714) );
OAI21x1_ASAP7_75t_L g715 ( .A1(n_570), .A2(n_96), .B(n_94), .Y(n_715) );
NOR2x1_ASAP7_75t_R g716 ( .A(n_668), .B(n_608), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_658), .Y(n_717) );
BUFx2_ASAP7_75t_L g718 ( .A(n_612), .Y(n_718) );
AO21x1_ASAP7_75t_L g719 ( .A1(n_656), .A2(n_102), .B(n_100), .Y(n_719) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_668), .Y(n_720) );
INVx1_ASAP7_75t_SL g721 ( .A(n_593), .Y(n_721) );
BUFx8_ASAP7_75t_L g722 ( .A(n_671), .Y(n_722) );
OAI22xp33_ASAP7_75t_L g723 ( .A1(n_588), .A2(n_45), .B1(n_46), .B2(n_48), .Y(n_723) );
AOI21x1_ASAP7_75t_L g724 ( .A1(n_674), .A2(n_159), .B(n_246), .Y(n_724) );
AO31x2_ASAP7_75t_L g725 ( .A1(n_678), .A2(n_45), .A3(n_46), .B(n_49), .Y(n_725) );
BUFx2_ASAP7_75t_SL g726 ( .A(n_625), .Y(n_726) );
AO31x2_ASAP7_75t_L g727 ( .A1(n_684), .A2(n_49), .A3(n_50), .B(n_51), .Y(n_727) );
OR2x6_ASAP7_75t_L g728 ( .A(n_612), .B(n_50), .Y(n_728) );
AO31x2_ASAP7_75t_L g729 ( .A1(n_655), .A2(n_51), .A3(n_52), .B(n_53), .Y(n_729) );
OAI21x1_ASAP7_75t_L g730 ( .A1(n_582), .A2(n_651), .B(n_674), .Y(n_730) );
OAI221xp5_ASAP7_75t_L g731 ( .A1(n_588), .A2(n_52), .B1(n_54), .B2(n_55), .C(n_56), .Y(n_731) );
OAI21xp5_ASAP7_75t_L g732 ( .A1(n_569), .A2(n_168), .B(n_243), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_634), .Y(n_733) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_669), .B(n_54), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_585), .B(n_57), .Y(n_735) );
A2O1A1Ixp33_ASAP7_75t_L g736 ( .A1(n_568), .A2(n_57), .B(n_58), .C(n_60), .Y(n_736) );
CKINVDCx11_ASAP7_75t_R g737 ( .A(n_606), .Y(n_737) );
AOI22xp5_ASAP7_75t_L g738 ( .A1(n_588), .A2(n_58), .B1(n_60), .B2(n_61), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g739 ( .A1(n_627), .A2(n_169), .B(n_242), .Y(n_739) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_653), .Y(n_740) );
INVx3_ASAP7_75t_L g741 ( .A(n_675), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_613), .B(n_62), .Y(n_742) );
AO21x1_ASAP7_75t_L g743 ( .A1(n_630), .A2(n_171), .B(n_241), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_596), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g745 ( .A1(n_642), .A2(n_163), .B(n_240), .Y(n_745) );
OAI22xp33_ASAP7_75t_L g746 ( .A1(n_608), .A2(n_62), .B1(n_63), .B2(n_64), .Y(n_746) );
NAND3xp33_ASAP7_75t_L g747 ( .A(n_619), .B(n_65), .C(n_66), .Y(n_747) );
BUFx6f_ASAP7_75t_L g748 ( .A(n_675), .Y(n_748) );
BUFx3_ASAP7_75t_L g749 ( .A(n_638), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_609), .B(n_67), .Y(n_750) );
OAI21x1_ASAP7_75t_L g751 ( .A1(n_571), .A2(n_176), .B(n_233), .Y(n_751) );
A2O1A1Ixp33_ASAP7_75t_L g752 ( .A1(n_624), .A2(n_68), .B(n_70), .C(n_71), .Y(n_752) );
OAI21x1_ASAP7_75t_L g753 ( .A1(n_572), .A2(n_156), .B(n_232), .Y(n_753) );
A2O1A1Ixp33_ASAP7_75t_L g754 ( .A1(n_589), .A2(n_68), .B(n_71), .C(n_72), .Y(n_754) );
AO32x2_ASAP7_75t_L g755 ( .A1(n_620), .A2(n_72), .A3(n_73), .B1(n_74), .B2(n_75), .Y(n_755) );
INVx2_ASAP7_75t_SL g756 ( .A(n_586), .Y(n_756) );
OAI21xp5_ASAP7_75t_L g757 ( .A1(n_577), .A2(n_180), .B(n_229), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_639), .Y(n_758) );
INVx2_ASAP7_75t_L g759 ( .A(n_639), .Y(n_759) );
OAI21x1_ASAP7_75t_L g760 ( .A1(n_584), .A2(n_179), .B(n_227), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_622), .B(n_73), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_623), .B(n_75), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_618), .Y(n_763) );
OR2x6_ASAP7_75t_L g764 ( .A(n_676), .B(n_76), .Y(n_764) );
A2O1A1Ixp33_ASAP7_75t_L g765 ( .A1(n_590), .A2(n_76), .B(n_77), .C(n_105), .Y(n_765) );
AND2x2_ASAP7_75t_L g766 ( .A(n_587), .B(n_77), .Y(n_766) );
BUFx5_ASAP7_75t_L g767 ( .A(n_654), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_687), .Y(n_768) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_617), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_580), .B(n_108), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_591), .A2(n_109), .B1(n_110), .B2(n_114), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_688), .Y(n_772) );
CKINVDCx6p67_ASAP7_75t_R g773 ( .A(n_633), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_628), .B(n_115), .Y(n_774) );
AO32x2_ASAP7_75t_L g775 ( .A1(n_621), .A2(n_122), .A3(n_123), .B1(n_124), .B2(n_125), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_645), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_689), .Y(n_777) );
O2A1O1Ixp33_ASAP7_75t_L g778 ( .A1(n_610), .A2(n_126), .B(n_127), .C(n_128), .Y(n_778) );
BUFx3_ASAP7_75t_L g779 ( .A(n_673), .Y(n_779) );
CKINVDCx16_ASAP7_75t_R g780 ( .A(n_632), .Y(n_780) );
BUFx3_ASAP7_75t_L g781 ( .A(n_673), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_664), .Y(n_782) );
A2O1A1Ixp33_ASAP7_75t_L g783 ( .A1(n_595), .A2(n_130), .B(n_132), .C(n_133), .Y(n_783) );
INVx2_ASAP7_75t_L g784 ( .A(n_650), .Y(n_784) );
OAI21xp5_ASAP7_75t_L g785 ( .A1(n_598), .A2(n_139), .B(n_142), .Y(n_785) );
AND2x2_ASAP7_75t_L g786 ( .A(n_682), .B(n_143), .Y(n_786) );
NOR2xp33_ASAP7_75t_SL g787 ( .A(n_630), .B(n_144), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_686), .A2(n_145), .B1(n_146), .B2(n_149), .Y(n_788) );
INVxp67_ASAP7_75t_SL g789 ( .A(n_662), .Y(n_789) );
BUFx3_ASAP7_75t_L g790 ( .A(n_640), .Y(n_790) );
AO31x2_ASAP7_75t_L g791 ( .A1(n_659), .A2(n_186), .A3(n_187), .B(n_190), .Y(n_791) );
AOI21xp5_ASAP7_75t_L g792 ( .A1(n_647), .A2(n_195), .B(n_198), .Y(n_792) );
OAI21xp5_ASAP7_75t_L g793 ( .A1(n_574), .A2(n_200), .B(n_201), .Y(n_793) );
O2A1O1Ixp33_ASAP7_75t_L g794 ( .A1(n_683), .A2(n_203), .B(n_204), .C(n_205), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_643), .A2(n_206), .B1(n_207), .B2(n_209), .Y(n_795) );
A2O1A1Ixp33_ASAP7_75t_L g796 ( .A1(n_644), .A2(n_210), .B(n_211), .C(n_212), .Y(n_796) );
AND2x6_ASAP7_75t_L g797 ( .A(n_660), .B(n_213), .Y(n_797) );
AO31x2_ASAP7_75t_L g798 ( .A1(n_646), .A2(n_216), .A3(n_217), .B(n_220), .Y(n_798) );
AND2x2_ASAP7_75t_SL g799 ( .A(n_597), .B(n_223), .Y(n_799) );
OAI21x1_ASAP7_75t_L g800 ( .A1(n_677), .A2(n_248), .B(n_224), .Y(n_800) );
AO31x2_ASAP7_75t_L g801 ( .A1(n_667), .A2(n_225), .A3(n_661), .B(n_601), .Y(n_801) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_649), .Y(n_802) );
AOI22xp33_ASAP7_75t_SL g803 ( .A1(n_599), .A2(n_611), .B1(n_615), .B2(n_666), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_635), .B(n_666), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_631), .B(n_641), .Y(n_805) );
O2A1O1Ixp33_ASAP7_75t_L g806 ( .A1(n_685), .A2(n_616), .B(n_603), .C(n_602), .Y(n_806) );
INVx2_ASAP7_75t_L g807 ( .A(n_576), .Y(n_807) );
AO22x2_ASAP7_75t_L g808 ( .A1(n_621), .A2(n_626), .B1(n_574), .B2(n_605), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g809 ( .A(n_637), .B(n_648), .Y(n_809) );
HB1xp67_ASAP7_75t_L g810 ( .A(n_670), .Y(n_810) );
CKINVDCx11_ASAP7_75t_R g811 ( .A(n_680), .Y(n_811) );
INVx2_ASAP7_75t_SL g812 ( .A(n_566), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_621), .B(n_626), .Y(n_813) );
INVx2_ASAP7_75t_SL g814 ( .A(n_626), .Y(n_814) );
OAI21x1_ASAP7_75t_L g815 ( .A1(n_570), .A2(n_582), .B(n_651), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_679), .Y(n_816) );
AOI21xp5_ASAP7_75t_L g817 ( .A1(n_652), .A2(n_494), .B(n_490), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_592), .A2(n_524), .B1(n_588), .B2(n_585), .Y(n_818) );
AO31x2_ASAP7_75t_L g819 ( .A1(n_573), .A2(n_678), .A3(n_684), .B(n_655), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_679), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_679), .Y(n_821) );
INVx3_ASAP7_75t_L g822 ( .A(n_671), .Y(n_822) );
O2A1O1Ixp33_ASAP7_75t_SL g823 ( .A1(n_573), .A2(n_607), .B(n_636), .C(n_657), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_625), .B(n_499), .Y(n_824) );
CKINVDCx20_ASAP7_75t_R g825 ( .A(n_617), .Y(n_825) );
OR2x2_ASAP7_75t_L g826 ( .A(n_681), .B(n_554), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_733), .Y(n_827) );
AO31x2_ASAP7_75t_L g828 ( .A1(n_813), .A2(n_719), .A3(n_743), .B(n_817), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_818), .A2(n_773), .B1(n_809), .B2(n_799), .Y(n_829) );
A2O1A1Ixp33_ASAP7_75t_L g830 ( .A1(n_805), .A2(n_803), .B(n_707), .C(n_806), .Y(n_830) );
OAI211xp5_ASAP7_75t_L g831 ( .A1(n_738), .A2(n_695), .B(n_731), .C(n_742), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_692), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_816), .Y(n_833) );
AOI21xp33_ASAP7_75t_L g834 ( .A1(n_778), .A2(n_794), .B(n_804), .Y(n_834) );
AOI22xp33_ASAP7_75t_SL g835 ( .A1(n_690), .A2(n_691), .B1(n_728), .B2(n_734), .Y(n_835) );
OAI21xp5_ASAP7_75t_L g836 ( .A1(n_814), .A2(n_698), .B(n_735), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_764), .A2(n_766), .B1(n_782), .B2(n_826), .Y(n_837) );
HB1xp67_ASAP7_75t_L g838 ( .A(n_824), .Y(n_838) );
OA21x2_ASAP7_75t_L g839 ( .A1(n_757), .A2(n_715), .B(n_753), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_710), .Y(n_840) );
AND2x2_ASAP7_75t_L g841 ( .A(n_802), .B(n_726), .Y(n_841) );
NOR2x1_ASAP7_75t_SL g842 ( .A(n_728), .B(n_701), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_714), .B(n_744), .Y(n_843) );
AOI21xp33_ASAP7_75t_L g844 ( .A1(n_750), .A2(n_762), .B(n_808), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_820), .Y(n_845) );
NAND2x1p5_ASAP7_75t_L g846 ( .A(n_721), .B(n_701), .Y(n_846) );
AO21x2_ASAP7_75t_L g847 ( .A1(n_793), .A2(n_724), .B(n_732), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_821), .Y(n_848) );
OA21x2_ASAP7_75t_L g849 ( .A1(n_751), .A2(n_800), .B(n_760), .Y(n_849) );
NOR2xp33_ASAP7_75t_L g850 ( .A(n_740), .B(n_756), .Y(n_850) );
AND2x4_ASAP7_75t_L g851 ( .A(n_789), .B(n_749), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_763), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_768), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_772), .Y(n_854) );
INVx2_ASAP7_75t_L g855 ( .A(n_777), .Y(n_855) );
AO21x2_ASAP7_75t_L g856 ( .A1(n_785), .A2(n_706), .B(n_700), .Y(n_856) );
HB1xp67_ASAP7_75t_L g857 ( .A(n_722), .Y(n_857) );
CKINVDCx14_ASAP7_75t_R g858 ( .A(n_737), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_761), .Y(n_859) );
NOR2xp33_ASAP7_75t_L g860 ( .A(n_769), .B(n_718), .Y(n_860) );
AOI21xp5_ASAP7_75t_L g861 ( .A1(n_787), .A2(n_812), .B(n_792), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_776), .B(n_699), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_767), .B(n_770), .Y(n_863) );
BUFx6f_ASAP7_75t_L g864 ( .A(n_701), .Y(n_864) );
BUFx6f_ASAP7_75t_L g865 ( .A(n_748), .Y(n_865) );
NOR2xp33_ASAP7_75t_L g866 ( .A(n_694), .B(n_702), .Y(n_866) );
OR2x2_ASAP7_75t_L g867 ( .A(n_780), .B(n_720), .Y(n_867) );
OA21x2_ASAP7_75t_L g868 ( .A1(n_796), .A2(n_745), .B(n_739), .Y(n_868) );
OAI21xp5_ASAP7_75t_L g869 ( .A1(n_696), .A2(n_736), .B(n_712), .Y(n_869) );
NAND2x1p5_ASAP7_75t_L g870 ( .A(n_748), .B(n_741), .Y(n_870) );
AOI22xp5_ASAP7_75t_L g871 ( .A1(n_825), .A2(n_703), .B1(n_764), .B2(n_811), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_767), .B(n_758), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_767), .B(n_759), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_697), .Y(n_874) );
OA21x2_ASAP7_75t_L g875 ( .A1(n_783), .A2(n_765), .B(n_752), .Y(n_875) );
NOR2x1p5_ASAP7_75t_L g876 ( .A(n_779), .B(n_781), .Y(n_876) );
AOI21xp5_ASAP7_75t_L g877 ( .A1(n_774), .A2(n_711), .B(n_786), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_767), .B(n_807), .Y(n_878) );
A2O1A1Ixp33_ASAP7_75t_L g879 ( .A1(n_704), .A2(n_747), .B(n_708), .C(n_754), .Y(n_879) );
OAI21xp5_ASAP7_75t_L g880 ( .A1(n_771), .A2(n_795), .B(n_788), .Y(n_880) );
OAI21x1_ASAP7_75t_L g881 ( .A1(n_822), .A2(n_713), .B(n_717), .Y(n_881) );
CKINVDCx5p33_ASAP7_75t_R g882 ( .A(n_709), .Y(n_882) );
BUFx3_ASAP7_75t_L g883 ( .A(n_722), .Y(n_883) );
OAI221xp5_ASAP7_75t_SL g884 ( .A1(n_723), .A2(n_746), .B1(n_790), .B2(n_716), .C(n_784), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_705), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_810), .B(n_819), .Y(n_886) );
OAI21xp5_ASAP7_75t_L g887 ( .A1(n_797), .A2(n_819), .B(n_693), .Y(n_887) );
A2O1A1Ixp33_ASAP7_75t_L g888 ( .A1(n_748), .A2(n_797), .B(n_705), .C(n_755), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_693), .B(n_797), .Y(n_889) );
AO21x2_ASAP7_75t_L g890 ( .A1(n_775), .A2(n_725), .B(n_727), .Y(n_890) );
AOI321xp33_ASAP7_75t_L g891 ( .A1(n_705), .A2(n_755), .A3(n_727), .B1(n_729), .B2(n_775), .C(n_709), .Y(n_891) );
AOI21xp5_ASAP7_75t_L g892 ( .A1(n_801), .A2(n_775), .B(n_791), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_755), .Y(n_893) );
NOR2x1_ASAP7_75t_R g894 ( .A(n_727), .B(n_729), .Y(n_894) );
AND2x2_ASAP7_75t_L g895 ( .A(n_729), .B(n_791), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_801), .B(n_798), .Y(n_896) );
OA21x2_ASAP7_75t_L g897 ( .A1(n_798), .A2(n_815), .B(n_730), .Y(n_897) );
AO31x2_ASAP7_75t_L g898 ( .A1(n_798), .A2(n_813), .A3(n_678), .B(n_684), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_692), .Y(n_899) );
NAND2xp5_ASAP7_75t_SL g900 ( .A(n_799), .B(n_604), .Y(n_900) );
OA21x2_ASAP7_75t_L g901 ( .A1(n_815), .A2(n_730), .B(n_582), .Y(n_901) );
INVx2_ASAP7_75t_L g902 ( .A(n_733), .Y(n_902) );
INVx2_ASAP7_75t_SL g903 ( .A(n_722), .Y(n_903) );
AO31x2_ASAP7_75t_L g904 ( .A1(n_813), .A2(n_678), .A3(n_684), .B(n_719), .Y(n_904) );
AO21x2_ASAP7_75t_L g905 ( .A1(n_813), .A2(n_684), .B(n_678), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_818), .A2(n_592), .B1(n_524), .B2(n_673), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_692), .Y(n_907) );
AOI221xp5_ASAP7_75t_L g908 ( .A1(n_818), .A2(n_455), .B1(n_585), .B2(n_550), .C(n_575), .Y(n_908) );
O2A1O1Ixp33_ASAP7_75t_L g909 ( .A1(n_805), .A2(n_455), .B(n_742), .C(n_712), .Y(n_909) );
AO21x2_ASAP7_75t_L g910 ( .A1(n_813), .A2(n_684), .B(n_678), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_692), .Y(n_911) );
INVx2_ASAP7_75t_L g912 ( .A(n_733), .Y(n_912) );
AND2x2_ASAP7_75t_L g913 ( .A(n_818), .B(n_681), .Y(n_913) );
AND2x4_ASAP7_75t_L g914 ( .A(n_789), .B(n_622), .Y(n_914) );
NOR2x1_ASAP7_75t_R g915 ( .A(n_737), .B(n_672), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_710), .B(n_714), .Y(n_916) );
INVx2_ASAP7_75t_SL g917 ( .A(n_722), .Y(n_917) );
INVx3_ASAP7_75t_SL g918 ( .A(n_721), .Y(n_918) );
AND2x4_ASAP7_75t_SL g919 ( .A(n_728), .B(n_625), .Y(n_919) );
CKINVDCx5p33_ASAP7_75t_R g920 ( .A(n_737), .Y(n_920) );
INVx2_ASAP7_75t_L g921 ( .A(n_733), .Y(n_921) );
OAI21xp5_ASAP7_75t_L g922 ( .A1(n_813), .A2(n_573), .B(n_477), .Y(n_922) );
BUFx3_ASAP7_75t_L g923 ( .A(n_722), .Y(n_923) );
OR2x2_ASAP7_75t_L g924 ( .A(n_826), .B(n_554), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_710), .B(n_714), .Y(n_925) );
OAI22xp5_ASAP7_75t_L g926 ( .A1(n_818), .A2(n_585), .B1(n_735), .B2(n_799), .Y(n_926) );
NOR2xp67_ASAP7_75t_SL g927 ( .A(n_780), .B(n_668), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_692), .Y(n_928) );
NOR2xp33_ASAP7_75t_L g929 ( .A(n_773), .B(n_524), .Y(n_929) );
INVx2_ASAP7_75t_L g930 ( .A(n_733), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_692), .Y(n_931) );
BUFx3_ASAP7_75t_L g932 ( .A(n_722), .Y(n_932) );
BUFx8_ASAP7_75t_L g933 ( .A(n_779), .Y(n_933) );
INVx3_ASAP7_75t_L g934 ( .A(n_722), .Y(n_934) );
OAI22xp33_ASAP7_75t_L g935 ( .A1(n_690), .A2(n_554), .B1(n_588), .B2(n_604), .Y(n_935) );
INVx1_ASAP7_75t_L g936 ( .A(n_692), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_692), .Y(n_937) );
INVx4_ASAP7_75t_L g938 ( .A(n_728), .Y(n_938) );
AOI21xp5_ASAP7_75t_L g939 ( .A1(n_823), .A2(n_674), .B(n_678), .Y(n_939) );
AND2x2_ASAP7_75t_L g940 ( .A(n_818), .B(n_681), .Y(n_940) );
AOI21xp5_ASAP7_75t_L g941 ( .A1(n_823), .A2(n_674), .B(n_678), .Y(n_941) );
AND2x2_ASAP7_75t_L g942 ( .A(n_818), .B(n_681), .Y(n_942) );
INVx2_ASAP7_75t_L g943 ( .A(n_733), .Y(n_943) );
HB1xp67_ASAP7_75t_L g944 ( .A(n_838), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_926), .A2(n_906), .B1(n_908), .B2(n_829), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_886), .Y(n_946) );
INVx1_ASAP7_75t_L g947 ( .A(n_885), .Y(n_947) );
CKINVDCx11_ASAP7_75t_R g948 ( .A(n_883), .Y(n_948) );
AND2x2_ASAP7_75t_L g949 ( .A(n_943), .B(n_827), .Y(n_949) );
HB1xp67_ASAP7_75t_L g950 ( .A(n_841), .Y(n_950) );
INVx2_ASAP7_75t_L g951 ( .A(n_905), .Y(n_951) );
AND2x2_ASAP7_75t_L g952 ( .A(n_902), .B(n_912), .Y(n_952) );
OR2x2_ASAP7_75t_L g953 ( .A(n_913), .B(n_942), .Y(n_953) );
OA21x2_ASAP7_75t_L g954 ( .A1(n_892), .A2(n_887), .B(n_896), .Y(n_954) );
INVxp33_ASAP7_75t_L g955 ( .A(n_927), .Y(n_955) );
AND2x2_ASAP7_75t_L g956 ( .A(n_921), .B(n_930), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_926), .A2(n_908), .B1(n_935), .B2(n_900), .Y(n_957) );
BUFx3_ASAP7_75t_L g958 ( .A(n_923), .Y(n_958) );
AND2x2_ASAP7_75t_L g959 ( .A(n_840), .B(n_855), .Y(n_959) );
OR2x2_ASAP7_75t_L g960 ( .A(n_940), .B(n_924), .Y(n_960) );
INVx2_ASAP7_75t_L g961 ( .A(n_910), .Y(n_961) );
HB1xp67_ASAP7_75t_L g962 ( .A(n_914), .Y(n_962) );
A2O1A1Ixp33_ASAP7_75t_L g963 ( .A1(n_909), .A2(n_830), .B(n_884), .C(n_874), .Y(n_963) );
BUFx3_ASAP7_75t_L g964 ( .A(n_932), .Y(n_964) );
AOI322xp5_ASAP7_75t_L g965 ( .A1(n_837), .A2(n_835), .A3(n_929), .B1(n_871), .B2(n_858), .C1(n_852), .C2(n_853), .Y(n_965) );
INVx1_ASAP7_75t_L g966 ( .A(n_893), .Y(n_966) );
NAND2xp5_ASAP7_75t_L g967 ( .A(n_854), .B(n_843), .Y(n_967) );
AOI22xp5_ASAP7_75t_L g968 ( .A1(n_831), .A2(n_938), .B1(n_859), .B2(n_869), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_843), .Y(n_969) );
BUFx3_ASAP7_75t_L g970 ( .A(n_934), .Y(n_970) );
AO21x2_ASAP7_75t_L g971 ( .A1(n_844), .A2(n_889), .B(n_922), .Y(n_971) );
AND2x4_ASAP7_75t_L g972 ( .A(n_872), .B(n_873), .Y(n_972) );
BUFx2_ASAP7_75t_L g973 ( .A(n_864), .Y(n_973) );
BUFx2_ASAP7_75t_L g974 ( .A(n_865), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_916), .Y(n_975) );
AO21x2_ASAP7_75t_L g976 ( .A1(n_922), .A2(n_941), .B(n_939), .Y(n_976) );
INVx3_ASAP7_75t_L g977 ( .A(n_865), .Y(n_977) );
OAI22xp5_ASAP7_75t_L g978 ( .A1(n_938), .A2(n_863), .B1(n_919), .B2(n_888), .Y(n_978) );
OAI22xp5_ASAP7_75t_L g979 ( .A1(n_863), .A2(n_918), .B1(n_916), .B2(n_925), .Y(n_979) );
OAI21xp5_ASAP7_75t_L g980 ( .A1(n_879), .A2(n_869), .B(n_834), .Y(n_980) );
INVx1_ASAP7_75t_L g981 ( .A(n_925), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_894), .Y(n_982) );
INVx2_ASAP7_75t_L g983 ( .A(n_901), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_832), .B(n_833), .Y(n_984) );
AND2x2_ASAP7_75t_L g985 ( .A(n_845), .B(n_848), .Y(n_985) );
OAI21xp33_ASAP7_75t_L g986 ( .A1(n_895), .A2(n_836), .B(n_866), .Y(n_986) );
INVxp67_ASAP7_75t_SL g987 ( .A(n_878), .Y(n_987) );
OR2x6_ASAP7_75t_L g988 ( .A(n_877), .B(n_836), .Y(n_988) );
BUFx2_ASAP7_75t_L g989 ( .A(n_878), .Y(n_989) );
OR2x2_ASAP7_75t_L g990 ( .A(n_862), .B(n_937), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_890), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_891), .Y(n_992) );
INVx1_ASAP7_75t_L g993 ( .A(n_891), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_872), .Y(n_994) );
OR2x6_ASAP7_75t_L g995 ( .A(n_880), .B(n_861), .Y(n_995) );
AND2x2_ASAP7_75t_L g996 ( .A(n_899), .B(n_936), .Y(n_996) );
OR2x6_ASAP7_75t_L g997 ( .A(n_880), .B(n_873), .Y(n_997) );
INVx4_ASAP7_75t_SL g998 ( .A(n_914), .Y(n_998) );
AND2x2_ASAP7_75t_L g999 ( .A(n_907), .B(n_931), .Y(n_999) );
OR2x6_ASAP7_75t_L g1000 ( .A(n_846), .B(n_881), .Y(n_1000) );
OAI22xp5_ASAP7_75t_L g1001 ( .A1(n_851), .A2(n_862), .B1(n_846), .B2(n_911), .Y(n_1001) );
INVx1_ASAP7_75t_L g1002 ( .A(n_928), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_842), .B(n_870), .Y(n_1003) );
OAI22xp5_ASAP7_75t_L g1004 ( .A1(n_851), .A2(n_860), .B1(n_867), .B2(n_850), .Y(n_1004) );
INVx2_ASAP7_75t_SL g1005 ( .A(n_876), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_898), .Y(n_1006) );
AOI322xp5_ASAP7_75t_L g1007 ( .A1(n_857), .A2(n_917), .A3(n_903), .B1(n_934), .B2(n_882), .C1(n_920), .C2(n_915), .Y(n_1007) );
INVx1_ASAP7_75t_L g1008 ( .A(n_898), .Y(n_1008) );
AND2x4_ASAP7_75t_L g1009 ( .A(n_856), .B(n_904), .Y(n_1009) );
INVx2_ASAP7_75t_L g1010 ( .A(n_898), .Y(n_1010) );
HB1xp67_ASAP7_75t_L g1011 ( .A(n_933), .Y(n_1011) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_856), .B(n_875), .Y(n_1012) );
CKINVDCx11_ASAP7_75t_R g1013 ( .A(n_933), .Y(n_1013) );
INVx3_ASAP7_75t_L g1014 ( .A(n_849), .Y(n_1014) );
OA21x2_ASAP7_75t_L g1015 ( .A1(n_828), .A2(n_897), .B(n_904), .Y(n_1015) );
INVx1_ASAP7_75t_L g1016 ( .A(n_828), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_828), .B(n_868), .Y(n_1017) );
NAND2xp33_ASAP7_75t_R g1018 ( .A(n_1003), .B(n_868), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_972), .B(n_847), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_972), .B(n_839), .Y(n_1020) );
INVx4_ASAP7_75t_R g1021 ( .A(n_958), .Y(n_1021) );
AND2x4_ASAP7_75t_L g1022 ( .A(n_982), .B(n_988), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_947), .Y(n_1023) );
INVx1_ASAP7_75t_L g1024 ( .A(n_947), .Y(n_1024) );
NAND2x1_ASAP7_75t_L g1025 ( .A(n_1000), .B(n_988), .Y(n_1025) );
INVxp67_ASAP7_75t_L g1026 ( .A(n_944), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_972), .B(n_992), .Y(n_1027) );
HB1xp67_ASAP7_75t_L g1028 ( .A(n_950), .Y(n_1028) );
AND2x4_ASAP7_75t_L g1029 ( .A(n_982), .B(n_988), .Y(n_1029) );
NOR2xp67_ASAP7_75t_L g1030 ( .A(n_968), .B(n_978), .Y(n_1030) );
OR2x2_ASAP7_75t_L g1031 ( .A(n_953), .B(n_960), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_992), .B(n_993), .Y(n_1032) );
NAND2xp5_ASAP7_75t_L g1033 ( .A(n_984), .B(n_985), .Y(n_1033) );
INVx1_ASAP7_75t_L g1034 ( .A(n_966), .Y(n_1034) );
AND2x4_ASAP7_75t_L g1035 ( .A(n_988), .B(n_997), .Y(n_1035) );
OR2x2_ASAP7_75t_L g1036 ( .A(n_953), .B(n_960), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_966), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_993), .B(n_994), .Y(n_1038) );
NAND2xp5_ASAP7_75t_L g1039 ( .A(n_984), .B(n_985), .Y(n_1039) );
HB1xp67_ASAP7_75t_L g1040 ( .A(n_989), .Y(n_1040) );
NOR2x1_ASAP7_75t_L g1041 ( .A(n_979), .B(n_1001), .Y(n_1041) );
AND2x2_ASAP7_75t_L g1042 ( .A(n_994), .B(n_989), .Y(n_1042) );
INVx2_ASAP7_75t_SL g1043 ( .A(n_998), .Y(n_1043) );
NAND2xp5_ASAP7_75t_L g1044 ( .A(n_996), .B(n_999), .Y(n_1044) );
AND2x4_ASAP7_75t_L g1045 ( .A(n_988), .B(n_997), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_959), .B(n_1012), .Y(n_1046) );
OR2x2_ASAP7_75t_L g1047 ( .A(n_946), .B(n_969), .Y(n_1047) );
AND2x2_ASAP7_75t_L g1048 ( .A(n_959), .B(n_1012), .Y(n_1048) );
HB1xp67_ASAP7_75t_L g1049 ( .A(n_990), .Y(n_1049) );
BUFx2_ASAP7_75t_L g1050 ( .A(n_987), .Y(n_1050) );
OAI22xp5_ASAP7_75t_L g1051 ( .A1(n_957), .A2(n_945), .B1(n_968), .B2(n_963), .Y(n_1051) );
BUFx2_ASAP7_75t_L g1052 ( .A(n_1000), .Y(n_1052) );
HB1xp67_ASAP7_75t_L g1053 ( .A(n_990), .Y(n_1053) );
INVx2_ASAP7_75t_L g1054 ( .A(n_983), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_997), .B(n_949), .Y(n_1055) );
BUFx2_ASAP7_75t_L g1056 ( .A(n_1000), .Y(n_1056) );
AO22x1_ASAP7_75t_L g1057 ( .A1(n_1005), .A2(n_955), .B1(n_1011), .B2(n_981), .Y(n_1057) );
INVx1_ASAP7_75t_SL g1058 ( .A(n_958), .Y(n_1058) );
NAND4xp25_ASAP7_75t_L g1059 ( .A(n_965), .B(n_1007), .C(n_980), .D(n_986), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g1060 ( .A(n_996), .B(n_999), .Y(n_1060) );
AND2x2_ASAP7_75t_L g1061 ( .A(n_997), .B(n_949), .Y(n_1061) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_997), .B(n_952), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_952), .B(n_956), .Y(n_1063) );
HB1xp67_ASAP7_75t_L g1064 ( .A(n_962), .Y(n_1064) );
INVx1_ASAP7_75t_L g1065 ( .A(n_991), .Y(n_1065) );
NAND2xp5_ASAP7_75t_R g1066 ( .A(n_1005), .B(n_1003), .Y(n_1066) );
BUFx2_ASAP7_75t_L g1067 ( .A(n_1000), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_956), .B(n_969), .Y(n_1068) );
AND2x2_ASAP7_75t_SL g1069 ( .A(n_998), .B(n_1009), .Y(n_1069) );
INVx2_ASAP7_75t_SL g1070 ( .A(n_998), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_975), .B(n_981), .Y(n_1071) );
HB1xp67_ASAP7_75t_L g1072 ( .A(n_975), .Y(n_1072) );
INVx4_ASAP7_75t_L g1073 ( .A(n_998), .Y(n_1073) );
HB1xp67_ASAP7_75t_L g1074 ( .A(n_967), .Y(n_1074) );
HB1xp67_ASAP7_75t_L g1075 ( .A(n_1002), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1046), .B(n_1009), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1023), .Y(n_1077) );
AND2x2_ASAP7_75t_L g1078 ( .A(n_1046), .B(n_1009), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_1048), .B(n_1009), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_1048), .B(n_971), .Y(n_1080) );
INVx2_ASAP7_75t_L g1081 ( .A(n_1054), .Y(n_1081) );
INVx1_ASAP7_75t_SL g1082 ( .A(n_1050), .Y(n_1082) );
NAND2xp5_ASAP7_75t_L g1083 ( .A(n_1063), .B(n_1049), .Y(n_1083) );
NAND2xp33_ASAP7_75t_SL g1084 ( .A(n_1073), .B(n_1004), .Y(n_1084) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1023), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_1063), .B(n_1053), .Y(n_1086) );
AND2x2_ASAP7_75t_L g1087 ( .A(n_1055), .B(n_971), .Y(n_1087) );
AND2x2_ASAP7_75t_L g1088 ( .A(n_1055), .B(n_971), .Y(n_1088) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1024), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1024), .Y(n_1090) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1034), .Y(n_1091) );
NAND2xp5_ASAP7_75t_L g1092 ( .A(n_1074), .B(n_1002), .Y(n_1092) );
OR2x2_ASAP7_75t_L g1093 ( .A(n_1031), .B(n_1006), .Y(n_1093) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1034), .Y(n_1094) );
OR2x2_ASAP7_75t_L g1095 ( .A(n_1031), .B(n_1008), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1096 ( .A(n_1061), .B(n_1008), .Y(n_1096) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_1061), .B(n_1017), .Y(n_1097) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1037), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_1059), .A2(n_995), .B1(n_970), .B2(n_964), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_1062), .B(n_1017), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1062), .B(n_1016), .Y(n_1101) );
HB1xp67_ASAP7_75t_L g1102 ( .A(n_1028), .Y(n_1102) );
OR2x2_ASAP7_75t_L g1103 ( .A(n_1036), .B(n_1016), .Y(n_1103) );
BUFx2_ASAP7_75t_L g1104 ( .A(n_1050), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_1019), .B(n_954), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_1019), .B(n_954), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_1027), .B(n_954), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1027), .B(n_954), .Y(n_1108) );
OR2x2_ASAP7_75t_L g1109 ( .A(n_1036), .B(n_1010), .Y(n_1109) );
NOR2xp33_ASAP7_75t_SL g1110 ( .A(n_1073), .B(n_1069), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_1020), .B(n_1015), .Y(n_1111) );
NAND2xp5_ASAP7_75t_L g1112 ( .A(n_1038), .B(n_970), .Y(n_1112) );
OR2x2_ASAP7_75t_L g1113 ( .A(n_1033), .B(n_961), .Y(n_1113) );
INVxp33_ASAP7_75t_L g1114 ( .A(n_1021), .Y(n_1114) );
OR2x2_ASAP7_75t_L g1115 ( .A(n_1039), .B(n_961), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1035), .B(n_1015), .Y(n_1116) );
HB1xp67_ASAP7_75t_L g1117 ( .A(n_1040), .Y(n_1117) );
INVx3_ASAP7_75t_L g1118 ( .A(n_1025), .Y(n_1118) );
NAND5xp2_ASAP7_75t_L g1119 ( .A(n_1021), .B(n_1013), .C(n_948), .D(n_964), .E(n_974), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_1035), .B(n_1015), .Y(n_1120) );
NAND2xp5_ASAP7_75t_L g1121 ( .A(n_1038), .B(n_976), .Y(n_1121) );
AND2x4_ASAP7_75t_L g1122 ( .A(n_1022), .B(n_995), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1065), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1124 ( .A(n_1035), .B(n_1015), .Y(n_1124) );
AND2x4_ASAP7_75t_L g1125 ( .A(n_1022), .B(n_995), .Y(n_1125) );
OR2x2_ASAP7_75t_L g1126 ( .A(n_1044), .B(n_951), .Y(n_1126) );
INVx2_ASAP7_75t_L g1127 ( .A(n_1081), .Y(n_1127) );
NOR2x1_ASAP7_75t_L g1128 ( .A(n_1119), .B(n_1058), .Y(n_1128) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1102), .Y(n_1129) );
NOR2xp33_ASAP7_75t_L g1130 ( .A(n_1112), .B(n_1059), .Y(n_1130) );
AND2x4_ASAP7_75t_L g1131 ( .A(n_1122), .B(n_1022), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1132 ( .A(n_1083), .B(n_1032), .Y(n_1132) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1092), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g1134 ( .A(n_1086), .B(n_1032), .Y(n_1134) );
AND3x2_ASAP7_75t_L g1135 ( .A(n_1110), .B(n_1067), .C(n_1052), .Y(n_1135) );
OR2x6_ASAP7_75t_L g1136 ( .A(n_1118), .B(n_1025), .Y(n_1136) );
OR2x2_ASAP7_75t_L g1137 ( .A(n_1109), .B(n_1093), .Y(n_1137) );
NOR2x1_ASAP7_75t_L g1138 ( .A(n_1119), .B(n_1073), .Y(n_1138) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1077), .Y(n_1139) );
NAND2xp5_ASAP7_75t_L g1140 ( .A(n_1107), .B(n_1108), .Y(n_1140) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1077), .Y(n_1141) );
OR2x2_ASAP7_75t_L g1142 ( .A(n_1109), .B(n_1060), .Y(n_1142) );
OR2x2_ASAP7_75t_L g1143 ( .A(n_1093), .B(n_1075), .Y(n_1143) );
INVx3_ASAP7_75t_SL g1144 ( .A(n_1082), .Y(n_1144) );
OR2x2_ASAP7_75t_L g1145 ( .A(n_1095), .B(n_1072), .Y(n_1145) );
INVx1_ASAP7_75t_SL g1146 ( .A(n_1082), .Y(n_1146) );
HB1xp67_ASAP7_75t_L g1147 ( .A(n_1104), .Y(n_1147) );
NAND2xp5_ASAP7_75t_L g1148 ( .A(n_1107), .B(n_1068), .Y(n_1148) );
OR2x6_ASAP7_75t_L g1149 ( .A(n_1118), .B(n_1073), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1150 ( .A(n_1108), .B(n_1068), .Y(n_1150) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_1105), .B(n_1035), .Y(n_1151) );
NOR2xp33_ASAP7_75t_L g1152 ( .A(n_1117), .B(n_1051), .Y(n_1152) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1085), .Y(n_1153) );
NAND2xp5_ASAP7_75t_L g1154 ( .A(n_1103), .B(n_1071), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1085), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_1097), .B(n_1022), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1103), .B(n_1071), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1089), .Y(n_1158) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_1105), .B(n_1045), .Y(n_1159) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1089), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1106), .B(n_1045), .Y(n_1161) );
INVx3_ASAP7_75t_L g1162 ( .A(n_1118), .Y(n_1162) );
NAND4xp25_ASAP7_75t_L g1163 ( .A(n_1099), .B(n_1041), .C(n_1030), .D(n_1018), .Y(n_1163) );
OR2x2_ASAP7_75t_L g1164 ( .A(n_1095), .B(n_1042), .Y(n_1164) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1090), .Y(n_1165) );
OR2x2_ASAP7_75t_L g1166 ( .A(n_1113), .B(n_1042), .Y(n_1166) );
NOR2xp33_ASAP7_75t_L g1167 ( .A(n_1121), .B(n_1026), .Y(n_1167) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1106), .B(n_1045), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1140), .B(n_1087), .Y(n_1169) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1137), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1151), .B(n_1087), .Y(n_1171) );
NAND2xp5_ASAP7_75t_L g1172 ( .A(n_1133), .B(n_1080), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1139), .Y(n_1173) );
NAND2xp5_ASAP7_75t_L g1174 ( .A(n_1167), .B(n_1080), .Y(n_1174) );
NAND2xp5_ASAP7_75t_L g1175 ( .A(n_1167), .B(n_1088), .Y(n_1175) );
OR2x2_ASAP7_75t_L g1176 ( .A(n_1148), .B(n_1113), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1151), .B(n_1088), .Y(n_1177) );
AND2x4_ASAP7_75t_L g1178 ( .A(n_1136), .B(n_1118), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1141), .Y(n_1179) );
AND2x4_ASAP7_75t_L g1180 ( .A(n_1136), .B(n_1131), .Y(n_1180) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1153), .Y(n_1181) );
INVx2_ASAP7_75t_L g1182 ( .A(n_1127), .Y(n_1182) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1152), .B(n_1096), .Y(n_1183) );
OR2x2_ASAP7_75t_L g1184 ( .A(n_1150), .B(n_1115), .Y(n_1184) );
INVx2_ASAP7_75t_L g1185 ( .A(n_1127), .Y(n_1185) );
HB1xp67_ASAP7_75t_L g1186 ( .A(n_1147), .Y(n_1186) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1166), .Y(n_1187) );
INVx1_ASAP7_75t_SL g1188 ( .A(n_1144), .Y(n_1188) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1155), .Y(n_1189) );
OAI21x1_ASAP7_75t_L g1190 ( .A1(n_1138), .A2(n_1041), .B(n_1014), .Y(n_1190) );
INVxp67_ASAP7_75t_L g1191 ( .A(n_1130), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1129), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1143), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1159), .B(n_1111), .Y(n_1194) );
NAND2xp5_ASAP7_75t_L g1195 ( .A(n_1152), .B(n_1096), .Y(n_1195) );
OR2x2_ASAP7_75t_L g1196 ( .A(n_1164), .B(n_1115), .Y(n_1196) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1158), .Y(n_1197) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1160), .Y(n_1198) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1165), .Y(n_1199) );
AOI22xp5_ASAP7_75t_L g1200 ( .A1(n_1191), .A2(n_1130), .B1(n_1128), .B2(n_1163), .Y(n_1200) );
NAND4xp25_ASAP7_75t_L g1201 ( .A(n_1188), .B(n_1030), .C(n_1084), .D(n_1110), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1196), .Y(n_1202) );
AOI22xp5_ASAP7_75t_L g1203 ( .A1(n_1183), .A2(n_1132), .B1(n_1134), .B2(n_1159), .Y(n_1203) );
AOI22xp5_ASAP7_75t_L g1204 ( .A1(n_1195), .A2(n_1193), .B1(n_1174), .B2(n_1170), .Y(n_1204) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1196), .Y(n_1205) );
NOR2x1_ASAP7_75t_L g1206 ( .A(n_1180), .B(n_1149), .Y(n_1206) );
AOI22xp5_ASAP7_75t_L g1207 ( .A1(n_1172), .A2(n_1168), .B1(n_1161), .B2(n_1131), .Y(n_1207) );
OR2x2_ASAP7_75t_L g1208 ( .A(n_1176), .B(n_1142), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1173), .Y(n_1209) );
OAI322xp33_ASAP7_75t_L g1210 ( .A1(n_1175), .A2(n_1145), .A3(n_1154), .B1(n_1157), .B2(n_1146), .C1(n_1144), .C2(n_1126), .Y(n_1210) );
NOR2xp33_ASAP7_75t_L g1211 ( .A(n_1192), .B(n_1114), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1212 ( .A(n_1169), .B(n_1147), .Y(n_1212) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1173), .Y(n_1213) );
NAND2xp5_ASAP7_75t_L g1214 ( .A(n_1169), .B(n_1161), .Y(n_1214) );
INVx1_ASAP7_75t_SL g1215 ( .A(n_1186), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1194), .B(n_1168), .Y(n_1216) );
NOR2xp33_ASAP7_75t_L g1217 ( .A(n_1187), .B(n_1057), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1194), .B(n_1156), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1179), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1179), .Y(n_1220) );
HB1xp67_ASAP7_75t_L g1221 ( .A(n_1215), .Y(n_1221) );
AOI211xp5_ASAP7_75t_L g1222 ( .A1(n_1210), .A2(n_1057), .B(n_1178), .C(n_1180), .Y(n_1222) );
OAI22xp5_ASAP7_75t_L g1223 ( .A1(n_1200), .A2(n_1180), .B1(n_1176), .B2(n_1184), .Y(n_1223) );
OAI21xp33_ASAP7_75t_SL g1224 ( .A1(n_1206), .A2(n_1149), .B(n_1190), .Y(n_1224) );
AOI22xp5_ASAP7_75t_L g1225 ( .A1(n_1217), .A2(n_1178), .B1(n_1131), .B2(n_1177), .Y(n_1225) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1209), .Y(n_1226) );
O2A1O1Ixp33_ASAP7_75t_L g1227 ( .A1(n_1215), .A2(n_1064), .B(n_1184), .C(n_1199), .Y(n_1227) );
AOI22xp33_ASAP7_75t_SL g1228 ( .A1(n_1211), .A2(n_1178), .B1(n_1104), .B2(n_1069), .Y(n_1228) );
AOI221xp5_ASAP7_75t_L g1229 ( .A1(n_1202), .A2(n_1171), .B1(n_1177), .B2(n_1189), .C(n_1198), .Y(n_1229) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1213), .Y(n_1230) );
OAI21xp5_ASAP7_75t_L g1231 ( .A1(n_1201), .A2(n_1190), .B(n_1149), .Y(n_1231) );
NAND2xp5_ASAP7_75t_L g1232 ( .A(n_1204), .B(n_1171), .Y(n_1232) );
AOI322xp5_ASAP7_75t_L g1233 ( .A1(n_1205), .A2(n_1076), .A3(n_1078), .B1(n_1079), .B2(n_1100), .C1(n_1097), .C2(n_1181), .Y(n_1233) );
AOI221xp5_ASAP7_75t_L g1234 ( .A1(n_1212), .A2(n_1198), .B1(n_1197), .B2(n_1189), .C(n_1181), .Y(n_1234) );
AOI21x1_ASAP7_75t_L g1235 ( .A1(n_1221), .A2(n_1136), .B(n_1216), .Y(n_1235) );
AND2x2_ASAP7_75t_SL g1236 ( .A(n_1224), .B(n_1069), .Y(n_1236) );
OAI222xp33_ASAP7_75t_L g1237 ( .A1(n_1228), .A2(n_1207), .B1(n_1203), .B2(n_1208), .C1(n_1214), .C2(n_1218), .Y(n_1237) );
NOR4xp75_ASAP7_75t_L g1238 ( .A(n_1223), .B(n_1214), .C(n_1043), .D(n_1070), .Y(n_1238) );
AOI221xp5_ASAP7_75t_L g1239 ( .A1(n_1222), .A2(n_1220), .B1(n_1219), .B2(n_1197), .C(n_1101), .Y(n_1239) );
NOR2x1_ASAP7_75t_L g1240 ( .A(n_1227), .B(n_1162), .Y(n_1240) );
OAI21xp5_ASAP7_75t_L g1241 ( .A1(n_1228), .A2(n_1070), .B(n_1043), .Y(n_1241) );
AOI21xp5_ASAP7_75t_L g1242 ( .A1(n_1231), .A2(n_1162), .B(n_1185), .Y(n_1242) );
AOI221xp5_ASAP7_75t_L g1243 ( .A1(n_1229), .A2(n_1101), .B1(n_1116), .B2(n_1120), .C(n_1124), .Y(n_1243) );
NOR2xp33_ASAP7_75t_L g1244 ( .A(n_1232), .B(n_1162), .Y(n_1244) );
NAND4xp25_ASAP7_75t_L g1245 ( .A(n_1239), .B(n_1225), .C(n_1233), .D(n_1234), .Y(n_1245) );
NAND3xp33_ASAP7_75t_SL g1246 ( .A(n_1238), .B(n_1230), .C(n_1226), .Y(n_1246) );
OAI221xp5_ASAP7_75t_L g1247 ( .A1(n_1240), .A2(n_1185), .B1(n_1182), .B2(n_1052), .C(n_1056), .Y(n_1247) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1244), .Y(n_1248) );
NAND3xp33_ASAP7_75t_SL g1249 ( .A(n_1241), .B(n_1066), .C(n_974), .Y(n_1249) );
NAND4xp25_ASAP7_75t_L g1250 ( .A(n_1243), .B(n_1029), .C(n_1122), .D(n_1125), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g1251 ( .A(n_1236), .B(n_1182), .Y(n_1251) );
NOR4xp25_ASAP7_75t_L g1252 ( .A(n_1245), .B(n_1237), .C(n_1235), .D(n_1242), .Y(n_1252) );
INVx2_ASAP7_75t_SL g1253 ( .A(n_1248), .Y(n_1253) );
NAND3xp33_ASAP7_75t_L g1254 ( .A(n_1250), .B(n_1135), .C(n_1123), .Y(n_1254) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1246), .Y(n_1255) );
NOR2x1p5_ASAP7_75t_L g1256 ( .A(n_1249), .B(n_1066), .Y(n_1256) );
AOI22xp5_ASAP7_75t_L g1257 ( .A1(n_1255), .A2(n_1251), .B1(n_1247), .B2(n_1029), .Y(n_1257) );
AOI22xp5_ASAP7_75t_L g1258 ( .A1(n_1252), .A2(n_1029), .B1(n_1125), .B2(n_1122), .Y(n_1258) );
OR2x2_ASAP7_75t_L g1259 ( .A(n_1253), .B(n_1126), .Y(n_1259) );
INVx3_ASAP7_75t_L g1260 ( .A(n_1256), .Y(n_1260) );
INVx2_ASAP7_75t_L g1261 ( .A(n_1259), .Y(n_1261) );
INVx2_ASAP7_75t_L g1262 ( .A(n_1260), .Y(n_1262) );
AND4x1_ASAP7_75t_L g1263 ( .A(n_1258), .B(n_1254), .C(n_1135), .D(n_1116), .Y(n_1263) );
HB1xp67_ASAP7_75t_L g1264 ( .A(n_1262), .Y(n_1264) );
INVx2_ASAP7_75t_L g1265 ( .A(n_1261), .Y(n_1265) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_1263), .B(n_1257), .Y(n_1266) );
AO21x2_ASAP7_75t_L g1267 ( .A1(n_1264), .A2(n_1029), .B(n_1094), .Y(n_1267) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1265), .Y(n_1268) );
OAI22xp5_ASAP7_75t_L g1269 ( .A1(n_1266), .A2(n_995), .B1(n_1047), .B2(n_1094), .Y(n_1269) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1268), .Y(n_1270) );
AO221x2_ASAP7_75t_L g1271 ( .A1(n_1270), .A2(n_1269), .B1(n_1267), .B2(n_1091), .C(n_1098), .Y(n_1271) );
AOI21xp5_ASAP7_75t_L g1272 ( .A1(n_1271), .A2(n_973), .B(n_977), .Y(n_1272) );
endmodule