module real_jpeg_13405_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_43;
wire n_8;
wire n_37;
wire n_21;
wire n_33;
wire n_38;
wire n_35;
wire n_29;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_48;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_0),
.B(n_20),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g9 ( 
.A(n_1),
.B(n_3),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_12),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_1),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_1),
.B(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_1),
.B(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_1),
.B(n_45),
.Y(n_49)
);

OR2x2_ASAP7_75t_SL g13 ( 
.A(n_2),
.B(n_14),
.Y(n_13)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_2),
.B(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_3),
.B(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_3),
.B(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_5),
.A2(n_17),
.B1(n_18),
.B2(n_23),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

AO21x1_ASAP7_75t_SL g27 ( 
.A1(n_5),
.A2(n_19),
.B(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g6 ( 
.A(n_7),
.Y(n_6)
);

AOI211xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_10),
.B(n_24),
.C(n_48),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_9),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_15),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_12),
.B(n_16),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_13),
.Y(n_12)
);

OR2x2_ASAP7_75t_SL g30 ( 
.A(n_14),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_14),
.B(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_18),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_21),
.Y(n_18)
);

OA21x2_ASAP7_75t_L g33 ( 
.A1(n_19),
.A2(n_23),
.B(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

NAND4xp25_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_37),
.C(n_42),
.D(n_46),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B1(n_32),
.B2(n_34),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_30),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_38),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_41),
.B(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);


endmodule