module fake_jpeg_18580_n_397 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_397);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_397;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_2),
.B(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_45),
.B(n_58),
.Y(n_115)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_25),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_51),
.Y(n_91)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_50),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_25),
.B(n_0),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_0),
.B(n_2),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_52),
.A2(n_59),
.B(n_26),
.C(n_28),
.Y(n_92)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_53),
.Y(n_138)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_22),
.B(n_14),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_55),
.B(n_64),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

OR2x2_ASAP7_75t_SL g59 ( 
.A(n_22),
.B(n_12),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_60),
.B(n_63),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_33),
.B(n_34),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_61),
.B(n_82),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_15),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_0),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_40),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_66),
.B(n_68),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_67),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_2),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_73),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_75),
.A2(n_87),
.B1(n_24),
.B2(n_42),
.Y(n_105)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_15),
.Y(n_80)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_19),
.B(n_23),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_83),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_137)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_15),
.Y(n_84)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_16),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_85),
.A2(n_86),
.B1(n_28),
.B2(n_26),
.Y(n_97)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_61),
.A2(n_52),
.B1(n_83),
.B2(n_75),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_90),
.A2(n_93),
.B1(n_96),
.B2(n_108),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_92),
.B(n_70),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_59),
.A2(n_38),
.B1(n_41),
.B2(n_23),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_48),
.A2(n_20),
.B1(n_41),
.B2(n_36),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_97),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_65),
.A2(n_24),
.B1(n_16),
.B2(n_32),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_98),
.A2(n_110),
.B1(n_113),
.B2(n_119),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_27),
.C(n_30),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_100),
.B(n_78),
.C(n_69),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_105),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_71),
.A2(n_79),
.B1(n_87),
.B2(n_77),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_49),
.A2(n_24),
.B1(n_32),
.B2(n_31),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_51),
.A2(n_36),
.B1(n_31),
.B2(n_20),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_55),
.A2(n_19),
.B(n_43),
.C(n_30),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_118),
.B(n_72),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_54),
.A2(n_27),
.B1(n_30),
.B2(n_43),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_58),
.A2(n_27),
.B1(n_43),
.B2(n_5),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_121),
.A2(n_50),
.B1(n_62),
.B2(n_44),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_76),
.A2(n_86),
.B1(n_53),
.B2(n_46),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_123),
.A2(n_131),
.B1(n_133),
.B2(n_9),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_85),
.A2(n_84),
.B1(n_3),
.B2(n_5),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_81),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_128),
.A2(n_99),
.B1(n_116),
.B2(n_136),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_73),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_73),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_139),
.A2(n_101),
.B1(n_124),
.B2(n_112),
.Y(n_189)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_141),
.Y(n_215)
);

INVx5_ASAP7_75t_SL g142 ( 
.A(n_94),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_142),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_143),
.B(n_151),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_57),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_144),
.B(n_168),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_134),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_146),
.B(n_148),
.Y(n_187)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_135),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_149),
.Y(n_205)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_152),
.A2(n_173),
.B1(n_175),
.B2(n_114),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_132),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_154),
.B(n_158),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_90),
.A2(n_56),
.B(n_78),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g219 ( 
.A(n_157),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_67),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_103),
.B(n_67),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_170),
.Y(n_186)
);

INVx11_ASAP7_75t_L g161 ( 
.A(n_94),
.Y(n_161)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_106),
.Y(n_163)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_163),
.Y(n_202)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_104),
.Y(n_164)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_164),
.Y(n_206)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

AOI21xp33_ASAP7_75t_L g166 ( 
.A1(n_91),
.A2(n_11),
.B(n_12),
.Y(n_166)
);

NOR3xp33_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_121),
.C(n_124),
.Y(n_184)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_167),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_92),
.B(n_47),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_169),
.B(n_175),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_134),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_91),
.B(n_74),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_174),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_120),
.B(n_11),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_176),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_98),
.A2(n_12),
.B1(n_110),
.B2(n_127),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_125),
.B(n_118),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_99),
.A2(n_127),
.B1(n_116),
.B2(n_136),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_126),
.B(n_115),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_177),
.A2(n_106),
.B1(n_138),
.B2(n_109),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_102),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_180),
.Y(n_209)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_108),
.Y(n_179)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_179),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_88),
.B(n_107),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_89),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_95),
.B(n_102),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_147),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_184),
.B(n_147),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_189),
.A2(n_200),
.B1(n_214),
.B2(n_153),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_179),
.A2(n_101),
.B1(n_112),
.B2(n_109),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_194),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_140),
.A2(n_114),
.B1(n_111),
.B2(n_122),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_196),
.A2(n_201),
.B1(n_212),
.B2(n_216),
.Y(n_233)
);

OAI22x1_ASAP7_75t_SL g199 ( 
.A1(n_145),
.A2(n_111),
.B1(n_122),
.B2(n_129),
.Y(n_199)
);

OA22x2_ASAP7_75t_L g239 ( 
.A1(n_199),
.A2(n_150),
.B1(n_161),
.B2(n_141),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_144),
.B(n_129),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_210),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_171),
.B(n_138),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_211),
.B(n_181),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_140),
.A2(n_145),
.B1(n_168),
.B2(n_143),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_182),
.A2(n_173),
.B1(n_155),
.B2(n_152),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_155),
.A2(n_174),
.B1(n_153),
.B2(n_159),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_170),
.B(n_151),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_169),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_220),
.A2(n_164),
.B1(n_142),
.B2(n_157),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_156),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_248),
.C(n_220),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_203),
.B(n_154),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_225),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_206),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_226),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_229),
.Y(n_255)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_218),
.Y(n_228)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_228),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_182),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_219),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_231),
.A2(n_235),
.B(n_239),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_204),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_237),
.Y(n_263)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_234),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_193),
.B(n_159),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_202),
.Y(n_236)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_236),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_146),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_195),
.B(n_148),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_238),
.B(n_248),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_240),
.A2(n_247),
.B1(n_253),
.B2(n_192),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_241),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_242),
.B(n_254),
.Y(n_268)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_202),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_243),
.Y(n_283)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_215),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_244),
.Y(n_256)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_245),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_197),
.B(n_178),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_246),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_214),
.A2(n_150),
.B1(n_142),
.B2(n_163),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_165),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_196),
.A2(n_220),
.B1(n_192),
.B2(n_216),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_249),
.A2(n_208),
.B1(n_191),
.B2(n_190),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_195),
.B(n_167),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_250),
.A2(n_185),
.B(n_213),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_251),
.Y(n_259)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_215),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_252),
.Y(n_277)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_221),
.Y(n_253)
);

MAJx2_ASAP7_75t_L g254 ( 
.A(n_193),
.B(n_181),
.C(n_186),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_257),
.B(n_273),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_258),
.A2(n_275),
.B1(n_239),
.B2(n_226),
.Y(n_295)
);

AO22x1_ASAP7_75t_L g260 ( 
.A1(n_229),
.A2(n_199),
.B1(n_210),
.B2(n_207),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_260),
.B(n_262),
.Y(n_308)
);

AO22x1_ASAP7_75t_L g262 ( 
.A1(n_237),
.A2(n_200),
.B1(n_205),
.B2(n_189),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_240),
.A2(n_205),
.B1(n_187),
.B2(n_209),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_265),
.A2(n_242),
.B1(n_224),
.B2(n_254),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_266),
.A2(n_271),
.B1(n_278),
.B2(n_252),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_222),
.A2(n_208),
.B(n_185),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_267),
.A2(n_279),
.B(n_272),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_233),
.A2(n_191),
.B1(n_190),
.B2(n_213),
.Y(n_271)
);

OAI22x1_ASAP7_75t_SL g275 ( 
.A1(n_233),
.A2(n_239),
.B1(n_247),
.B2(n_249),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_276),
.A2(n_235),
.B1(n_228),
.B2(n_234),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_227),
.A2(n_188),
.B1(n_221),
.B2(n_219),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_230),
.A2(n_188),
.B(n_219),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_276),
.Y(n_284)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_284),
.Y(n_309)
);

INVx8_ASAP7_75t_L g285 ( 
.A(n_275),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_286),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_264),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_281),
.Y(n_287)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_287),
.Y(n_312)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_281),
.Y(n_288)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_288),
.Y(n_317)
);

BUFx12f_ASAP7_75t_SL g289 ( 
.A(n_267),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_289),
.B(n_302),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_290),
.A2(n_292),
.B1(n_303),
.B2(n_304),
.Y(n_315)
);

OAI32xp33_ASAP7_75t_L g291 ( 
.A1(n_255),
.A2(n_232),
.A3(n_250),
.B1(n_273),
.B2(n_263),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_291),
.B(n_306),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_293),
.A2(n_294),
.B1(n_295),
.B2(n_297),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_258),
.A2(n_224),
.B1(n_225),
.B2(n_239),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_261),
.B(n_231),
.Y(n_296)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_296),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_255),
.A2(n_235),
.B1(n_238),
.B2(n_236),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_257),
.B(n_243),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_305),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_264),
.Y(n_300)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_300),
.Y(n_323)
);

A2O1A1O1Ixp25_ASAP7_75t_L g301 ( 
.A1(n_268),
.A2(n_244),
.B(n_245),
.C(n_253),
.D(n_263),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_301),
.B(n_278),
.Y(n_313)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_269),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_269),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_268),
.B(n_265),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_272),
.B(n_270),
.Y(n_306)
);

AO22x1_ASAP7_75t_SL g307 ( 
.A1(n_260),
.A2(n_262),
.B1(n_271),
.B2(n_266),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_307),
.A2(n_283),
.B1(n_277),
.B2(n_256),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_313),
.B(n_325),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_285),
.A2(n_260),
.B1(n_262),
.B2(n_259),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_314),
.B(n_326),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_279),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_316),
.B(n_318),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_305),
.B(n_282),
.Y(n_318)
);

FAx1_ASAP7_75t_SL g319 ( 
.A(n_297),
.B(n_282),
.CI(n_259),
.CON(n_319),
.SN(n_319)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_319),
.B(n_307),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_298),
.B(n_270),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_294),
.A2(n_280),
.B1(n_277),
.B2(n_283),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_327),
.A2(n_306),
.B1(n_308),
.B2(n_289),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_299),
.B(n_274),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_328),
.B(n_329),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_293),
.B(n_274),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_320),
.B(n_308),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_330),
.B(n_334),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_331),
.A2(n_343),
.B1(n_336),
.B2(n_345),
.Y(n_357)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_323),
.Y(n_332)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_332),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_319),
.B(n_302),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_322),
.A2(n_304),
.B(n_306),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_335),
.A2(n_342),
.B(n_339),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_292),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_337),
.Y(n_353)
);

NAND4xp25_ASAP7_75t_L g338 ( 
.A(n_314),
.B(n_301),
.C(n_290),
.D(n_291),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_338),
.B(n_339),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_311),
.B(n_307),
.Y(n_340)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_340),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_322),
.A2(n_309),
.B(n_313),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_316),
.A2(n_315),
.B1(n_312),
.B2(n_317),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_324),
.B(n_321),
.Y(n_345)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_345),
.Y(n_358)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_324),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_346),
.B(n_333),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_325),
.B(n_310),
.C(n_328),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_310),
.C(n_318),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_348),
.B(n_354),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_340),
.B(n_336),
.Y(n_350)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_350),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_342),
.A2(n_329),
.B1(n_335),
.B2(n_331),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_351),
.A2(n_358),
.B1(n_353),
.B2(n_360),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_347),
.B(n_341),
.C(n_333),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_355),
.B(n_341),
.C(n_344),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_357),
.B(n_360),
.Y(n_362)
);

INVx11_ASAP7_75t_L g361 ( 
.A(n_343),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_361),
.A2(n_356),
.B1(n_353),
.B2(n_350),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_364),
.B(n_372),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_359),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_365),
.B(n_371),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_349),
.B(n_344),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_366),
.A2(n_358),
.B(n_356),
.Y(n_374)
);

BUFx4f_ASAP7_75t_SL g367 ( 
.A(n_352),
.Y(n_367)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_367),
.Y(n_376)
);

BUFx4f_ASAP7_75t_SL g369 ( 
.A(n_352),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_369),
.B(n_370),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_349),
.A2(n_359),
.B(n_354),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_374),
.A2(n_378),
.B(n_369),
.Y(n_387)
);

INVx6_ASAP7_75t_L g375 ( 
.A(n_362),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_375),
.B(n_381),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_368),
.B(n_357),
.Y(n_377)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_377),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_366),
.A2(n_361),
.B(n_348),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_367),
.A2(n_361),
.B1(n_369),
.B2(n_363),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_373),
.B(n_363),
.Y(n_383)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_383),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_376),
.B(n_367),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_384),
.A2(n_386),
.B(n_385),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_379),
.B(n_364),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_387),
.A2(n_384),
.B(n_380),
.Y(n_391)
);

AOI31xp67_ASAP7_75t_SL g388 ( 
.A1(n_382),
.A2(n_381),
.A3(n_378),
.B(n_374),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_388),
.B(n_390),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_391),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_393),
.B(n_389),
.C(n_380),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_394),
.A2(n_395),
.B(n_355),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_392),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_396),
.B(n_375),
.Y(n_397)
);


endmodule