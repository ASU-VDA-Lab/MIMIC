module fake_jpeg_13371_n_298 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

BUFx10_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_0),
.B(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

CKINVDCx6p67_ASAP7_75t_R g94 ( 
.A(n_47),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_49),
.B(n_67),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_50),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_51),
.Y(n_130)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_52),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

HAxp5_ASAP7_75t_SL g56 ( 
.A(n_16),
.B(n_0),
.CON(n_56),
.SN(n_56)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_56),
.B(n_60),
.Y(n_126)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_26),
.B(n_9),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_68),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_26),
.B(n_9),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_28),
.B(n_9),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_64),
.B(n_79),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_27),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_73),
.Y(n_98)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_28),
.B(n_39),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_36),
.Y(n_91)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_76),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_78),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_35),
.B(n_8),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_81),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_83),
.Y(n_106)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_85),
.Y(n_108)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_31),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_56),
.A2(n_23),
.B1(n_27),
.B2(n_44),
.Y(n_88)
);

OAI22x1_ASAP7_75t_L g153 ( 
.A1(n_88),
.A2(n_89),
.B1(n_92),
.B2(n_123),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_47),
.A2(n_24),
.B1(n_44),
.B2(n_25),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_24),
.B1(n_20),
.B2(n_37),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_90),
.A2(n_128),
.B1(n_135),
.B2(n_94),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_91),
.B(n_119),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_53),
.A2(n_20),
.B1(n_25),
.B2(n_37),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_86),
.A2(n_31),
.B1(n_29),
.B2(n_17),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_109),
.A2(n_115),
.B1(n_122),
.B2(n_133),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_110),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_81),
.A2(n_48),
.B1(n_76),
.B2(n_66),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_49),
.B(n_29),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_118),
.B(n_120),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_60),
.B(n_36),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_64),
.B(n_39),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_79),
.A2(n_35),
.B1(n_65),
.B2(n_58),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_84),
.A2(n_41),
.B1(n_1),
.B2(n_4),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_50),
.B(n_3),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_124),
.B(n_128),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_67),
.A2(n_41),
.B1(n_4),
.B2(n_6),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_68),
.A2(n_41),
.B1(n_4),
.B2(n_6),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_129),
.A2(n_131),
.B1(n_113),
.B2(n_94),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_69),
.A2(n_41),
.B1(n_10),
.B2(n_11),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_49),
.A2(n_3),
.B1(n_12),
.B2(n_15),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_80),
.A2(n_3),
.B1(n_12),
.B2(n_81),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_136),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_145),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_138),
.B(n_142),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_126),
.A2(n_118),
.B(n_91),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_139),
.A2(n_172),
.B(n_173),
.Y(n_196)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

AO22x1_ASAP7_75t_SL g141 ( 
.A1(n_117),
.A2(n_126),
.B1(n_97),
.B2(n_134),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_168),
.Y(n_178)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_143),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_107),
.B(n_120),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_144),
.B(n_167),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_99),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_96),
.B(n_106),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_146),
.Y(n_193)
);

NOR2x1_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_171),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_102),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_154),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_130),
.Y(n_149)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_149),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_150),
.A2(n_151),
.B1(n_157),
.B2(n_161),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_124),
.A2(n_90),
.B1(n_104),
.B2(n_103),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_94),
.B(n_93),
.Y(n_154)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_94),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_159),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_93),
.B(n_105),
.Y(n_159)
);

INVx11_ASAP7_75t_L g160 ( 
.A(n_101),
.Y(n_160)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_108),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_163),
.Y(n_187)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_105),
.B(n_114),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_L g164 ( 
.A1(n_109),
.A2(n_130),
.B(n_97),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_166),
.Y(n_198)
);

AO22x1_ASAP7_75t_L g165 ( 
.A1(n_134),
.A2(n_127),
.B1(n_103),
.B2(n_112),
.Y(n_165)
);

O2A1O1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_165),
.A2(n_172),
.B(n_160),
.C(n_140),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_95),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_95),
.B(n_87),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_87),
.B(n_112),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_174),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_121),
.Y(n_170)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_121),
.Y(n_171)
);

NAND2xp33_ASAP7_75t_SL g172 ( 
.A(n_100),
.B(n_132),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_125),
.A2(n_100),
.B(n_132),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_125),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_155),
.A2(n_142),
.B1(n_151),
.B2(n_145),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_180),
.A2(n_191),
.B1(n_192),
.B2(n_194),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_185),
.Y(n_210)
);

OAI32xp33_ASAP7_75t_L g185 ( 
.A1(n_167),
.A2(n_144),
.A3(n_141),
.B1(n_139),
.B2(n_138),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_138),
.B(n_148),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_162),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_190),
.A2(n_178),
.B1(n_196),
.B2(n_192),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_155),
.A2(n_150),
.B1(n_141),
.B2(n_153),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_153),
.A2(n_173),
.B1(n_174),
.B2(n_170),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_158),
.A2(n_137),
.B1(n_165),
.B2(n_171),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_202),
.A2(n_166),
.B1(n_165),
.B2(n_156),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_188),
.B(n_136),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_205),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_216),
.Y(n_226)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_197),
.Y(n_209)
);

OAI21xp33_ASAP7_75t_SL g234 ( 
.A1(n_209),
.A2(n_175),
.B(n_189),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_211),
.A2(n_195),
.B1(n_184),
.B2(n_189),
.Y(n_230)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_201),
.Y(n_212)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_190),
.A2(n_143),
.B1(n_152),
.B2(n_149),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_213),
.A2(n_217),
.B1(n_206),
.B2(n_205),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_149),
.Y(n_214)
);

NAND3xp33_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_215),
.C(n_218),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_187),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_180),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_200),
.Y(n_218)
);

NOR3xp33_ASAP7_75t_SL g219 ( 
.A(n_178),
.B(n_185),
.C(n_181),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_219),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_194),
.A2(n_196),
.B1(n_202),
.B2(n_191),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_220),
.A2(n_208),
.B1(n_221),
.B2(n_216),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_181),
.Y(n_221)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_221),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_177),
.B(n_193),
.Y(n_222)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_222),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_223),
.Y(n_237)
);

A2O1A1O1Ixp25_ASAP7_75t_L g224 ( 
.A1(n_186),
.A2(n_197),
.B(n_201),
.C(n_203),
.D(n_199),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_224),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_199),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_195),
.C(n_184),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_225),
.A2(n_186),
.B(n_175),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_228),
.A2(n_213),
.B(n_223),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_230),
.A2(n_243),
.B1(n_235),
.B2(n_226),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_239),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_236),
.B(n_220),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_204),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_240),
.A2(n_208),
.B1(n_211),
.B2(n_224),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_222),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_219),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_210),
.C(n_217),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_245),
.C(n_256),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_247),
.A2(n_232),
.B1(n_240),
.B2(n_230),
.Y(n_261)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_207),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_251),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_250),
.A2(n_257),
.B(n_258),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_233),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_252),
.B(n_254),
.Y(n_259)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_227),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_253),
.A2(n_255),
.B1(n_237),
.B2(n_231),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_233),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_227),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_212),
.C(n_209),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_226),
.Y(n_257)
);

AO21x1_ASAP7_75t_L g258 ( 
.A1(n_238),
.A2(n_243),
.B(n_229),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_261),
.A2(n_263),
.B1(n_269),
.B2(n_258),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_247),
.A2(n_232),
.B1(n_237),
.B2(n_231),
.Y(n_263)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_264),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_241),
.C(n_244),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_262),
.Y(n_271)
);

NOR3xp33_ASAP7_75t_SL g267 ( 
.A(n_248),
.B(n_246),
.C(n_249),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_267),
.B(n_253),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_251),
.A2(n_254),
.B1(n_250),
.B2(n_246),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_266),
.A2(n_257),
.B1(n_256),
.B2(n_252),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_270),
.A2(n_273),
.B1(n_275),
.B2(n_268),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_271),
.A2(n_272),
.B(n_263),
.Y(n_282)
);

FAx1_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_258),
.CI(n_255),
.CON(n_272),
.SN(n_272)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_274),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_260),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_267),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_269),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_262),
.C(n_265),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_278),
.A2(n_276),
.B(n_277),
.Y(n_286)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_279),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_281),
.A2(n_272),
.B1(n_277),
.B2(n_283),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_283),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_261),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_280),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_279),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_278),
.Y(n_291)
);

INVxp33_ASAP7_75t_L g290 ( 
.A(n_287),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_291),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_288),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_293),
.B(n_290),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_294),
.Y(n_296)
);

AND2x4_ASAP7_75t_L g295 ( 
.A(n_292),
.B(n_285),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_295),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_293),
.Y(n_298)
);


endmodule