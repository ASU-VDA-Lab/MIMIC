module fake_jpeg_23217_n_93 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_93);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_93;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

BUFx10_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx2_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_8),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

OAI21xp33_ASAP7_75t_L g21 ( 
.A1(n_13),
.A2(n_0),
.B(n_1),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_21),
.A2(n_23),
.B1(n_27),
.B2(n_18),
.Y(n_33)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_25),
.Y(n_39)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_28),
.Y(n_30)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_20),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_L g32 ( 
.A1(n_22),
.A2(n_18),
.B1(n_17),
.B2(n_16),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_34),
.B1(n_36),
.B2(n_17),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_25),
.B1(n_28),
.B2(n_11),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_27),
.A2(n_18),
.B1(n_13),
.B2(n_19),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_26),
.A2(n_19),
.B1(n_10),
.B2(n_14),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

O2A1O1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_50),
.B(n_48),
.C(n_41),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_33),
.B(n_30),
.C(n_20),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_45),
.B(n_47),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_37),
.A2(n_25),
.B(n_28),
.C(n_24),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_50),
.B1(n_29),
.B2(n_20),
.Y(n_55)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_30),
.B(n_10),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_25),
.B1(n_28),
.B2(n_12),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_48),
.A2(n_11),
.B1(n_2),
.B2(n_3),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_31),
.B(n_14),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_20),
.Y(n_52)
);

FAx1_ASAP7_75t_SL g61 ( 
.A(n_52),
.B(n_0),
.CI(n_2),
.CON(n_61),
.SN(n_61)
);

AND2x6_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_7),
.Y(n_53)
);

XNOR2x1_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_56),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_55),
.B1(n_60),
.B2(n_56),
.Y(n_63)
);

OR2x4_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_20),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_11),
.B(n_2),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_61),
.C(n_44),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_SL g70 ( 
.A(n_62),
.B(n_61),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_64),
.Y(n_72)
);

NOR3xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_51),
.C(n_43),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_68),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_6),
.C(n_9),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_68),
.Y(n_79)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_71),
.B(n_76),
.Y(n_80)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_72),
.A2(n_66),
.B(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_78),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_SL g78 ( 
.A1(n_75),
.A2(n_65),
.B(n_54),
.C(n_61),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_81),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_58),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_58),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_84),
.A2(n_71),
.B(n_74),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_73),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_83),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_86),
.B(n_9),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_78),
.C(n_75),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_89),
.B(n_90),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_87),
.A2(n_0),
.B(n_3),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_91),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_88),
.Y(n_93)
);


endmodule