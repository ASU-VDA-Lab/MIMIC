module fake_jpeg_16693_n_350 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_350);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_350;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_22),
.Y(n_65)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_48),
.Y(n_62)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_60),
.Y(n_93)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_22),
.B1(n_29),
.B2(n_23),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_63),
.A2(n_26),
.B1(n_34),
.B2(n_31),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_65),
.Y(n_82)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_76),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_37),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_71),
.B(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_37),
.Y(n_73)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_35),
.Y(n_76)
);

CKINVDCx5p33_ASAP7_75t_R g78 ( 
.A(n_39),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_80),
.Y(n_110)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_35),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_85),
.Y(n_116)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_68),
.A2(n_29),
.B1(n_44),
.B2(n_48),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_87),
.A2(n_57),
.B1(n_39),
.B2(n_49),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_63),
.A2(n_29),
.B1(n_48),
.B2(n_49),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_88),
.A2(n_107),
.B1(n_111),
.B2(n_112),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_23),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_94),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_59),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g96 ( 
.A1(n_70),
.A2(n_24),
.B(n_28),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_96),
.A2(n_30),
.B(n_33),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_33),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_102),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_45),
.Y(n_124)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_66),
.Y(n_100)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_33),
.Y(n_102)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_55),
.A2(n_24),
.B1(n_18),
.B2(n_31),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_70),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_109),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_55),
.A2(n_34),
.B1(n_26),
.B2(n_28),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_74),
.A2(n_52),
.B1(n_51),
.B2(n_47),
.Y(n_111)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_117),
.A2(n_129),
.B1(n_134),
.B2(n_139),
.Y(n_152)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_94),
.A2(n_42),
.B(n_18),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_136),
.Y(n_154)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_124),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_89),
.B(n_45),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_137),
.Y(n_151)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_30),
.B(n_32),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_74),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_133),
.Y(n_162)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_103),
.B(n_20),
.Y(n_135)
);

BUFx24_ASAP7_75t_SL g147 ( 
.A(n_135),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_82),
.B(n_42),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_92),
.B(n_45),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_93),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_140),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_84),
.B(n_77),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_88),
.A2(n_57),
.B1(n_47),
.B2(n_51),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_141),
.A2(n_101),
.B1(n_86),
.B2(n_105),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_85),
.B(n_32),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_142),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_97),
.B(n_102),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_42),
.Y(n_167)
);

FAx1_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_87),
.CI(n_112),
.CON(n_144),
.SN(n_144)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_144),
.B(n_141),
.Y(n_171)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_145),
.A2(n_115),
.B1(n_117),
.B2(n_131),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_139),
.B1(n_134),
.B2(n_115),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_129),
.A2(n_101),
.B1(n_91),
.B2(n_90),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_155),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_113),
.A2(n_101),
.B1(n_106),
.B2(n_90),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_158),
.A2(n_159),
.B1(n_163),
.B2(n_119),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_120),
.A2(n_86),
.B1(n_91),
.B2(n_95),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_126),
.A2(n_95),
.B1(n_98),
.B2(n_100),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_127),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_168),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_166),
.B(n_132),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_120),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_127),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_169),
.A2(n_145),
.B1(n_164),
.B2(n_165),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_SL g194 ( 
.A(n_170),
.B(n_172),
.C(n_176),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_171),
.A2(n_178),
.B(n_149),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_149),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_173),
.B(n_184),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_136),
.C(n_143),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_190),
.C(n_157),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_156),
.Y(n_175)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_175),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_144),
.A2(n_126),
.B1(n_140),
.B2(n_137),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_177),
.A2(n_192),
.B1(n_52),
.B2(n_47),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_130),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_181),
.A2(n_146),
.B1(n_158),
.B2(n_162),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_128),
.Y(n_182)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_156),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_150),
.Y(n_185)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_187),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_128),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_189),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_144),
.B(n_163),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_138),
.C(n_122),
.Y(n_190)
);

OA21x2_ASAP7_75t_L g191 ( 
.A1(n_144),
.A2(n_128),
.B(n_116),
.Y(n_191)
);

OA22x2_ASAP7_75t_L g220 ( 
.A1(n_191),
.A2(n_52),
.B1(n_46),
.B2(n_67),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_152),
.A2(n_125),
.B1(n_121),
.B2(n_123),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_195),
.A2(n_210),
.B1(n_213),
.B2(n_215),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_189),
.A2(n_155),
.B(n_162),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_196),
.A2(n_201),
.B(n_220),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_218),
.C(n_172),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_159),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_164),
.Y(n_203)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_179),
.Y(n_204)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

AO22x1_ASAP7_75t_L g206 ( 
.A1(n_191),
.A2(n_145),
.B1(n_161),
.B2(n_160),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_211),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_208),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_186),
.Y(n_209)
);

INVxp33_ASAP7_75t_SL g234 ( 
.A(n_209),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_181),
.A2(n_168),
.B1(n_148),
.B2(n_153),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_173),
.Y(n_212)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_193),
.A2(n_148),
.B1(n_125),
.B2(n_121),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_214),
.B(n_177),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_169),
.A2(n_147),
.B1(n_108),
.B2(n_51),
.Y(n_215)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_216),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_174),
.B(n_42),
.C(n_77),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_191),
.A2(n_67),
.B1(n_61),
.B2(n_127),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_219),
.A2(n_182),
.B1(n_179),
.B2(n_180),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_227),
.C(n_218),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_224),
.B(n_238),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_190),
.Y(n_227)
);

NAND3xp33_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_188),
.C(n_193),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_236),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_178),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_242),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_195),
.A2(n_191),
.B1(n_183),
.B2(n_185),
.Y(n_231)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_233),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_210),
.A2(n_192),
.B1(n_180),
.B2(n_170),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_235),
.A2(n_201),
.B1(n_217),
.B2(n_205),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_197),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_202),
.A2(n_178),
.B1(n_187),
.B2(n_32),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_237),
.A2(n_240),
.B1(n_244),
.B2(n_25),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_196),
.A2(n_12),
.B(n_17),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_243),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_201),
.A2(n_194),
.B1(n_211),
.B2(n_212),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_202),
.B(n_33),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_200),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_206),
.A2(n_0),
.B(n_1),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_245),
.A2(n_241),
.B(n_244),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_248),
.C(n_254),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_205),
.C(n_217),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_226),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_255),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_252),
.A2(n_256),
.B1(n_258),
.B2(n_221),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_219),
.C(n_216),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_229),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_239),
.A2(n_194),
.B1(n_206),
.B2(n_220),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_241),
.A2(n_220),
.B1(n_212),
.B2(n_207),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_198),
.C(n_220),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_266),
.C(n_25),
.Y(n_283)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_234),
.Y(n_260)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_260),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_262),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_223),
.Y(n_263)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

FAx1_ASAP7_75t_SL g264 ( 
.A(n_237),
.B(n_33),
.CI(n_25),
.CON(n_264),
.SN(n_264)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_267),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_265),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_224),
.B(n_25),
.C(n_20),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_240),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_267),
.A2(n_225),
.B1(n_232),
.B2(n_245),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_270),
.A2(n_272),
.B1(n_280),
.B2(n_281),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_246),
.A2(n_221),
.B1(n_238),
.B2(n_242),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_274),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_10),
.Y(n_277)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_277),
.Y(n_297)
);

NOR2xp67_ASAP7_75t_SL g278 ( 
.A(n_248),
.B(n_10),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_278),
.A2(n_283),
.B(n_9),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_25),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_285),
.C(n_266),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_261),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_256),
.A2(n_251),
.B1(n_258),
.B2(n_252),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_249),
.B(n_21),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_284),
.B(n_249),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_21),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_253),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_265),
.Y(n_290)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_287),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_254),
.C(n_257),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_291),
.C(n_299),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_284),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_298),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_257),
.C(n_264),
.Y(n_291)
);

XOR2x2_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_264),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_293),
.A2(n_294),
.B(n_296),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_275),
.A2(n_9),
.B(n_15),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_271),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_9),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_276),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_300),
.A2(n_286),
.B(n_269),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_30),
.C(n_4),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_30),
.C(n_4),
.Y(n_313)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_280),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_3),
.Y(n_312)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_303),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_282),
.Y(n_306)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_306),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_297),
.B(n_281),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_309),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_270),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_311),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_283),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_312),
.B(n_4),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_301),
.C(n_287),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_293),
.A2(n_12),
.B(n_5),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_315),
.A2(n_300),
.B(n_5),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_12),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_14),
.Y(n_323)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_319),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_321),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_322),
.B(n_4),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_323),
.B(n_326),
.Y(n_331)
);

NOR2xp67_ASAP7_75t_L g325 ( 
.A(n_305),
.B(n_289),
.Y(n_325)
);

OAI21x1_ASAP7_75t_SL g333 ( 
.A1(n_325),
.A2(n_315),
.B(n_311),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_308),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_314),
.A2(n_291),
.B1(n_6),
.B2(n_11),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_327),
.B(n_313),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_330),
.B(n_332),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_304),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_335),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_317),
.A2(n_304),
.B(n_310),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_334),
.B(n_318),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_324),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_336),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_338),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_319),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_340),
.A2(n_329),
.B(n_13),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_335),
.Y(n_342)
);

OAI21x1_ASAP7_75t_L g344 ( 
.A1(n_342),
.A2(n_328),
.B(n_320),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_344),
.A2(n_345),
.B(n_337),
.Y(n_346)
);

OAI211xp5_ASAP7_75t_L g347 ( 
.A1(n_346),
.A2(n_343),
.B(n_341),
.C(n_339),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_347),
.A2(n_11),
.B(n_13),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_14),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_349),
.B(n_30),
.Y(n_350)
);


endmodule