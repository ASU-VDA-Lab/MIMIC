module fake_jpeg_5442_n_51 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_51);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_51;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx10_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_17),
.Y(n_22)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_18),
.A2(n_13),
.B1(n_10),
.B2(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_24),
.B(n_26),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_16),
.Y(n_25)
);

OAI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_25),
.A2(n_27),
.B1(n_14),
.B2(n_22),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_15),
.B1(n_19),
.B2(n_17),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_30),
.B(n_32),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_25),
.A2(n_15),
.B1(n_19),
.B2(n_14),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_21),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_21),
.B1(n_9),
.B2(n_11),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_35),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_31),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_33),
.B(n_10),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_37),
.B(n_38),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_29),
.C(n_18),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

AO21x1_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_43),
.B(n_12),
.Y(n_45)
);

AO221x1_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_12),
.B1(n_8),
.B2(n_3),
.C(n_1),
.Y(n_43)
);

OAI322xp33_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_40),
.A3(n_12),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_3),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_4),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_41),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_47),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_6),
.C(n_2),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_50),
.B(n_2),
.Y(n_51)
);


endmodule