module fake_jpeg_1730_n_148 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_148);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_59),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_58),
.Y(n_66)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_60),
.A2(n_43),
.B1(n_47),
.B2(n_45),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_50),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_52),
.B(n_53),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_69),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_38),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_70),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_56),
.A2(n_51),
.B1(n_48),
.B2(n_45),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_51),
.B1(n_50),
.B2(n_49),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_60),
.B1(n_54),
.B2(n_61),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_57),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_75),
.B(n_80),
.Y(n_98)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_81),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_40),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_40),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_84),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_61),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_0),
.Y(n_102)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_17),
.B1(n_32),
.B2(n_31),
.Y(n_95)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_26),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_55),
.B1(n_61),
.B2(n_42),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_99),
.B1(n_85),
.B2(n_77),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_39),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_91),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_77),
.Y(n_91)
);

INVxp67_ASAP7_75t_SL g104 ( 
.A(n_95),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_16),
.B1(n_30),
.B2(n_29),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_102),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_73),
.B(n_87),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_103),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_37),
.B1(n_28),
.B2(n_27),
.Y(n_99)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_0),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_12),
.B1(n_104),
.B2(n_111),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_93),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_109),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_89),
.C(n_90),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_110),
.Y(n_124)
);

AND2x6_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_25),
.Y(n_108)
);

AND2x6_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_120),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_1),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_24),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_92),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_114),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_2),
.B(n_3),
.Y(n_116)
);

NOR3xp33_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_121),
.C(n_7),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_4),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_5),
.Y(n_118)
);

AND2x6_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_22),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_90),
.A2(n_5),
.B(n_6),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_125),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_15),
.C(n_18),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_127),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_20),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_21),
.C(n_10),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_132),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_119),
.Y(n_135)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_135),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_124),
.C(n_115),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_138),
.C(n_126),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_115),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_140),
.B(n_141),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_139),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_134),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_143),
.A2(n_133),
.B(n_104),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_125),
.B(n_128),
.Y(n_145)
);

AOI21x1_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_108),
.B(n_120),
.Y(n_146)
);

BUFx24_ASAP7_75t_SL g147 ( 
.A(n_146),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_130),
.Y(n_148)
);


endmodule