module fake_jpeg_22081_n_187 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_187);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_15),
.B(n_17),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_32),
.B(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_0),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_26),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_42),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_3),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_31),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_4),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_4),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_4),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_45),
.A2(n_29),
.B1(n_28),
.B2(n_19),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_29),
.B1(n_28),
.B2(n_27),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_47),
.A2(n_70),
.B1(n_8),
.B2(n_9),
.Y(n_89)
);

OR2x2_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_27),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_49),
.A2(n_64),
.B(n_11),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_51),
.Y(n_88)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_69),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_53),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_91)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_58),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_29),
.B1(n_19),
.B2(n_31),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_67),
.B1(n_20),
.B2(n_18),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_63),
.Y(n_94)
);

MAJx2_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_27),
.C(n_22),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_10),
.Y(n_93)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_27),
.B(n_30),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_39),
.A2(n_25),
.B1(n_24),
.B2(n_23),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_71),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_22),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_37),
.A2(n_25),
.B1(n_24),
.B2(n_23),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_14),
.C(n_13),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_73),
.B(n_5),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_21),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_21),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_20),
.Y(n_78)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_82),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_81),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_93),
.Y(n_104)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_5),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_75),
.B(n_7),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_85),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_7),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_86),
.Y(n_111)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_8),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_60),
.B1(n_13),
.B2(n_12),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_91),
.A2(n_52),
.B1(n_47),
.B2(n_65),
.Y(n_103)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_49),
.Y(n_95)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_10),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_54),
.Y(n_118)
);

NAND2xp33_ASAP7_75t_SL g97 ( 
.A(n_62),
.B(n_69),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_97),
.A2(n_99),
.B(n_72),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_59),
.B(n_12),
.Y(n_101)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_93),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_56),
.C(n_51),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_79),
.C(n_84),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_113),
.B1(n_115),
.B2(n_96),
.Y(n_134)
);

CKINVDCx10_ASAP7_75t_R g112 ( 
.A(n_92),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_114),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_77),
.A2(n_87),
.B1(n_97),
.B2(n_91),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_94),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_72),
.B1(n_63),
.B2(n_55),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_86),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_118),
.B(n_76),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_54),
.B(n_46),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_46),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_123),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_48),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_112),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_124),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_119),
.A2(n_98),
.B1(n_100),
.B2(n_88),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_120),
.B1(n_103),
.B2(n_113),
.Y(n_144)
);

AOI221xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_134),
.B1(n_104),
.B2(n_105),
.C(n_115),
.Y(n_155)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_127),
.B(n_128),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_114),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_81),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_107),
.B(n_109),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_106),
.C(n_105),
.Y(n_156)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_116),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_110),
.Y(n_137)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_78),
.Y(n_138)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_90),
.Y(n_139)
);

OAI322xp33_ASAP7_75t_L g153 ( 
.A1(n_139),
.A2(n_140),
.A3(n_141),
.B1(n_107),
.B2(n_104),
.C1(n_120),
.C2(n_108),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_121),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_76),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_142),
.B(n_117),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_153),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_149),
.B(n_141),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_155),
.Y(n_166)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_154),
.A2(n_132),
.B(n_140),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_133),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_129),
.B1(n_134),
.B2(n_132),
.Y(n_158)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_162),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_163),
.Y(n_170)
);

AOI322xp5_ASAP7_75t_SL g162 ( 
.A1(n_150),
.A2(n_126),
.A3(n_128),
.B1(n_142),
.B2(n_144),
.C1(n_136),
.C2(n_156),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_165),
.C(n_152),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_169),
.C(n_172),
.Y(n_178)
);

MAJx2_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_126),
.C(n_154),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_139),
.C(n_138),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_127),
.C(n_135),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_160),
.Y(n_175)
);

AOI322xp5_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_161),
.A3(n_131),
.B1(n_165),
.B2(n_159),
.C1(n_147),
.C2(n_148),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_175),
.C(n_176),
.Y(n_181)
);

AOI322xp5_ASAP7_75t_L g176 ( 
.A1(n_171),
.A2(n_161),
.A3(n_131),
.B1(n_148),
.B2(n_157),
.C1(n_146),
.C2(n_151),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_146),
.Y(n_177)
);

NAND3xp33_ASAP7_75t_SL g180 ( 
.A(n_177),
.B(n_137),
.C(n_102),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_170),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_178),
.B(n_102),
.Y(n_182)
);

FAx1_ASAP7_75t_SL g183 ( 
.A(n_180),
.B(n_169),
.CI(n_122),
.CON(n_183),
.SN(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_48),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_183),
.A2(n_181),
.B(n_85),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_184),
.B(n_80),
.C(n_183),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_185),
.B(n_186),
.Y(n_187)
);


endmodule