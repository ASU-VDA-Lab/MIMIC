module fake_jpeg_8328_n_96 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_96);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_96;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_62;
wire n_43;
wire n_82;

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_40),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_34),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_8),
.B(n_33),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_3),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_0),
.Y(n_60)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

BUFx24_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_5),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_SL g76 ( 
.A(n_68),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

OR2x2_ASAP7_75t_SL g75 ( 
.A(n_69),
.B(n_70),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_6),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_58),
.B1(n_59),
.B2(n_55),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_77),
.A2(n_45),
.B1(n_50),
.B2(n_10),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_57),
.B1(n_51),
.B2(n_49),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_80),
.A2(n_81),
.B1(n_83),
.B2(n_76),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_7),
.C(n_9),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_71),
.B(n_11),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_12),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_13),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_88),
.A2(n_85),
.B1(n_75),
.B2(n_73),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_72),
.B1(n_19),
.B2(n_21),
.Y(n_90)
);

NAND4xp25_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_16),
.C(n_22),
.D(n_24),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_29),
.B(n_30),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_35),
.C(n_36),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_37),
.B(n_38),
.Y(n_95)
);

FAx1_ASAP7_75t_SL g96 ( 
.A(n_95),
.B(n_39),
.CI(n_74),
.CON(n_96),
.SN(n_96)
);


endmodule