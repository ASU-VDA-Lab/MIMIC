module fake_netlist_5_845_n_989 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_225, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_223, n_188, n_190, n_8, n_201, n_158, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_222, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_989);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_222;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_989;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_785;
wire n_316;
wire n_855;
wire n_389;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_916;
wire n_452;
wire n_885;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_841;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_526;
wire n_915;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_859;
wire n_864;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_932;
wire n_417;
wire n_946;
wire n_612;
wire n_385;
wire n_516;
wire n_498;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_509;
wire n_568;
wire n_936;
wire n_373;
wire n_947;
wire n_757;
wire n_820;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_394;
wire n_250;
wire n_579;
wire n_938;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_325;
wire n_449;
wire n_862;
wire n_900;
wire n_856;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_271;
wire n_934;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_654;
wire n_370;
wire n_976;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_961;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_255;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_680;
wire n_974;
wire n_395;
wire n_432;
wire n_553;
wire n_839;
wire n_901;
wire n_727;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_903;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_228;
wire n_283;
wire n_383;
wire n_781;
wire n_834;
wire n_711;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_963;
wire n_954;
wire n_627;
wire n_767;
wire n_440;
wire n_793;
wire n_478;
wire n_726;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_970;
wire n_911;
wire n_557;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_707;
wire n_710;
wire n_795;
wire n_695;
wire n_832;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_561;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_233;
wire n_404;
wire n_686;
wire n_366;
wire n_572;
wire n_754;
wire n_712;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_808;
wire n_409;
wire n_797;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_536;
wire n_531;
wire n_935;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_960;
wire n_759;
wire n_438;
wire n_806;
wire n_713;
wire n_904;
wire n_985;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_626;
wire n_925;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_67),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_161),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_207),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_109),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_33),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_74),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_136),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_48),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_210),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_127),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_56),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_21),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_205),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_142),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_175),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_214),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_93),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_100),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_94),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_213),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_209),
.Y(n_246)
);

BUFx5_ASAP7_75t_L g247 ( 
.A(n_170),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_39),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_112),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_35),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_221),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_7),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_96),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_8),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_186),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_115),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_196),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_200),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_204),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_179),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_172),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_208),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_225),
.Y(n_263)
);

BUFx2_ASAP7_75t_SL g264 ( 
.A(n_8),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_168),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_206),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_197),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_11),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_31),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_211),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_153),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_192),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_176),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_185),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_199),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_166),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_159),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_145),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_25),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_101),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_28),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_140),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_212),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_178),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_23),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_193),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_188),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_97),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_82),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_259),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_268),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_269),
.Y(n_292)
);

NOR2xp67_ASAP7_75t_L g293 ( 
.A(n_229),
.B(n_0),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_247),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_281),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_226),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_273),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_227),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_228),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_230),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_287),
.Y(n_302)
);

INVxp67_ASAP7_75t_SL g303 ( 
.A(n_231),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_272),
.B(n_276),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_234),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_232),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_235),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_285),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_281),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_233),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_239),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_236),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_238),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_247),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_240),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_237),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_244),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_L g318 ( 
.A(n_229),
.B(n_0),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_252),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_241),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_254),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_246),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_250),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_264),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_255),
.Y(n_325)
);

BUFx6f_ASAP7_75t_SL g326 ( 
.A(n_274),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_256),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_257),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_262),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_267),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_278),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_279),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_316),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_294),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_299),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_324),
.B(n_274),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_291),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_292),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_297),
.B(n_275),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_306),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_300),
.B(n_275),
.Y(n_341)
);

NOR2x1_ASAP7_75t_L g342 ( 
.A(n_305),
.B(n_280),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_310),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_295),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_312),
.Y(n_345)
);

INVxp33_ASAP7_75t_SL g346 ( 
.A(n_301),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_295),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_317),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_308),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_314),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_298),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_322),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_314),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_323),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_325),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_327),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_328),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_329),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_304),
.B(n_260),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_330),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_311),
.B(n_289),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_331),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_290),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_303),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_313),
.Y(n_365)
);

AND2x4_ASAP7_75t_L g366 ( 
.A(n_293),
.B(n_289),
.Y(n_366)
);

NOR2x1_ASAP7_75t_L g367 ( 
.A(n_307),
.B(n_282),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_326),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_326),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_302),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_318),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_319),
.Y(n_372)
);

BUFx8_ASAP7_75t_L g373 ( 
.A(n_296),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_320),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_315),
.Y(n_375)
);

AND2x4_ASAP7_75t_L g376 ( 
.A(n_316),
.B(n_283),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_321),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_332),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_321),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_332),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_296),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_359),
.B(n_242),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_359),
.B(n_243),
.Y(n_383)
);

INVx5_ASAP7_75t_L g384 ( 
.A(n_337),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_349),
.B(n_245),
.Y(n_385)
);

BUFx10_ASAP7_75t_L g386 ( 
.A(n_376),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_349),
.Y(n_387)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_353),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_336),
.B(n_248),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_344),
.B(n_347),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_372),
.B(n_249),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_353),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_335),
.Y(n_393)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_353),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_340),
.Y(n_395)
);

NAND2x1p5_ASAP7_75t_L g396 ( 
.A(n_374),
.B(n_284),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_371),
.Y(n_397)
);

INVx4_ASAP7_75t_L g398 ( 
.A(n_353),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_343),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_344),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_347),
.B(n_247),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_345),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_348),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_350),
.B(n_247),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_334),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_339),
.B(n_251),
.Y(n_406)
);

OR2x2_ASAP7_75t_SL g407 ( 
.A(n_378),
.B(n_288),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_346),
.Y(n_408)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_356),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_352),
.Y(n_410)
);

NAND2xp33_ASAP7_75t_L g411 ( 
.A(n_341),
.B(n_274),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_362),
.Y(n_412)
);

BUFx10_ASAP7_75t_L g413 ( 
.A(n_376),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_378),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_346),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_350),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_356),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_356),
.Y(n_418)
);

NAND2xp33_ASAP7_75t_L g419 ( 
.A(n_361),
.B(n_274),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_356),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_334),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_357),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_357),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_337),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_351),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_364),
.B(n_365),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_357),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_L g428 ( 
.A1(n_366),
.A2(n_247),
.B1(n_258),
.B2(n_253),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_366),
.B(n_247),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_351),
.B(n_261),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_342),
.B(n_263),
.Y(n_431)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_357),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_358),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_358),
.Y(n_434)
);

INVx5_ASAP7_75t_L g435 ( 
.A(n_337),
.Y(n_435)
);

INVx2_ASAP7_75t_SL g436 ( 
.A(n_336),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_358),
.Y(n_437)
);

INVx5_ASAP7_75t_L g438 ( 
.A(n_337),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_358),
.Y(n_439)
);

BUFx6f_ASAP7_75t_SL g440 ( 
.A(n_376),
.Y(n_440)
);

AND2x2_ASAP7_75t_SL g441 ( 
.A(n_333),
.B(n_309),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g442 ( 
.A(n_380),
.B(n_265),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_360),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_360),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_360),
.B(n_266),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_360),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_338),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_338),
.Y(n_448)
);

NAND2x1p5_ASAP7_75t_L g449 ( 
.A(n_421),
.B(n_367),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_400),
.Y(n_450)
);

OAI21xp33_ASAP7_75t_L g451 ( 
.A1(n_436),
.A2(n_369),
.B(n_368),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_390),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_418),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_390),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_416),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_406),
.B(n_366),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_393),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_395),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_408),
.Y(n_459)
);

INVxp67_ASAP7_75t_SL g460 ( 
.A(n_392),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_399),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_431),
.A2(n_375),
.B1(n_380),
.B2(n_271),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_402),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_403),
.Y(n_464)
);

NAND2x1p5_ASAP7_75t_L g465 ( 
.A(n_425),
.B(n_363),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_410),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_406),
.B(n_354),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_412),
.Y(n_468)
);

AO22x2_ASAP7_75t_L g469 ( 
.A1(n_414),
.A2(n_379),
.B1(n_377),
.B2(n_370),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_387),
.Y(n_470)
);

AO22x2_ASAP7_75t_L g471 ( 
.A1(n_414),
.A2(n_381),
.B1(n_309),
.B2(n_3),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_429),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g473 ( 
.A(n_385),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_426),
.B(n_354),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_428),
.A2(n_277),
.B1(n_286),
.B2(n_270),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_429),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_392),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_401),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_392),
.Y(n_479)
);

AO22x2_ASAP7_75t_L g480 ( 
.A1(n_431),
.A2(n_381),
.B1(n_3),
.B2(n_1),
.Y(n_480)
);

NAND2xp33_ASAP7_75t_L g481 ( 
.A(n_396),
.B(n_338),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_382),
.B(n_338),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_401),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_383),
.B(n_355),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_426),
.B(n_355),
.Y(n_485)
);

AO22x2_ASAP7_75t_L g486 ( 
.A1(n_442),
.A2(n_4),
.B1(n_1),
.B2(n_2),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_404),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_415),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_404),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_396),
.A2(n_373),
.B1(n_5),
.B2(n_2),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_405),
.Y(n_491)
);

CKINVDCx14_ASAP7_75t_R g492 ( 
.A(n_386),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_445),
.B(n_32),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_424),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_441),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_440),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_405),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_424),
.Y(n_498)
);

AO22x2_ASAP7_75t_L g499 ( 
.A1(n_389),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_397),
.B(n_391),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_397),
.A2(n_373),
.B1(n_36),
.B2(n_37),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_418),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_445),
.B(n_34),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_427),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_437),
.Y(n_505)
);

OA22x2_ASAP7_75t_L g506 ( 
.A1(n_407),
.A2(n_9),
.B1(n_6),
.B2(n_7),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_443),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_448),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_430),
.B(n_9),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_417),
.B(n_38),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_422),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_418),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_433),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_386),
.B(n_10),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_440),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_434),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_420),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_428),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_439),
.B(n_40),
.Y(n_519)
);

NAND2x1p5_ASAP7_75t_L g520 ( 
.A(n_409),
.B(n_41),
.Y(n_520)
);

AO22x2_ASAP7_75t_L g521 ( 
.A1(n_413),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_521)
);

NAND2xp33_ASAP7_75t_SL g522 ( 
.A(n_514),
.B(n_420),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_473),
.B(n_413),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_500),
.B(n_420),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_456),
.B(n_423),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_509),
.B(n_423),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_467),
.B(n_423),
.Y(n_527)
);

NAND2xp33_ASAP7_75t_SL g528 ( 
.A(n_518),
.B(n_444),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_474),
.B(n_485),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_491),
.B(n_444),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_452),
.B(n_446),
.Y(n_531)
);

NAND2xp33_ASAP7_75t_SL g532 ( 
.A(n_488),
.B(n_444),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_497),
.B(n_409),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_484),
.B(n_432),
.Y(n_534)
);

NAND2xp33_ASAP7_75t_SL g535 ( 
.A(n_459),
.B(n_447),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_470),
.B(n_432),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_452),
.B(n_388),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_457),
.B(n_384),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_458),
.B(n_384),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_461),
.B(n_384),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_449),
.B(n_465),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_463),
.B(n_438),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_464),
.B(n_388),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_466),
.B(n_468),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_472),
.B(n_435),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_454),
.B(n_394),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_476),
.B(n_435),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_454),
.B(n_394),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_462),
.B(n_438),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_482),
.B(n_438),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_478),
.B(n_435),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_483),
.B(n_398),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_475),
.B(n_398),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_487),
.B(n_411),
.Y(n_554)
);

NAND2xp33_ASAP7_75t_SL g555 ( 
.A(n_495),
.B(n_419),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_501),
.B(n_42),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_487),
.B(n_43),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_489),
.B(n_44),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_489),
.B(n_451),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_493),
.B(n_45),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_503),
.B(n_46),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_450),
.B(n_47),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_455),
.B(n_49),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_455),
.B(n_50),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_SL g565 ( 
.A(n_496),
.B(n_13),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_511),
.B(n_513),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_453),
.B(n_51),
.Y(n_567)
);

NAND2xp33_ASAP7_75t_SL g568 ( 
.A(n_512),
.B(n_14),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_453),
.B(n_52),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_502),
.B(n_53),
.Y(n_570)
);

NAND2xp33_ASAP7_75t_SL g571 ( 
.A(n_517),
.B(n_15),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_502),
.B(n_54),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_516),
.B(n_55),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_516),
.B(n_57),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_506),
.B(n_58),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_494),
.B(n_59),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_504),
.B(n_15),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_515),
.B(n_60),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_498),
.B(n_477),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_479),
.B(n_61),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_505),
.B(n_62),
.Y(n_581)
);

NAND2xp33_ASAP7_75t_SL g582 ( 
.A(n_510),
.B(n_16),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_504),
.B(n_16),
.Y(n_583)
);

INVxp67_ASAP7_75t_L g584 ( 
.A(n_541),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_543),
.B(n_490),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_537),
.A2(n_481),
.B(n_460),
.Y(n_586)
);

O2A1O1Ixp33_ASAP7_75t_SL g587 ( 
.A1(n_557),
.A2(n_519),
.B(n_508),
.C(n_507),
.Y(n_587)
);

AO21x1_ASAP7_75t_L g588 ( 
.A1(n_558),
.A2(n_520),
.B(n_499),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_543),
.Y(n_589)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_546),
.A2(n_492),
.B(n_499),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_544),
.B(n_17),
.Y(n_591)
);

AO31x2_ASAP7_75t_L g592 ( 
.A1(n_577),
.A2(n_469),
.A3(n_480),
.B(n_486),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_L g593 ( 
.A1(n_529),
.A2(n_469),
.B(n_480),
.Y(n_593)
);

NOR2xp67_ASAP7_75t_L g594 ( 
.A(n_554),
.B(n_548),
.Y(n_594)
);

AOI31xp67_ASAP7_75t_L g595 ( 
.A1(n_525),
.A2(n_486),
.A3(n_521),
.B(n_471),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_L g596 ( 
.A1(n_531),
.A2(n_471),
.B(n_521),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_578),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_SL g598 ( 
.A1(n_553),
.A2(n_64),
.B(n_63),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_575),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_566),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_583),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_579),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_559),
.B(n_18),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_L g604 ( 
.A1(n_556),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_604)
);

O2A1O1Ixp33_ASAP7_75t_SL g605 ( 
.A1(n_560),
.A2(n_157),
.B(n_223),
.C(n_222),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_524),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_578),
.B(n_20),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_534),
.A2(n_66),
.B(n_65),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_536),
.B(n_523),
.Y(n_609)
);

BUFx12f_ASAP7_75t_L g610 ( 
.A(n_535),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_528),
.A2(n_552),
.B(n_527),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_L g612 ( 
.A1(n_526),
.A2(n_69),
.B(n_68),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_545),
.B(n_22),
.Y(n_613)
);

AOI21x1_ASAP7_75t_L g614 ( 
.A1(n_550),
.A2(n_561),
.B(n_551),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_547),
.B(n_22),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_530),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_582),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_549),
.B(n_538),
.Y(n_618)
);

O2A1O1Ixp5_ASAP7_75t_L g619 ( 
.A1(n_522),
.A2(n_160),
.B(n_220),
.C(n_219),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_533),
.B(n_23),
.Y(n_620)
);

OAI21x1_ASAP7_75t_L g621 ( 
.A1(n_573),
.A2(n_71),
.B(n_70),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_539),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_540),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_532),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_574),
.A2(n_73),
.B(n_72),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_542),
.Y(n_626)
);

NAND3x1_ASAP7_75t_L g627 ( 
.A(n_565),
.B(n_24),
.C(n_25),
.Y(n_627)
);

AO21x2_ASAP7_75t_L g628 ( 
.A1(n_563),
.A2(n_76),
.B(n_75),
.Y(n_628)
);

OA21x2_ASAP7_75t_L g629 ( 
.A1(n_564),
.A2(n_78),
.B(n_77),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_555),
.B(n_24),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_L g631 ( 
.A1(n_567),
.A2(n_80),
.B(n_79),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_569),
.B(n_26),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_568),
.A2(n_571),
.B1(n_572),
.B2(n_570),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_SL g634 ( 
.A(n_580),
.B(n_81),
.Y(n_634)
);

OAI21x1_ASAP7_75t_L g635 ( 
.A1(n_576),
.A2(n_84),
.B(n_83),
.Y(n_635)
);

INVx3_ASAP7_75t_SL g636 ( 
.A(n_581),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_562),
.Y(n_637)
);

OA22x2_ASAP7_75t_L g638 ( 
.A1(n_575),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_541),
.B(n_27),
.Y(n_639)
);

OAI21x1_ASAP7_75t_L g640 ( 
.A1(n_531),
.A2(n_86),
.B(n_85),
.Y(n_640)
);

OAI21x1_ASAP7_75t_L g641 ( 
.A1(n_531),
.A2(n_88),
.B(n_87),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_529),
.B(n_29),
.Y(n_642)
);

BUFx8_ASAP7_75t_L g643 ( 
.A(n_610),
.Y(n_643)
);

OAI21x1_ASAP7_75t_L g644 ( 
.A1(n_611),
.A2(n_90),
.B(n_89),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_624),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_601),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_600),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_584),
.Y(n_648)
);

NAND3xp33_ASAP7_75t_L g649 ( 
.A(n_591),
.B(n_30),
.C(n_91),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_L g650 ( 
.A1(n_594),
.A2(n_92),
.B(n_95),
.Y(n_650)
);

OA21x2_ASAP7_75t_L g651 ( 
.A1(n_586),
.A2(n_98),
.B(n_99),
.Y(n_651)
);

BUFx2_ASAP7_75t_L g652 ( 
.A(n_597),
.Y(n_652)
);

AO31x2_ASAP7_75t_L g653 ( 
.A1(n_588),
.A2(n_102),
.A3(n_103),
.B(n_104),
.Y(n_653)
);

CKINVDCx6p67_ASAP7_75t_R g654 ( 
.A(n_636),
.Y(n_654)
);

OAI21x1_ASAP7_75t_L g655 ( 
.A1(n_614),
.A2(n_105),
.B(n_106),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_SL g656 ( 
.A(n_617),
.B(n_107),
.Y(n_656)
);

AOI221xp5_ASAP7_75t_SL g657 ( 
.A1(n_590),
.A2(n_108),
.B1(n_110),
.B2(n_111),
.C(n_113),
.Y(n_657)
);

INVx1_ASAP7_75t_SL g658 ( 
.A(n_639),
.Y(n_658)
);

NAND2x1p5_ASAP7_75t_L g659 ( 
.A(n_589),
.B(n_114),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_602),
.Y(n_660)
);

OA21x2_ASAP7_75t_L g661 ( 
.A1(n_640),
.A2(n_116),
.B(n_117),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_606),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_585),
.B(n_118),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_604),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_664)
);

NAND3xp33_ASAP7_75t_L g665 ( 
.A(n_604),
.B(n_122),
.C(n_123),
.Y(n_665)
);

OAI21x1_ASAP7_75t_L g666 ( 
.A1(n_621),
.A2(n_124),
.B(n_125),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_609),
.B(n_224),
.Y(n_667)
);

OAI21xp5_ASAP7_75t_L g668 ( 
.A1(n_594),
.A2(n_126),
.B(n_128),
.Y(n_668)
);

OAI21x1_ASAP7_75t_L g669 ( 
.A1(n_641),
.A2(n_635),
.B(n_612),
.Y(n_669)
);

CKINVDCx6p67_ASAP7_75t_R g670 ( 
.A(n_607),
.Y(n_670)
);

OR2x6_ASAP7_75t_L g671 ( 
.A(n_609),
.B(n_129),
.Y(n_671)
);

OAI22xp5_ASAP7_75t_L g672 ( 
.A1(n_596),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_672)
);

OAI21x1_ASAP7_75t_L g673 ( 
.A1(n_619),
.A2(n_133),
.B(n_134),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_616),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_603),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_626),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_622),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_642),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_622),
.Y(n_679)
);

INVx1_ASAP7_75t_SL g680 ( 
.A(n_613),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_638),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_615),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_622),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_599),
.A2(n_135),
.B1(n_137),
.B2(n_138),
.Y(n_684)
);

AOI22x1_ASAP7_75t_L g685 ( 
.A1(n_637),
.A2(n_631),
.B1(n_625),
.B2(n_618),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_596),
.B(n_139),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_593),
.B(n_592),
.Y(n_687)
);

NAND3xp33_ASAP7_75t_L g688 ( 
.A(n_593),
.B(n_141),
.C(n_143),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_630),
.B(n_620),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_623),
.Y(n_690)
);

OAI21x1_ASAP7_75t_L g691 ( 
.A1(n_631),
.A2(n_144),
.B(n_146),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_587),
.A2(n_147),
.B(n_148),
.Y(n_692)
);

INVx1_ASAP7_75t_SL g693 ( 
.A(n_632),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_648),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_687),
.B(n_675),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_644),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_660),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_647),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_676),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_666),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_653),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_672),
.A2(n_599),
.B1(n_637),
.B2(n_633),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_653),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_674),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_667),
.B(n_628),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_672),
.A2(n_633),
.B1(n_634),
.B2(n_628),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_667),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_691),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_674),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_662),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_655),
.Y(n_711)
);

OAI21x1_ASAP7_75t_SL g712 ( 
.A1(n_692),
.A2(n_668),
.B(n_650),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_678),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_651),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_669),
.Y(n_715)
);

NAND2x1p5_ASAP7_75t_L g716 ( 
.A(n_685),
.B(n_629),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_651),
.Y(n_717)
);

AO31x2_ASAP7_75t_L g718 ( 
.A1(n_692),
.A2(n_595),
.A3(n_592),
.B(n_598),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_671),
.B(n_592),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_693),
.B(n_634),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_677),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_661),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_673),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_661),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_682),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_681),
.Y(n_726)
);

OA21x2_ASAP7_75t_L g727 ( 
.A1(n_657),
.A2(n_605),
.B(n_629),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_650),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_668),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_659),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_686),
.B(n_689),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_659),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_688),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_679),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_677),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_671),
.Y(n_736)
);

INVx4_ASAP7_75t_L g737 ( 
.A(n_671),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_677),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_677),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_658),
.B(n_608),
.Y(n_740)
);

OA21x2_ASAP7_75t_L g741 ( 
.A1(n_665),
.A2(n_627),
.B(n_150),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_690),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_689),
.A2(n_149),
.B1(n_151),
.B2(n_152),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_663),
.B(n_154),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_648),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_663),
.B(n_218),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_646),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_SL g748 ( 
.A(n_654),
.B(n_656),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_645),
.Y(n_749)
);

BUFx2_ASAP7_75t_L g750 ( 
.A(n_652),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_680),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_646),
.Y(n_752)
);

OR2x2_ASAP7_75t_L g753 ( 
.A(n_670),
.B(n_155),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_R g754 ( 
.A(n_748),
.B(n_683),
.Y(n_754)
);

NAND2xp33_ASAP7_75t_R g755 ( 
.A(n_731),
.B(n_643),
.Y(n_755)
);

AND2x4_ASAP7_75t_L g756 ( 
.A(n_749),
.B(n_645),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_R g757 ( 
.A(n_749),
.B(n_643),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_749),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_731),
.B(n_649),
.Y(n_759)
);

XNOR2xp5_ASAP7_75t_L g760 ( 
.A(n_753),
.B(n_664),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_695),
.B(n_684),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_694),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_750),
.B(n_707),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_704),
.Y(n_764)
);

NAND2xp33_ASAP7_75t_R g765 ( 
.A(n_720),
.B(n_156),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_751),
.B(n_684),
.Y(n_766)
);

XNOR2xp5_ASAP7_75t_L g767 ( 
.A(n_753),
.B(n_664),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_745),
.Y(n_768)
);

INVxp67_ASAP7_75t_L g769 ( 
.A(n_745),
.Y(n_769)
);

XNOR2xp5_ASAP7_75t_L g770 ( 
.A(n_736),
.B(n_217),
.Y(n_770)
);

OR2x6_ASAP7_75t_L g771 ( 
.A(n_737),
.B(n_158),
.Y(n_771)
);

XNOR2xp5_ASAP7_75t_L g772 ( 
.A(n_744),
.B(n_162),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_704),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_707),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_709),
.Y(n_775)
);

OR2x6_ASAP7_75t_L g776 ( 
.A(n_737),
.B(n_163),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_R g777 ( 
.A(n_707),
.B(n_216),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_707),
.B(n_164),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_725),
.B(n_165),
.Y(n_779)
);

NAND2xp33_ASAP7_75t_R g780 ( 
.A(n_744),
.B(n_167),
.Y(n_780)
);

INVxp67_ASAP7_75t_L g781 ( 
.A(n_742),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_736),
.B(n_169),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_697),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_695),
.B(n_713),
.Y(n_784)
);

CKINVDCx20_ASAP7_75t_R g785 ( 
.A(n_746),
.Y(n_785)
);

NAND2xp33_ASAP7_75t_R g786 ( 
.A(n_746),
.B(n_741),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_R g787 ( 
.A(n_721),
.B(n_215),
.Y(n_787)
);

NAND2xp33_ASAP7_75t_R g788 ( 
.A(n_741),
.B(n_171),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_721),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_721),
.B(n_173),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_697),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_738),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_713),
.B(n_174),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_710),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_740),
.B(n_177),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_783),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_791),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_794),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_760),
.A2(n_767),
.B1(n_702),
.B2(n_706),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_768),
.B(n_710),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_763),
.B(n_719),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_764),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_773),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_769),
.B(n_719),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_775),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_784),
.Y(n_806)
);

OR2x6_ASAP7_75t_L g807 ( 
.A(n_771),
.B(n_776),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_762),
.B(n_699),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_759),
.B(n_719),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_777),
.B(n_728),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_758),
.B(n_719),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_781),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_758),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_761),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_766),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_793),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_756),
.B(n_785),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_779),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_789),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_774),
.B(n_708),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_792),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_782),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_757),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_795),
.B(n_698),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_770),
.B(n_735),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_771),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_776),
.B(n_708),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_786),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_772),
.B(n_698),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_772),
.B(n_735),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_778),
.B(n_708),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_788),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_790),
.Y(n_833)
);

INVxp67_ASAP7_75t_SL g834 ( 
.A(n_780),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_754),
.B(n_728),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_755),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_765),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_787),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_783),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_783),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_764),
.Y(n_841)
);

OR2x2_ASAP7_75t_L g842 ( 
.A(n_784),
.B(n_701),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_802),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_797),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_815),
.B(n_729),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_799),
.A2(n_729),
.B1(n_712),
.B2(n_733),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_797),
.Y(n_847)
);

BUFx2_ASAP7_75t_L g848 ( 
.A(n_828),
.Y(n_848)
);

OAI22xp5_ASAP7_75t_L g849 ( 
.A1(n_834),
.A2(n_743),
.B1(n_747),
.B2(n_752),
.Y(n_849)
);

INVxp67_ASAP7_75t_SL g850 ( 
.A(n_802),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_SL g851 ( 
.A1(n_834),
.A2(n_712),
.B1(n_741),
.B2(n_747),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_807),
.A2(n_733),
.B1(n_741),
.B2(n_705),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_812),
.B(n_752),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_828),
.B(n_814),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_841),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_827),
.B(n_796),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_798),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_841),
.Y(n_858)
);

INVxp67_ASAP7_75t_L g859 ( 
.A(n_806),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_796),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_798),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_839),
.Y(n_862)
);

NOR3xp33_ASAP7_75t_SL g863 ( 
.A(n_810),
.B(n_703),
.C(n_714),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_804),
.B(n_714),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_803),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_803),
.B(n_717),
.Y(n_866)
);

NAND4xp25_ASAP7_75t_L g867 ( 
.A(n_829),
.B(n_726),
.C(n_734),
.D(n_739),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_805),
.B(n_717),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_839),
.Y(n_869)
);

NOR2xp67_ASAP7_75t_L g870 ( 
.A(n_832),
.B(n_700),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_796),
.Y(n_871)
);

AOI211xp5_ASAP7_75t_L g872 ( 
.A1(n_832),
.A2(n_726),
.B(n_732),
.C(n_730),
.Y(n_872)
);

OAI221xp5_ASAP7_75t_L g873 ( 
.A1(n_810),
.A2(n_732),
.B1(n_730),
.B2(n_734),
.C(n_716),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_816),
.B(n_705),
.Y(n_874)
);

OR2x2_ASAP7_75t_L g875 ( 
.A(n_848),
.B(n_809),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_854),
.B(n_842),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_865),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_856),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_844),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_843),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_854),
.B(n_801),
.Y(n_881)
);

INVx2_ASAP7_75t_SL g882 ( 
.A(n_856),
.Y(n_882)
);

AND2x4_ASAP7_75t_SL g883 ( 
.A(n_863),
.B(n_807),
.Y(n_883)
);

NAND2xp33_ASAP7_75t_SL g884 ( 
.A(n_846),
.B(n_837),
.Y(n_884)
);

NOR2xp67_ASAP7_75t_L g885 ( 
.A(n_859),
.B(n_836),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_856),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_864),
.B(n_805),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_864),
.B(n_817),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_855),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_844),
.Y(n_890)
);

INVx1_ASAP7_75t_SL g891 ( 
.A(n_874),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_858),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_860),
.B(n_811),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_870),
.B(n_827),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_871),
.B(n_811),
.Y(n_895)
);

NAND2x1_ASAP7_75t_L g896 ( 
.A(n_847),
.B(n_807),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_845),
.B(n_816),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_853),
.B(n_818),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_850),
.B(n_857),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_857),
.B(n_840),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_888),
.B(n_823),
.Y(n_901)
);

OAI22xp33_ASAP7_75t_L g902 ( 
.A1(n_896),
.A2(n_852),
.B1(n_837),
.B2(n_873),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_891),
.B(n_851),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_885),
.B(n_898),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_897),
.B(n_846),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_880),
.B(n_861),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_889),
.B(n_861),
.Y(n_907)
);

NAND2xp33_ASAP7_75t_SL g908 ( 
.A(n_875),
.B(n_823),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_884),
.A2(n_826),
.B1(n_867),
.B2(n_827),
.Y(n_909)
);

CKINVDCx20_ASAP7_75t_R g910 ( 
.A(n_884),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_892),
.B(n_862),
.Y(n_911)
);

OAI22xp33_ASAP7_75t_L g912 ( 
.A1(n_882),
.A2(n_835),
.B1(n_849),
.B2(n_838),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_887),
.B(n_862),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_887),
.B(n_869),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_899),
.B(n_869),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_906),
.Y(n_916)
);

AOI222xp33_ASAP7_75t_L g917 ( 
.A1(n_910),
.A2(n_905),
.B1(n_902),
.B2(n_903),
.C1(n_912),
.C2(n_883),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_904),
.B(n_878),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_907),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_911),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_915),
.B(n_877),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_913),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_901),
.B(n_878),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_914),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_909),
.B(n_882),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_908),
.B(n_886),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_917),
.B(n_894),
.Y(n_927)
);

NAND3xp33_ASAP7_75t_L g928 ( 
.A(n_917),
.B(n_872),
.C(n_824),
.Y(n_928)
);

AOI21xp33_ASAP7_75t_L g929 ( 
.A1(n_916),
.A2(n_821),
.B(n_819),
.Y(n_929)
);

OAI21xp33_ASAP7_75t_SL g930 ( 
.A1(n_926),
.A2(n_886),
.B(n_881),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_918),
.B(n_893),
.Y(n_931)
);

OR2x2_ASAP7_75t_L g932 ( 
.A(n_924),
.B(n_876),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_919),
.B(n_881),
.Y(n_933)
);

OAI32xp33_ASAP7_75t_L g934 ( 
.A1(n_925),
.A2(n_838),
.A3(n_900),
.B1(n_895),
.B2(n_893),
.Y(n_934)
);

OAI22xp33_ASAP7_75t_L g935 ( 
.A1(n_928),
.A2(n_922),
.B1(n_920),
.B2(n_921),
.Y(n_935)
);

AOI22xp33_ASAP7_75t_L g936 ( 
.A1(n_927),
.A2(n_922),
.B1(n_923),
.B2(n_883),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_933),
.A2(n_921),
.B1(n_894),
.B2(n_895),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_929),
.B(n_894),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_931),
.B(n_830),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_935),
.B(n_932),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_939),
.Y(n_941)
);

INVxp33_ASAP7_75t_SL g942 ( 
.A(n_936),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_938),
.B(n_930),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_937),
.Y(n_944)
);

NOR3xp33_ASAP7_75t_L g945 ( 
.A(n_940),
.B(n_934),
.C(n_808),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_941),
.B(n_825),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_944),
.B(n_879),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_943),
.B(n_879),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_942),
.B(n_890),
.Y(n_949)
);

NAND3xp33_ASAP7_75t_SL g950 ( 
.A(n_940),
.B(n_813),
.C(n_822),
.Y(n_950)
);

AOI221xp5_ASAP7_75t_L g951 ( 
.A1(n_945),
.A2(n_950),
.B1(n_949),
.B2(n_948),
.C(n_947),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_946),
.Y(n_952)
);

XNOR2x1_ASAP7_75t_L g953 ( 
.A(n_946),
.B(n_820),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_949),
.Y(n_954)
);

AO22x1_ASAP7_75t_L g955 ( 
.A1(n_954),
.A2(n_952),
.B1(n_951),
.B2(n_953),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_952),
.Y(n_956)
);

AND3x4_ASAP7_75t_L g957 ( 
.A(n_954),
.B(n_811),
.C(n_820),
.Y(n_957)
);

XOR2xp5_ASAP7_75t_L g958 ( 
.A(n_954),
.B(n_833),
.Y(n_958)
);

NAND4xp75_ASAP7_75t_L g959 ( 
.A(n_952),
.B(n_800),
.C(n_868),
.D(n_866),
.Y(n_959)
);

NAND2xp33_ASAP7_75t_SL g960 ( 
.A(n_957),
.B(n_833),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_956),
.B(n_958),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_R g962 ( 
.A(n_959),
.B(n_180),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_955),
.B(n_868),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_R g964 ( 
.A(n_956),
.B(n_181),
.Y(n_964)
);

XNOR2x1_ASAP7_75t_L g965 ( 
.A(n_955),
.B(n_182),
.Y(n_965)
);

AOI22xp5_ASAP7_75t_L g966 ( 
.A1(n_960),
.A2(n_831),
.B1(n_820),
.B2(n_705),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_965),
.A2(n_831),
.B(n_723),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_964),
.B(n_831),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_963),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_962),
.Y(n_970)
);

OR2x2_ASAP7_75t_L g971 ( 
.A(n_961),
.B(n_718),
.Y(n_971)
);

XNOR2xp5_ASAP7_75t_L g972 ( 
.A(n_965),
.B(n_183),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_970),
.A2(n_696),
.B1(n_711),
.B2(n_700),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_969),
.B(n_184),
.Y(n_974)
);

INVx1_ASAP7_75t_SL g975 ( 
.A(n_972),
.Y(n_975)
);

NOR3xp33_ASAP7_75t_L g976 ( 
.A(n_968),
.B(n_696),
.C(n_711),
.Y(n_976)
);

OAI21xp5_ASAP7_75t_L g977 ( 
.A1(n_967),
.A2(n_724),
.B(n_722),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_971),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_974),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_975),
.B(n_966),
.Y(n_980)
);

CKINVDCx20_ASAP7_75t_R g981 ( 
.A(n_978),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_L g982 ( 
.A1(n_981),
.A2(n_976),
.B1(n_977),
.B2(n_973),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_L g983 ( 
.A1(n_979),
.A2(n_727),
.B1(n_715),
.B2(n_187),
.Y(n_983)
);

XNOR2xp5_ASAP7_75t_L g984 ( 
.A(n_982),
.B(n_980),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_984),
.Y(n_985)
);

AOI222xp33_ASAP7_75t_L g986 ( 
.A1(n_984),
.A2(n_983),
.B1(n_715),
.B2(n_190),
.C1(n_191),
.C2(n_194),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_985),
.Y(n_987)
);

AOI221xp5_ASAP7_75t_L g988 ( 
.A1(n_987),
.A2(n_986),
.B1(n_189),
.B2(n_195),
.C(n_198),
.Y(n_988)
);

AOI211xp5_ASAP7_75t_L g989 ( 
.A1(n_988),
.A2(n_201),
.B(n_202),
.C(n_203),
.Y(n_989)
);


endmodule