module real_aes_1800_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_733;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g525 ( .A(n_0), .B(n_222), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_1), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g156 ( .A(n_2), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_3), .B(n_528), .Y(n_547) );
NAND2xp33_ASAP7_75t_SL g518 ( .A(n_4), .B(n_177), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_5), .B(n_190), .Y(n_213) );
INVx1_ASAP7_75t_L g510 ( .A(n_6), .Y(n_510) );
INVx1_ASAP7_75t_L g247 ( .A(n_7), .Y(n_247) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_8), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_9), .Y(n_264) );
AND2x2_ASAP7_75t_L g545 ( .A(n_10), .B(n_146), .Y(n_545) );
AOI22xp33_ASAP7_75t_SL g798 ( .A1(n_11), .A2(n_792), .B1(n_799), .B2(n_801), .Y(n_798) );
INVx2_ASAP7_75t_L g147 ( .A(n_12), .Y(n_147) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_13), .Y(n_114) );
INVx1_ASAP7_75t_L g223 ( .A(n_14), .Y(n_223) );
AOI221x1_ASAP7_75t_L g513 ( .A1(n_15), .A2(n_179), .B1(n_514), .B2(n_516), .C(n_517), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_16), .B(n_528), .Y(n_581) );
INVx1_ASAP7_75t_L g110 ( .A(n_17), .Y(n_110) );
INVx1_ASAP7_75t_L g220 ( .A(n_18), .Y(n_220) );
INVx1_ASAP7_75t_SL g168 ( .A(n_19), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_20), .B(n_171), .Y(n_193) );
AOI33xp33_ASAP7_75t_L g238 ( .A1(n_21), .A2(n_49), .A3(n_153), .B1(n_164), .B2(n_239), .B3(n_240), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_22), .A2(n_516), .B(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_23), .B(n_222), .Y(n_550) );
AOI221xp5_ASAP7_75t_SL g590 ( .A1(n_24), .A2(n_40), .B1(n_516), .B2(n_528), .C(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g257 ( .A(n_25), .Y(n_257) );
OR2x2_ASAP7_75t_L g148 ( .A(n_26), .B(n_91), .Y(n_148) );
OA21x2_ASAP7_75t_L g181 ( .A1(n_26), .A2(n_91), .B(n_147), .Y(n_181) );
INVxp67_ASAP7_75t_L g512 ( .A(n_27), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_28), .B(n_225), .Y(n_585) );
AND2x2_ASAP7_75t_L g539 ( .A(n_29), .B(n_145), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_30), .B(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_31), .A2(n_516), .B(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_32), .B(n_225), .Y(n_592) );
AND2x2_ASAP7_75t_L g158 ( .A(n_33), .B(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g163 ( .A(n_33), .Y(n_163) );
AND2x2_ASAP7_75t_L g177 ( .A(n_33), .B(n_156), .Y(n_177) );
NOR3xp33_ASAP7_75t_L g111 ( .A(n_34), .B(n_112), .C(n_114), .Y(n_111) );
OR2x6_ASAP7_75t_L g128 ( .A(n_34), .B(n_129), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g259 ( .A(n_35), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g827 ( .A(n_36), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_37), .B(n_151), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_38), .A2(n_180), .B1(n_186), .B2(n_190), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_39), .B(n_195), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_41), .A2(n_83), .B1(n_161), .B2(n_516), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_42), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_43), .B(n_222), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_44), .B(n_197), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_45), .B(n_171), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_46), .Y(n_189) );
AND2x2_ASAP7_75t_L g529 ( .A(n_47), .B(n_145), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_48), .B(n_145), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_50), .B(n_171), .Y(n_288) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_51), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g816 ( .A1(n_51), .A2(n_63), .B1(n_436), .B2(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g154 ( .A(n_52), .Y(n_154) );
INVx1_ASAP7_75t_L g173 ( .A(n_52), .Y(n_173) );
AOI22x1_ASAP7_75t_L g792 ( .A1(n_53), .A2(n_793), .B1(n_794), .B2(n_795), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_53), .Y(n_793) );
AND2x2_ASAP7_75t_L g289 ( .A(n_54), .B(n_145), .Y(n_289) );
AOI221xp5_ASAP7_75t_L g245 ( .A1(n_55), .A2(n_76), .B1(n_151), .B2(n_161), .C(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_56), .B(n_151), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_57), .B(n_528), .Y(n_538) );
OAI21xp5_ASAP7_75t_L g803 ( .A1(n_58), .A2(n_804), .B(n_819), .Y(n_803) );
INVx1_ASAP7_75t_L g822 ( .A(n_58), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_59), .B(n_180), .Y(n_266) );
AOI21xp5_ASAP7_75t_SL g202 ( .A1(n_60), .A2(n_161), .B(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g566 ( .A(n_61), .B(n_145), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_62), .B(n_225), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_63), .Y(n_817) );
INVx1_ASAP7_75t_L g216 ( .A(n_64), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_65), .B(n_222), .Y(n_564) );
AND2x2_ASAP7_75t_SL g586 ( .A(n_66), .B(n_146), .Y(n_586) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_67), .A2(n_516), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g287 ( .A(n_68), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_69), .B(n_225), .Y(n_551) );
AND2x2_ASAP7_75t_SL g558 ( .A(n_70), .B(n_197), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_71), .A2(n_103), .B1(n_796), .B2(n_797), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_71), .Y(n_796) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_72), .A2(n_161), .B(n_286), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_73), .A2(n_815), .B1(n_816), .B2(n_818), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_73), .Y(n_815) );
INVx1_ASAP7_75t_L g159 ( .A(n_74), .Y(n_159) );
INVx1_ASAP7_75t_L g175 ( .A(n_74), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_75), .B(n_151), .Y(n_241) );
AND2x2_ASAP7_75t_L g178 ( .A(n_77), .B(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g217 ( .A(n_78), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_79), .A2(n_161), .B(n_167), .Y(n_160) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_80), .A2(n_161), .B(n_192), .C(n_196), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_81), .A2(n_86), .B1(n_151), .B2(n_528), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_82), .B(n_528), .Y(n_565) );
INVx1_ASAP7_75t_L g109 ( .A(n_84), .Y(n_109) );
AND2x2_ASAP7_75t_SL g200 ( .A(n_85), .B(n_179), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g235 ( .A1(n_87), .A2(n_161), .B1(n_236), .B2(n_237), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_88), .B(n_222), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_89), .B(n_222), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_90), .A2(n_516), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g204 ( .A(n_92), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_93), .B(n_225), .Y(n_563) );
AND2x2_ASAP7_75t_L g242 ( .A(n_94), .B(n_179), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_95), .A2(n_255), .B(n_256), .C(n_258), .Y(n_254) );
INVxp67_ASAP7_75t_L g515 ( .A(n_96), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_97), .B(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_98), .B(n_225), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_99), .A2(n_516), .B(n_583), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_100), .Y(n_124) );
BUFx2_ASAP7_75t_L g120 ( .A(n_101), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_102), .B(n_171), .Y(n_205) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_103), .Y(n_797) );
AOI21xp33_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_115), .B(n_826), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g828 ( .A(n_106), .Y(n_828) );
INVx3_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_SL g107 ( .A(n_108), .B(n_111), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_109), .B(n_110), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_114), .B(n_127), .Y(n_126) );
AND2x6_ASAP7_75t_SL g500 ( .A(n_114), .B(n_128), .Y(n_500) );
OR2x6_ASAP7_75t_SL g791 ( .A(n_114), .B(n_127), .Y(n_791) );
OR2x2_ASAP7_75t_L g802 ( .A(n_114), .B(n_128), .Y(n_802) );
OA22x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_130), .B1(n_803), .B2(n_824), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_121), .Y(n_116) );
CKINVDCx11_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
BUFx3_ASAP7_75t_L g825 ( .A(n_118), .Y(n_825) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g121 ( .A(n_122), .Y(n_121) );
HB1xp67_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g819 ( .A1(n_123), .A2(n_820), .B(n_821), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
INVx1_ASAP7_75t_L g823 ( .A(n_125), .Y(n_823) );
BUFx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
BUFx3_ASAP7_75t_L g807 ( .A(n_126), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_128), .Y(n_127) );
OAI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_792), .B(n_798), .Y(n_130) );
INVxp67_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
OAI22x1_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_499), .B1(n_501), .B2(n_789), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OAI22xp5_ASAP7_75t_L g799 ( .A1(n_134), .A2(n_499), .B1(n_502), .B2(n_800), .Y(n_799) );
AND3x1_ASAP7_75t_L g134 ( .A(n_135), .B(n_493), .C(n_496), .Y(n_134) );
NAND5xp2_ASAP7_75t_L g135 ( .A(n_136), .B(n_393), .C(n_423), .D(n_437), .E(n_463), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OAI21xp33_ASAP7_75t_L g493 ( .A1(n_137), .A2(n_436), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g811 ( .A(n_137), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_342), .Y(n_137) );
NOR3xp33_ASAP7_75t_SL g138 ( .A(n_139), .B(n_290), .C(n_324), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_207), .B(n_229), .C(n_268), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_182), .Y(n_140) );
BUFx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_142), .B(n_280), .Y(n_345) );
AND2x2_ASAP7_75t_L g432 ( .A(n_142), .B(n_210), .Y(n_432) );
HB1xp67_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
OR2x2_ASAP7_75t_L g228 ( .A(n_143), .B(n_199), .Y(n_228) );
INVx1_ASAP7_75t_L g270 ( .A(n_143), .Y(n_270) );
INVx2_ASAP7_75t_L g275 ( .A(n_143), .Y(n_275) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_143), .Y(n_303) );
INVx1_ASAP7_75t_L g317 ( .A(n_143), .Y(n_317) );
AND2x2_ASAP7_75t_L g321 ( .A(n_143), .B(n_212), .Y(n_321) );
AND2x2_ASAP7_75t_L g402 ( .A(n_143), .B(n_211), .Y(n_402) );
AO21x2_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_149), .B(n_178), .Y(n_143) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_144), .A2(n_533), .B(n_539), .Y(n_532) );
AO21x2_ASAP7_75t_L g559 ( .A1(n_144), .A2(n_560), .B(n_566), .Y(n_559) );
AO21x2_ASAP7_75t_L g597 ( .A1(n_144), .A2(n_533), .B(n_539), .Y(n_597) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_145), .Y(n_144) );
OA21x2_ASAP7_75t_L g589 ( .A1(n_145), .A2(n_590), .B(n_594), .Y(n_589) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_SL g146 ( .A(n_147), .B(n_148), .Y(n_146) );
AND2x4_ASAP7_75t_L g190 ( .A(n_147), .B(n_148), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_150), .B(n_160), .Y(n_149) );
INVx1_ASAP7_75t_L g267 ( .A(n_151), .Y(n_267) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_151), .A2(n_161), .B1(n_509), .B2(n_511), .Y(n_508) );
AND2x4_ASAP7_75t_L g151 ( .A(n_152), .B(n_157), .Y(n_151) );
INVx1_ASAP7_75t_L g187 ( .A(n_152), .Y(n_187) );
AND2x2_ASAP7_75t_L g152 ( .A(n_153), .B(n_155), .Y(n_152) );
OR2x6_ASAP7_75t_L g169 ( .A(n_153), .B(n_165), .Y(n_169) );
INVxp33_ASAP7_75t_L g239 ( .A(n_153), .Y(n_239) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_L g166 ( .A(n_154), .B(n_156), .Y(n_166) );
AND2x4_ASAP7_75t_L g225 ( .A(n_154), .B(n_174), .Y(n_225) );
HB1xp67_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g188 ( .A(n_157), .Y(n_188) );
BUFx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AND2x6_ASAP7_75t_L g516 ( .A(n_158), .B(n_166), .Y(n_516) );
INVx2_ASAP7_75t_L g165 ( .A(n_159), .Y(n_165) );
AND2x6_ASAP7_75t_L g222 ( .A(n_159), .B(n_172), .Y(n_222) );
INVxp67_ASAP7_75t_L g265 ( .A(n_161), .Y(n_265) );
AND2x4_ASAP7_75t_L g161 ( .A(n_162), .B(n_166), .Y(n_161) );
NOR2x1p5_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
INVx1_ASAP7_75t_L g240 ( .A(n_164), .Y(n_240) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
O2A1O1Ixp33_ASAP7_75t_SL g167 ( .A1(n_168), .A2(n_169), .B(n_170), .C(n_176), .Y(n_167) );
INVx2_ASAP7_75t_L g195 ( .A(n_169), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_L g203 ( .A1(n_169), .A2(n_176), .B(n_204), .C(n_205), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g215 ( .A1(n_169), .A2(n_216), .B1(n_217), .B2(n_218), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_SL g246 ( .A1(n_169), .A2(n_176), .B(n_247), .C(n_248), .Y(n_246) );
INVxp67_ASAP7_75t_L g255 ( .A(n_169), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_L g286 ( .A1(n_169), .A2(n_176), .B(n_287), .C(n_288), .Y(n_286) );
INVx1_ASAP7_75t_L g218 ( .A(n_171), .Y(n_218) );
AND2x4_ASAP7_75t_L g528 ( .A(n_171), .B(n_177), .Y(n_528) );
AND2x4_ASAP7_75t_L g171 ( .A(n_172), .B(n_174), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_176), .A2(n_193), .B(n_194), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_176), .B(n_190), .Y(n_226) );
INVx1_ASAP7_75t_L g236 ( .A(n_176), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_176), .A2(n_525), .B(n_526), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_176), .A2(n_536), .B(n_537), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_176), .A2(n_550), .B(n_551), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_176), .A2(n_563), .B(n_564), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g583 ( .A1(n_176), .A2(n_584), .B(n_585), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g591 ( .A1(n_176), .A2(n_592), .B(n_593), .Y(n_591) );
INVx5_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_177), .Y(n_258) );
OAI22xp5_ASAP7_75t_L g253 ( .A1(n_179), .A2(n_254), .B1(n_259), .B2(n_260), .Y(n_253) );
INVx3_ASAP7_75t_L g260 ( .A(n_179), .Y(n_260) );
INVx4_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_180), .B(n_263), .Y(n_262) );
AOI21x1_ASAP7_75t_L g521 ( .A1(n_180), .A2(n_522), .B(n_529), .Y(n_521) );
INVx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
BUFx4f_ASAP7_75t_L g197 ( .A(n_181), .Y(n_197) );
AND2x4_ASAP7_75t_SL g182 ( .A(n_183), .B(n_198), .Y(n_182) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g227 ( .A(n_184), .Y(n_227) );
AND2x2_ASAP7_75t_L g271 ( .A(n_184), .B(n_212), .Y(n_271) );
AND2x2_ASAP7_75t_L g292 ( .A(n_184), .B(n_199), .Y(n_292) );
INVx1_ASAP7_75t_L g315 ( .A(n_184), .Y(n_315) );
AND2x4_ASAP7_75t_L g382 ( .A(n_184), .B(n_211), .Y(n_382) );
AND2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_191), .Y(n_184) );
NOR3xp33_ASAP7_75t_L g186 ( .A(n_187), .B(n_188), .C(n_189), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_190), .A2(n_202), .B(n_206), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_190), .B(n_510), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_190), .B(n_512), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_190), .B(n_515), .Y(n_514) );
NOR3xp33_ASAP7_75t_L g517 ( .A(n_190), .B(n_218), .C(n_518), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_190), .A2(n_547), .B(n_548), .Y(n_546) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_196), .A2(n_234), .B(n_242), .Y(n_233) );
AO21x2_ASAP7_75t_L g297 ( .A1(n_196), .A2(n_234), .B(n_242), .Y(n_297) );
AOI21x1_ASAP7_75t_L g554 ( .A1(n_196), .A2(n_555), .B(n_558), .Y(n_554) );
INVx2_ASAP7_75t_SL g196 ( .A(n_197), .Y(n_196) );
OA21x2_ASAP7_75t_L g244 ( .A1(n_197), .A2(n_245), .B(n_249), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_197), .A2(n_581), .B(n_582), .Y(n_580) );
AND2x4_ASAP7_75t_L g398 ( .A(n_198), .B(n_315), .Y(n_398) );
OR2x2_ASAP7_75t_L g439 ( .A(n_198), .B(n_440), .Y(n_439) );
NOR2xp67_ASAP7_75t_SL g458 ( .A(n_198), .B(n_331), .Y(n_458) );
NOR2x1_ASAP7_75t_L g476 ( .A(n_198), .B(n_390), .Y(n_476) );
INVx4_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NOR2x1_ASAP7_75t_SL g276 ( .A(n_199), .B(n_212), .Y(n_276) );
AND2x4_ASAP7_75t_L g314 ( .A(n_199), .B(n_315), .Y(n_314) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_199), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_199), .B(n_274), .Y(n_352) );
INVx2_ASAP7_75t_L g366 ( .A(n_199), .Y(n_366) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_199), .B(n_318), .Y(n_388) );
AND2x2_ASAP7_75t_L g480 ( .A(n_199), .B(n_338), .Y(n_480) );
OR2x6_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NOR2x1_ASAP7_75t_L g208 ( .A(n_209), .B(n_228), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_210), .B(n_317), .Y(n_331) );
AND2x2_ASAP7_75t_SL g340 ( .A(n_210), .B(n_320), .Y(n_340) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_227), .Y(n_210) );
INVx1_ASAP7_75t_L g318 ( .A(n_211), .Y(n_318) );
INVx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g338 ( .A(n_212), .Y(n_338) );
AND2x4_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
OAI21xp5_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_219), .B(n_226), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_218), .B(n_257), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B1(n_223), .B2(n_224), .Y(n_219) );
INVxp67_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVxp67_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g371 ( .A(n_227), .Y(n_371) );
INVx2_ASAP7_75t_SL g416 ( .A(n_228), .Y(n_416) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_250), .Y(n_230) );
NAND2x1p5_ASAP7_75t_L g325 ( .A(n_231), .B(n_326), .Y(n_325) );
BUFx2_ASAP7_75t_L g362 ( .A(n_231), .Y(n_362) );
AND2x2_ASAP7_75t_L g486 ( .A(n_231), .B(n_311), .Y(n_486) );
AND2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_243), .Y(n_231) );
AND2x4_ASAP7_75t_L g299 ( .A(n_232), .B(n_281), .Y(n_299) );
INVx1_ASAP7_75t_L g310 ( .A(n_232), .Y(n_310) );
AND2x2_ASAP7_75t_L g341 ( .A(n_232), .B(n_296), .Y(n_341) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_233), .B(n_244), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_233), .B(n_282), .Y(n_373) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_235), .B(n_241), .Y(n_234) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVxp67_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g279 ( .A(n_244), .Y(n_279) );
AND2x4_ASAP7_75t_L g347 ( .A(n_244), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g359 ( .A(n_244), .Y(n_359) );
INVx1_ASAP7_75t_L g401 ( .A(n_244), .Y(n_401) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_244), .Y(n_413) );
AND2x2_ASAP7_75t_L g429 ( .A(n_244), .B(n_252), .Y(n_429) );
BUFx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g376 ( .A(n_251), .B(n_334), .Y(n_376) );
INVx1_ASAP7_75t_SL g378 ( .A(n_251), .Y(n_378) );
AND2x2_ASAP7_75t_L g399 ( .A(n_251), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x4_ASAP7_75t_L g278 ( .A(n_252), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g306 ( .A(n_252), .Y(n_306) );
INVx2_ASAP7_75t_L g312 ( .A(n_252), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_252), .B(n_282), .Y(n_327) );
OR2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_261), .Y(n_252) );
AO21x2_ASAP7_75t_L g282 ( .A1(n_260), .A2(n_283), .B(n_289), .Y(n_282) );
AO21x2_ASAP7_75t_L g296 ( .A1(n_260), .A2(n_283), .B(n_289), .Y(n_296) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_265), .B1(n_266), .B2(n_267), .Y(n_261) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OAI21xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_272), .B(n_277), .Y(n_268) );
INVx1_ASAP7_75t_L g408 ( .A(n_269), .Y(n_408) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx2_ASAP7_75t_L g328 ( .A(n_271), .Y(n_328) );
AND2x2_ASAP7_75t_L g384 ( .A(n_271), .B(n_320), .Y(n_384) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_276), .Y(n_272) );
INVx1_ASAP7_75t_L g298 ( .A(n_273), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_273), .B(n_314), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_273), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g405 ( .A(n_273), .B(n_398), .Y(n_405) );
AND2x2_ASAP7_75t_L g479 ( .A(n_273), .B(n_480), .Y(n_479) );
INVx3_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_274), .Y(n_467) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_275), .Y(n_387) );
AND2x2_ASAP7_75t_L g300 ( .A(n_276), .B(n_301), .Y(n_300) );
OAI21xp33_ASAP7_75t_L g488 ( .A1(n_276), .A2(n_489), .B(n_491), .Y(n_488) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
INVx3_ASAP7_75t_L g374 ( .A(n_278), .Y(n_374) );
NAND2x1_ASAP7_75t_SL g418 ( .A(n_278), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g421 ( .A(n_278), .B(n_299), .Y(n_421) );
AND2x2_ASAP7_75t_L g333 ( .A(n_280), .B(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g470 ( .A(n_280), .B(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g481 ( .A(n_280), .B(n_429), .Y(n_481) );
INVx3_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2x1p5_ASAP7_75t_L g357 ( .A(n_281), .B(n_358), .Y(n_357) );
INVx3_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g412 ( .A(n_282), .B(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
OAI21xp5_ASAP7_75t_SL g290 ( .A1(n_291), .A2(n_304), .B(n_307), .Y(n_290) );
AOI22xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_293), .B1(n_299), .B2(n_300), .Y(n_291) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_292), .Y(n_349) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_298), .Y(n_293) );
AND2x2_ASAP7_75t_L g322 ( .A(n_294), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g428 ( .A(n_294), .B(n_429), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_294), .A2(n_447), .B1(n_448), .B2(n_449), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_294), .B(n_455), .Y(n_454) );
AND2x4_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g311 ( .A(n_296), .B(n_312), .Y(n_311) );
NOR2xp67_ASAP7_75t_L g392 ( .A(n_296), .B(n_312), .Y(n_392) );
NOR2x1_ASAP7_75t_L g400 ( .A(n_296), .B(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g348 ( .A(n_297), .Y(n_348) );
AND2x2_ASAP7_75t_L g356 ( .A(n_297), .B(n_312), .Y(n_356) );
INVx1_ASAP7_75t_L g419 ( .A(n_297), .Y(n_419) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2x1_ASAP7_75t_L g337 ( .A(n_302), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g449 ( .A(n_305), .B(n_334), .Y(n_449) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g323 ( .A(n_306), .Y(n_323) );
AND2x2_ASAP7_75t_L g346 ( .A(n_306), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g434 ( .A(n_306), .B(n_341), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_313), .B1(n_319), .B2(n_322), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g442 ( .A(n_309), .B(n_443), .Y(n_442) );
NAND2x1p5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
AND2x2_ASAP7_75t_L g472 ( .A(n_312), .B(n_359), .Y(n_472) );
AND2x2_ASAP7_75t_SL g313 ( .A(n_314), .B(n_316), .Y(n_313) );
INVx2_ASAP7_75t_L g339 ( .A(n_314), .Y(n_339) );
OAI21xp33_ASAP7_75t_SL g485 ( .A1(n_314), .A2(n_486), .B(n_487), .Y(n_485) );
AND2x4_ASAP7_75t_SL g316 ( .A(n_317), .B(n_318), .Y(n_316) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_317), .Y(n_475) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
O2A1O1Ixp33_ASAP7_75t_SL g417 ( .A1(n_320), .A2(n_418), .B(n_420), .C(n_422), .Y(n_417) );
AND2x2_ASAP7_75t_SL g369 ( .A(n_321), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g422 ( .A(n_321), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_321), .B(n_398), .Y(n_462) );
INVx1_ASAP7_75t_SL g329 ( .A(n_322), .Y(n_329) );
AND2x2_ASAP7_75t_L g410 ( .A(n_323), .B(n_347), .Y(n_410) );
INVx1_ASAP7_75t_L g455 ( .A(n_323), .Y(n_455) );
OAI221xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_328), .B1(n_329), .B2(n_330), .C(n_332), .Y(n_324) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_325), .Y(n_444) );
INVx2_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g492 ( .A(n_327), .B(n_335), .Y(n_492) );
OR2x2_ASAP7_75t_L g351 ( .A(n_328), .B(n_352), .Y(n_351) );
NOR2x1_ASAP7_75t_L g364 ( .A(n_328), .B(n_365), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_328), .B(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g490 ( .A(n_328), .B(n_387), .Y(n_490) );
BUFx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AOI32xp33_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_336), .A3(n_339), .B1(n_340), .B2(n_341), .Y(n_332) );
INVx1_ASAP7_75t_L g353 ( .A(n_334), .Y(n_353) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_336), .B(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g448 ( .A(n_337), .Y(n_448) );
OAI22xp33_ASAP7_75t_SL g430 ( .A1(n_339), .A2(n_431), .B1(n_433), .B2(n_435), .Y(n_430) );
INVx1_ASAP7_75t_L g461 ( .A(n_340), .Y(n_461) );
AOI211x1_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_349), .B(n_350), .C(n_367), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_344), .B(n_429), .Y(n_435) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_L g391 ( .A(n_347), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g457 ( .A(n_347), .Y(n_457) );
OAI222xp33_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_353), .B1(n_354), .B2(n_360), .C1(n_361), .C2(n_363), .Y(n_350) );
INVxp67_ASAP7_75t_L g447 ( .A(n_351), .Y(n_447) );
OR2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_357), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_355), .B(n_440), .Y(n_487) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g403 ( .A(n_356), .B(n_400), .Y(n_403) );
INVx3_ASAP7_75t_L g443 ( .A(n_358), .Y(n_443) );
BUFx3_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g381 ( .A(n_366), .B(n_382), .Y(n_381) );
OAI221xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_372), .B1(n_375), .B2(n_380), .C(n_383), .Y(n_367) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
OAI21xp5_ASAP7_75t_L g425 ( .A1(n_369), .A2(n_426), .B(n_428), .Y(n_425) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
OR2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVx1_ASAP7_75t_L g379 ( .A(n_373), .Y(n_379) );
OR2x2_ASAP7_75t_L g483 ( .A(n_374), .B(n_419), .Y(n_483) );
NOR2xp67_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_377), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
OAI21xp5_ASAP7_75t_L g477 ( .A1(n_380), .A2(n_409), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OAI21xp5_ASAP7_75t_L g459 ( .A1(n_381), .A2(n_453), .B(n_460), .Y(n_459) );
INVx4_ASAP7_75t_L g390 ( .A(n_382), .Y(n_390) );
OAI31xp33_ASAP7_75t_SL g383 ( .A1(n_384), .A2(n_385), .A3(n_389), .B(n_391), .Y(n_383) );
INVx1_ASAP7_75t_L g441 ( .A(n_385), .Y(n_441) );
NOR2x1_ASAP7_75t_L g385 ( .A(n_386), .B(n_388), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g415 ( .A(n_390), .Y(n_415) );
AND2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_406), .Y(n_393) );
NAND4xp25_ASAP7_75t_L g494 ( .A(n_394), .B(n_406), .C(n_425), .D(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_404), .Y(n_394) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_399), .B1(n_402), .B2(n_403), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g466 ( .A(n_398), .B(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_399), .B(n_419), .Y(n_427) );
INVx1_ASAP7_75t_SL g440 ( .A(n_402), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_407), .B(n_417), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .B1(n_411), .B2(n_414), .Y(n_407) );
INVx3_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVxp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NAND2x1_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_416), .A2(n_479), .B1(n_481), .B2(n_482), .Y(n_478) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NOR3xp33_ASAP7_75t_L g423 ( .A(n_424), .B(n_430), .C(n_436), .Y(n_423) );
INVxp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g495 ( .A(n_430), .Y(n_495) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI21xp33_ASAP7_75t_L g496 ( .A1(n_436), .A2(n_497), .B(n_498), .Y(n_496) );
INVxp33_ASAP7_75t_L g497 ( .A(n_437), .Y(n_497) );
AND2x2_ASAP7_75t_L g810 ( .A(n_437), .B(n_463), .Y(n_810) );
NOR2xp67_ASAP7_75t_L g437 ( .A(n_438), .B(n_445), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_441), .B1(n_442), .B2(n_444), .Y(n_438) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_442), .A2(n_465), .B(n_468), .Y(n_464) );
INVx2_ASAP7_75t_L g452 ( .A(n_443), .Y(n_452) );
NAND3xp33_ASAP7_75t_SL g445 ( .A(n_446), .B(n_450), .C(n_459), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_453), .B1(n_456), .B2(n_458), .Y(n_450) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
INVxp33_ASAP7_75t_SL g498 ( .A(n_463), .Y(n_498) );
NOR3x1_ASAP7_75t_L g463 ( .A(n_464), .B(n_477), .C(n_484), .Y(n_463) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_473), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_485), .B(n_488), .Y(n_484) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g812 ( .A(n_494), .Y(n_812) );
CKINVDCx11_ASAP7_75t_R g499 ( .A(n_500), .Y(n_499) );
INVx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_503), .B(n_666), .Y(n_502) );
NOR4xp25_ASAP7_75t_L g503 ( .A(n_504), .B(n_609), .C(n_648), .D(n_655), .Y(n_503) );
OAI221xp5_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_530), .B1(n_567), .B2(n_576), .C(n_595), .Y(n_504) );
OR2x2_ASAP7_75t_L g739 ( .A(n_505), .B(n_601), .Y(n_739) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g654 ( .A(n_506), .B(n_579), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_506), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_SL g719 ( .A(n_506), .B(n_720), .Y(n_719) );
AND2x4_ASAP7_75t_L g506 ( .A(n_507), .B(n_519), .Y(n_506) );
AND2x4_ASAP7_75t_SL g578 ( .A(n_507), .B(n_579), .Y(n_578) );
INVx3_ASAP7_75t_L g600 ( .A(n_507), .Y(n_600) );
AND2x2_ASAP7_75t_L g635 ( .A(n_507), .B(n_608), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_507), .B(n_520), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_507), .B(n_602), .Y(n_687) );
OR2x2_ASAP7_75t_L g765 ( .A(n_507), .B(n_579), .Y(n_765) );
AND2x4_ASAP7_75t_L g507 ( .A(n_508), .B(n_513), .Y(n_507) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g587 ( .A(n_520), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_520), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g613 ( .A(n_520), .Y(n_613) );
OR2x2_ASAP7_75t_L g618 ( .A(n_520), .B(n_602), .Y(n_618) );
AND2x2_ASAP7_75t_L g631 ( .A(n_520), .B(n_589), .Y(n_631) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_520), .Y(n_634) );
INVx1_ASAP7_75t_L g646 ( .A(n_520), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_520), .B(n_600), .Y(n_711) );
INVx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_527), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_531), .B(n_540), .Y(n_530) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
OR2x2_ASAP7_75t_L g575 ( .A(n_532), .B(n_559), .Y(n_575) );
AND2x4_ASAP7_75t_L g605 ( .A(n_532), .B(n_544), .Y(n_605) );
INVx2_ASAP7_75t_L g639 ( .A(n_532), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_532), .B(n_559), .Y(n_697) );
AND2x2_ASAP7_75t_L g744 ( .A(n_532), .B(n_573), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_538), .Y(n_533) );
AOI222xp33_ASAP7_75t_L g732 ( .A1(n_540), .A2(n_604), .B1(n_647), .B2(n_707), .C1(n_733), .C2(n_735), .Y(n_732) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_552), .Y(n_541) );
AND2x2_ASAP7_75t_L g651 ( .A(n_542), .B(n_571), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_542), .B(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g780 ( .A(n_542), .B(n_620), .Y(n_780) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_543), .A2(n_611), .B(n_615), .Y(n_610) );
AND2x2_ASAP7_75t_L g691 ( .A(n_543), .B(n_574), .Y(n_691) );
OR2x2_ASAP7_75t_L g716 ( .A(n_543), .B(n_575), .Y(n_716) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx5_ASAP7_75t_L g570 ( .A(n_544), .Y(n_570) );
AND2x2_ASAP7_75t_L g657 ( .A(n_544), .B(n_639), .Y(n_657) );
AND2x2_ASAP7_75t_L g683 ( .A(n_544), .B(n_559), .Y(n_683) );
OR2x2_ASAP7_75t_L g686 ( .A(n_544), .B(n_573), .Y(n_686) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_544), .Y(n_704) );
AND2x4_ASAP7_75t_SL g761 ( .A(n_544), .B(n_638), .Y(n_761) );
OR2x2_ASAP7_75t_L g770 ( .A(n_544), .B(n_597), .Y(n_770) );
OR2x6_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
INVx1_ASAP7_75t_L g603 ( .A(n_552), .Y(n_603) );
AOI221xp5_ASAP7_75t_SL g721 ( .A1(n_552), .A2(n_605), .B1(n_722), .B2(n_724), .C(n_725), .Y(n_721) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_559), .Y(n_552) );
OR2x2_ASAP7_75t_L g660 ( .A(n_553), .B(n_630), .Y(n_660) );
OR2x2_ASAP7_75t_L g670 ( .A(n_553), .B(n_671), .Y(n_670) );
OR2x2_ASAP7_75t_L g696 ( .A(n_553), .B(n_697), .Y(n_696) );
AND2x4_ASAP7_75t_L g702 ( .A(n_553), .B(n_621), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_553), .B(n_685), .Y(n_714) );
INVx2_ASAP7_75t_L g727 ( .A(n_553), .Y(n_727) );
NAND2xp5_ASAP7_75t_SL g748 ( .A(n_553), .B(n_605), .Y(n_748) );
AND2x2_ASAP7_75t_L g752 ( .A(n_553), .B(n_574), .Y(n_752) );
AND2x2_ASAP7_75t_L g760 ( .A(n_553), .B(n_761), .Y(n_760) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g573 ( .A(n_554), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_559), .B(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g604 ( .A(n_559), .B(n_573), .Y(n_604) );
INVx2_ASAP7_75t_L g621 ( .A(n_559), .Y(n_621) );
AND2x4_ASAP7_75t_L g638 ( .A(n_559), .B(n_639), .Y(n_638) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_559), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_565), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_568), .B(n_571), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g750 ( .A(n_569), .B(n_572), .Y(n_750) );
AND2x4_ASAP7_75t_L g596 ( .A(n_570), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g637 ( .A(n_570), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g664 ( .A(n_570), .B(n_604), .Y(n_664) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
AND2x2_ASAP7_75t_L g768 ( .A(n_572), .B(n_769), .Y(n_768) );
BUFx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g620 ( .A(n_573), .B(n_621), .Y(n_620) );
OAI21xp5_ASAP7_75t_SL g640 ( .A1(n_574), .A2(n_641), .B(n_647), .Y(n_640) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_587), .Y(n_577) );
INVx1_ASAP7_75t_SL g694 ( .A(n_578), .Y(n_694) );
AND2x2_ASAP7_75t_L g724 ( .A(n_578), .B(n_634), .Y(n_724) );
AND2x4_ASAP7_75t_L g735 ( .A(n_578), .B(n_736), .Y(n_735) );
OR2x2_ASAP7_75t_L g601 ( .A(n_579), .B(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g608 ( .A(n_579), .Y(n_608) );
AND2x4_ASAP7_75t_L g614 ( .A(n_579), .B(n_600), .Y(n_614) );
INVx2_ASAP7_75t_L g625 ( .A(n_579), .Y(n_625) );
INVx1_ASAP7_75t_L g674 ( .A(n_579), .Y(n_674) );
OR2x2_ASAP7_75t_L g695 ( .A(n_579), .B(n_679), .Y(n_695) );
OR2x2_ASAP7_75t_L g709 ( .A(n_579), .B(n_589), .Y(n_709) );
HB1xp67_ASAP7_75t_L g775 ( .A(n_579), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_579), .B(n_631), .Y(n_781) );
OR2x6_ASAP7_75t_L g579 ( .A(n_580), .B(n_586), .Y(n_579) );
INVx1_ASAP7_75t_L g626 ( .A(n_587), .Y(n_626) );
AND2x2_ASAP7_75t_L g759 ( .A(n_587), .B(n_625), .Y(n_759) );
AND2x2_ASAP7_75t_L g784 ( .A(n_587), .B(n_614), .Y(n_784) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g602 ( .A(n_589), .Y(n_602) );
BUFx3_ASAP7_75t_L g644 ( .A(n_589), .Y(n_644) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_589), .Y(n_671) );
INVx1_ASAP7_75t_L g680 ( .A(n_589), .Y(n_680) );
AOI33xp33_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_598), .A3(n_603), .B1(n_604), .B2(n_605), .B3(n_606), .Y(n_595) );
AOI21x1_ASAP7_75t_SL g698 ( .A1(n_596), .A2(n_620), .B(n_682), .Y(n_698) );
INVx2_ASAP7_75t_L g728 ( .A(n_596), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_596), .B(n_727), .Y(n_734) );
AND2x2_ASAP7_75t_L g682 ( .A(n_597), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
AND2x2_ASAP7_75t_L g645 ( .A(n_600), .B(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g746 ( .A(n_601), .Y(n_746) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_602), .Y(n_736) );
OAI32xp33_ASAP7_75t_L g785 ( .A1(n_603), .A2(n_605), .A3(n_781), .B1(n_786), .B2(n_788), .Y(n_785) );
AND2x2_ASAP7_75t_L g703 ( .A(n_604), .B(n_704), .Y(n_703) );
INVx2_ASAP7_75t_SL g693 ( .A(n_605), .Y(n_693) );
AND2x2_ASAP7_75t_L g758 ( .A(n_605), .B(n_702), .Y(n_758) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OAI221xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_619), .B1(n_622), .B2(n_636), .C(n_640), .Y(n_609) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_613), .B(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_614), .B(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_614), .B(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_614), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g663 ( .A(n_618), .Y(n_663) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NOR3xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_627), .C(n_632), .Y(n_622) );
INVx1_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
OAI22xp33_ASAP7_75t_L g725 ( .A1(n_624), .A2(n_686), .B1(n_726), .B2(n_729), .Y(n_725) );
OR2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
INVx1_ASAP7_75t_L g629 ( .A(n_625), .Y(n_629) );
NOR2x1p5_ASAP7_75t_L g643 ( .A(n_625), .B(n_644), .Y(n_643) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_625), .Y(n_665) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OAI322xp33_ASAP7_75t_L g692 ( .A1(n_628), .A2(n_670), .A3(n_693), .B1(n_694), .B2(n_695), .C1(n_696), .C2(n_698), .Y(n_692) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
A2O1A1Ixp33_ASAP7_75t_L g648 ( .A1(n_630), .A2(n_649), .B(n_650), .C(n_652), .Y(n_648) );
OR2x2_ASAP7_75t_L g740 ( .A(n_630), .B(n_694), .Y(n_740) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g647 ( .A(n_631), .B(n_635), .Y(n_647) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g653 ( .A(n_637), .B(n_654), .Y(n_653) );
INVx3_ASAP7_75t_SL g685 ( .A(n_638), .Y(n_685) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_642), .B(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
INVx1_ASAP7_75t_SL g689 ( .A(n_645), .Y(n_689) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_646), .Y(n_731) );
OR2x6_ASAP7_75t_SL g786 ( .A(n_649), .B(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVxp67_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AOI211xp5_ASAP7_75t_L g776 ( .A1(n_654), .A2(n_777), .B(n_778), .C(n_785), .Y(n_776) );
O2A1O1Ixp33_ASAP7_75t_SL g655 ( .A1(n_656), .A2(n_658), .B(n_661), .C(n_665), .Y(n_655) );
OAI211xp5_ASAP7_75t_SL g667 ( .A1(n_656), .A2(n_668), .B(n_675), .C(n_699), .Y(n_667) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx3_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVxp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
NOR3xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_712), .C(n_756), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_672), .Y(n_668) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_671), .Y(n_763) );
INVx1_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g718 ( .A(n_674), .Y(n_718) );
NOR3xp33_ASAP7_75t_SL g675 ( .A(n_676), .B(n_688), .C(n_692), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_681), .B1(n_684), .B2(n_687), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g720 ( .A(n_680), .Y(n_720) );
INVxp67_ASAP7_75t_SL g787 ( .A(n_680), .Y(n_787) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
OR2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
INVx1_ASAP7_75t_SL g773 ( .A(n_686), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
OR2x2_ASAP7_75t_L g723 ( .A(n_689), .B(n_709), .Y(n_723) );
OR2x2_ASAP7_75t_L g774 ( .A(n_689), .B(n_775), .Y(n_774) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g772 ( .A(n_697), .Y(n_772) );
OR2x2_ASAP7_75t_L g788 ( .A(n_697), .B(n_727), .Y(n_788) );
OAI21xp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_703), .B(n_705), .Y(n_699) );
OAI31xp33_ASAP7_75t_L g713 ( .A1(n_700), .A2(n_714), .A3(n_715), .B(n_717), .Y(n_713) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_710), .Y(n_707) );
INVx1_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
AND2x4_ASAP7_75t_L g745 ( .A(n_710), .B(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
NAND4xp25_ASAP7_75t_SL g712 ( .A(n_713), .B(n_721), .C(n_732), .D(n_737), .Y(n_712) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
HB1xp67_ASAP7_75t_L g755 ( .A(n_720), .Y(n_755) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
OR2x2_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
INVxp67_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
AOI221xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_741), .B1(n_745), .B2(n_747), .C(n_749), .Y(n_737) );
NAND2xp33_ASAP7_75t_SL g738 ( .A(n_739), .B(n_740), .Y(n_738) );
INVx1_ASAP7_75t_L g782 ( .A(n_741), .Y(n_782) );
AND2x2_ASAP7_75t_SL g741 ( .A(n_742), .B(n_744), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
AOI21xp33_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_751), .B(n_753), .Y(n_749) );
INVx1_ASAP7_75t_L g777 ( .A(n_751), .Y(n_777) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
NAND2xp5_ASAP7_75t_SL g756 ( .A(n_757), .B(n_776), .Y(n_756) );
AOI221xp5_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_759), .B1(n_760), .B2(n_762), .C(n_766), .Y(n_757) );
AND2x2_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
INVx1_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
AOI21xp33_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_771), .B(n_774), .Y(n_766) );
INVxp33_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_SL g769 ( .A(n_770), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_772), .B(n_773), .Y(n_771) );
OAI22xp5_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_781), .B1(n_782), .B2(n_783), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
CKINVDCx5p33_ASAP7_75t_R g789 ( .A(n_790), .Y(n_789) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_790), .Y(n_800) );
CKINVDCx11_ASAP7_75t_R g790 ( .A(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx2_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_805), .B(n_808), .Y(n_804) );
CKINVDCx11_ASAP7_75t_R g805 ( .A(n_806), .Y(n_805) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_807), .Y(n_806) );
INVxp67_ASAP7_75t_SL g820 ( .A(n_808), .Y(n_820) );
XNOR2xp5_ASAP7_75t_L g808 ( .A(n_809), .B(n_813), .Y(n_808) );
NAND3x1_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .C(n_812), .Y(n_809) );
CKINVDCx5p33_ASAP7_75t_R g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g818 ( .A(n_816), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g821 ( .A(n_822), .B(n_823), .Y(n_821) );
CKINVDCx5p33_ASAP7_75t_R g824 ( .A(n_825), .Y(n_824) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .Y(n_826) );
endmodule