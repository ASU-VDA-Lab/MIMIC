module fake_ariane_1546_n_1236 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1236);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1236;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_423;
wire n_603;
wire n_373;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_187;
wire n_817;
wire n_924;
wire n_781;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_524;
wire n_1214;
wire n_634;
wire n_1138;
wire n_214;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_232;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1018;
wire n_259;
wire n_953;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_200;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_868;
wire n_884;
wire n_1034;
wire n_1085;
wire n_277;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_929;
wire n_206;
wire n_899;
wire n_352;
wire n_611;
wire n_365;
wire n_238;
wire n_1013;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_440;
wire n_273;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_461;
wire n_1121;
wire n_209;
wire n_490;
wire n_225;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_676;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_555;
wire n_804;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_513;
wire n_288;
wire n_1178;
wire n_1026;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_1083;
wire n_967;
wire n_746;
wire n_292;
wire n_1079;
wire n_615;
wire n_1139;
wire n_517;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_470;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_299;
wire n_836;
wire n_564;
wire n_205;
wire n_1029;
wire n_760;
wire n_522;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_598;
wire n_345;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_776;
wire n_424;
wire n_466;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_553;
wire n_814;
wire n_578;
wire n_405;
wire n_320;
wire n_1134;
wire n_647;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_218;
wire n_247;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_233;
wire n_957;
wire n_388;
wire n_1218;
wire n_321;
wire n_221;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_845;
wire n_888;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_769;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_999;
wire n_456;
wire n_852;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_317;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_687;
wire n_797;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_393;
wire n_474;
wire n_805;
wire n_295;
wire n_190;
wire n_1072;
wire n_695;
wire n_180;
wire n_730;
wire n_386;
wire n_516;
wire n_1137;
wire n_197;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_752;
wire n_985;
wire n_421;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_649;
wire n_374;
wire n_643;
wire n_226;
wire n_682;
wire n_819;
wire n_586;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_272;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_224;
wire n_894;
wire n_420;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_181;
wire n_617;
wire n_543;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_613;
wire n_1022;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_213;
wire n_1014;
wire n_724;
wire n_493;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_1183;
wire n_981;
wire n_1110;
wire n_243;
wire n_185;
wire n_1204;
wire n_994;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_828;
wire n_322;
wire n_558;
wire n_653;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1167;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_244;
wire n_679;
wire n_220;
wire n_663;
wire n_443;
wire n_528;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_385;
wire n_917;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1064;
wire n_633;
wire n_900;
wire n_1093;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_835;
wire n_446;
wire n_1076;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_188;
wire n_323;
wire n_550;
wire n_997;
wire n_635;
wire n_694;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_228;
wire n_671;
wire n_1148;
wire n_654;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_658;
wire n_630;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_196;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1229;
wire n_415;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_895;
wire n_304;
wire n_583;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_265;
wire n_208;
wire n_275;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_963;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1001;
wire n_1115;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_250;
wire n_773;
wire n_1010;
wire n_882;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_548;
wire n_289;
wire n_523;
wire n_457;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_573;
wire n_796;
wire n_531;
wire n_675;

INVx1_ASAP7_75t_L g180 ( 
.A(n_77),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_162),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_15),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_81),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_169),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_124),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_118),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_119),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_38),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_1),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_34),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_23),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_108),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_132),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_36),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_172),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_41),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_12),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_87),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_97),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_128),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_46),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_138),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_75),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_171),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_68),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_167),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_120),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_13),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_155),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_70),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_85),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_90),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_163),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_121),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_141),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_99),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_56),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_80),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_160),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_22),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_115),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_157),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_57),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_76),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_84),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_123),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_13),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_156),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_60),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_37),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_42),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_150),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_5),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_83),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_50),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_148),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_147),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_66),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_65),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_158),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_5),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_143),
.Y(n_245)
);

BUFx5_ASAP7_75t_L g246 ( 
.A(n_89),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_53),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_24),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_61),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_107),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_73),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_125),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_41),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_30),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_178),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_25),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_9),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_102),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_31),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_34),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_144),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_139),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_154),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_11),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_28),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_31),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_170),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_149),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_135),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_48),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_133),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_96),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_21),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_33),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_0),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_7),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_179),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_146),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_69),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_174),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_23),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_161),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_27),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_152),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_165),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_117),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_95),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_43),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_103),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_112),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_145),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_43),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_140),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_38),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_16),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_3),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_51),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_27),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_10),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_72),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_274),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_192),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_184),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_193),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_194),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_275),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_200),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_218),
.B(n_0),
.Y(n_308)
);

INVxp33_ASAP7_75t_SL g309 ( 
.A(n_190),
.Y(n_309)
);

NOR2xp67_ASAP7_75t_L g310 ( 
.A(n_190),
.B(n_1),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_253),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_257),
.Y(n_312)
);

NOR2xp67_ASAP7_75t_L g313 ( 
.A(n_197),
.B(n_2),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_192),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_264),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_264),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_273),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_265),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_197),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_206),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_198),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_180),
.B(n_2),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_211),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_223),
.Y(n_324)
);

INVxp33_ASAP7_75t_SL g325 ( 
.A(n_199),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_230),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_266),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_233),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_206),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_281),
.B(n_3),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_186),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_283),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_292),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_299),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_199),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_234),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_273),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_236),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_186),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_240),
.Y(n_340)
);

BUFx2_ASAP7_75t_L g341 ( 
.A(n_288),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_273),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_182),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_240),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_288),
.Y(n_345)
);

INVxp33_ASAP7_75t_L g346 ( 
.A(n_227),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_294),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_191),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_196),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_300),
.B(n_4),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_204),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_205),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_249),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_294),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_209),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_241),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_245),
.Y(n_357)
);

BUFx10_ASAP7_75t_L g358 ( 
.A(n_181),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_219),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_245),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_295),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_222),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_187),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_244),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_295),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_248),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_225),
.B(n_4),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_226),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_296),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_254),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_296),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_256),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_228),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_259),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_239),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_242),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_260),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_243),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_249),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_247),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_276),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_298),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_261),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_185),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_263),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_201),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_272),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_286),
.Y(n_388)
);

INVxp67_ASAP7_75t_SL g389 ( 
.A(n_285),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_285),
.Y(n_390)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_227),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_353),
.B(n_293),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_384),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_329),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_343),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_348),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_329),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_339),
.B(n_235),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_349),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_351),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_352),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_386),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_357),
.Y(n_403)
);

AND3x2_ASAP7_75t_L g404 ( 
.A(n_317),
.B(n_258),
.C(n_237),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_R g405 ( 
.A(n_363),
.B(n_202),
.Y(n_405)
);

BUFx8_ASAP7_75t_L g406 ( 
.A(n_335),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_361),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_355),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_359),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_362),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_379),
.B(n_181),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_368),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_357),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_373),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_375),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_376),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_331),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_378),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_361),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_363),
.B(n_187),
.Y(n_420)
);

AND2x6_ASAP7_75t_L g421 ( 
.A(n_320),
.B(n_237),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_380),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_383),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_385),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_339),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_320),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_387),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_340),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_388),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_346),
.B(n_214),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_391),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_303),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_321),
.B(n_188),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_304),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_340),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_371),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_389),
.B(n_214),
.Y(n_437)
);

INVxp67_ASAP7_75t_SL g438 ( 
.A(n_337),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_305),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_341),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_307),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_358),
.B(n_251),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_321),
.B(n_188),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_344),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_371),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_311),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_312),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_318),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_333),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_344),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_360),
.Y(n_451)
);

BUFx10_ASAP7_75t_L g452 ( 
.A(n_356),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_372),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_334),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_322),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_360),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_350),
.Y(n_457)
);

OA21x2_ASAP7_75t_L g458 ( 
.A1(n_367),
.A2(n_269),
.B(n_258),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_327),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_358),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_323),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_405),
.B(n_356),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_426),
.Y(n_463)
);

INVx4_ASAP7_75t_L g464 ( 
.A(n_427),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_426),
.B(n_358),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_397),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_397),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_426),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_460),
.B(n_324),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_394),
.Y(n_470)
);

BUFx4f_ASAP7_75t_L g471 ( 
.A(n_458),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_417),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_460),
.B(n_326),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_455),
.A2(n_308),
.B1(n_457),
.B2(n_325),
.Y(n_474)
);

NAND2xp33_ASAP7_75t_L g475 ( 
.A(n_460),
.B(n_246),
.Y(n_475)
);

OAI221xp5_ASAP7_75t_L g476 ( 
.A1(n_455),
.A2(n_330),
.B1(n_332),
.B2(n_306),
.C(n_310),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_426),
.B(n_328),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_394),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_394),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_457),
.A2(n_325),
.B1(n_309),
.B2(n_459),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_397),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_399),
.Y(n_482)
);

NOR3xp33_ASAP7_75t_L g483 ( 
.A(n_453),
.B(n_365),
.C(n_354),
.Y(n_483)
);

AND2x6_ASAP7_75t_L g484 ( 
.A(n_430),
.B(n_269),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_397),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_397),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_393),
.B(n_402),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_461),
.B(n_309),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_397),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_427),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_459),
.B(n_342),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_452),
.B(n_336),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_420),
.B(n_338),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_452),
.B(n_364),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_427),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_452),
.B(n_366),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_427),
.Y(n_497)
);

AND2x2_ASAP7_75t_SL g498 ( 
.A(n_458),
.B(n_278),
.Y(n_498)
);

NAND2xp33_ASAP7_75t_L g499 ( 
.A(n_442),
.B(n_246),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_452),
.B(n_370),
.Y(n_500)
);

NAND2xp33_ASAP7_75t_SL g501 ( 
.A(n_433),
.B(n_382),
.Y(n_501)
);

BUFx10_ASAP7_75t_L g502 ( 
.A(n_403),
.Y(n_502)
);

INVxp33_ASAP7_75t_L g503 ( 
.A(n_398),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_431),
.B(n_369),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_427),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_427),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_431),
.B(n_390),
.Y(n_507)
);

BUFx10_ASAP7_75t_L g508 ( 
.A(n_395),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_L g509 ( 
.A1(n_458),
.A2(n_390),
.B1(n_301),
.B2(n_347),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_440),
.Y(n_510)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_441),
.Y(n_511)
);

OR2x6_ASAP7_75t_L g512 ( 
.A(n_412),
.B(n_313),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_441),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_441),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_430),
.B(n_345),
.Y(n_515)
);

INVx4_ASAP7_75t_L g516 ( 
.A(n_441),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_411),
.B(n_319),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_441),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_437),
.B(n_189),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_453),
.B(n_372),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_441),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_399),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_438),
.B(n_381),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_395),
.B(n_396),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_413),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_399),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_392),
.B(n_189),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_434),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_434),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_400),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_L g531 ( 
.A1(n_458),
.A2(n_381),
.B1(n_377),
.B2(n_374),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_396),
.B(n_195),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_475),
.A2(n_465),
.B(n_477),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_480),
.A2(n_443),
.B1(n_423),
.B2(n_410),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_507),
.B(n_374),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_524),
.B(n_434),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_504),
.B(n_434),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_524),
.B(n_454),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_524),
.B(n_454),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_508),
.B(n_454),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_470),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_524),
.B(n_454),
.Y(n_542)
);

AO22x1_ASAP7_75t_L g543 ( 
.A1(n_523),
.A2(n_406),
.B1(n_451),
.B2(n_450),
.Y(n_543)
);

AND2x6_ASAP7_75t_SL g544 ( 
.A(n_493),
.B(n_302),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_510),
.B(n_401),
.Y(n_545)
);

INVxp67_ASAP7_75t_SL g546 ( 
.A(n_463),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_474),
.B(n_401),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_508),
.B(n_410),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_482),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_508),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_470),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_474),
.B(n_414),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_482),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_463),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_508),
.B(n_414),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_510),
.B(n_377),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_526),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_480),
.B(n_407),
.Y(n_558)
);

NOR3xp33_ASAP7_75t_L g559 ( 
.A(n_525),
.B(n_445),
.C(n_436),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_468),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_478),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_526),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_530),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_475),
.A2(n_423),
.B(n_415),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_528),
.B(n_415),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_528),
.B(n_424),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_530),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_484),
.A2(n_491),
.B1(n_512),
.B2(n_476),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_528),
.Y(n_569)
);

A2O1A1Ixp33_ASAP7_75t_L g570 ( 
.A1(n_471),
.A2(n_529),
.B(n_491),
.C(n_515),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_471),
.B(n_424),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_529),
.B(n_400),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_478),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_479),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_529),
.B(n_400),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_479),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_471),
.B(n_408),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_527),
.B(n_408),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_517),
.B(n_408),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_468),
.Y(n_580)
);

O2A1O1Ixp33_ASAP7_75t_L g581 ( 
.A1(n_532),
.A2(n_449),
.B(n_448),
.C(n_447),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_522),
.Y(n_582)
);

BUFx6f_ASAP7_75t_SL g583 ( 
.A(n_502),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_491),
.B(n_409),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_522),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_484),
.A2(n_416),
.B1(n_422),
.B2(n_409),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_469),
.B(n_473),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_491),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_519),
.A2(n_432),
.B1(n_449),
.B2(n_448),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_490),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_512),
.B(n_412),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_525),
.Y(n_592)
);

OAI221xp5_ASAP7_75t_L g593 ( 
.A1(n_509),
.A2(n_432),
.B1(n_447),
.B2(n_418),
.C(n_429),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_472),
.B(n_419),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_506),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_484),
.B(n_409),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_520),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_464),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_520),
.B(n_445),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_484),
.B(n_416),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_484),
.B(n_416),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_498),
.B(n_418),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_506),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_484),
.B(n_418),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_513),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_513),
.Y(n_606)
);

NOR3xp33_ASAP7_75t_L g607 ( 
.A(n_487),
.B(n_428),
.C(n_425),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_498),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_484),
.B(n_422),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_490),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_498),
.B(n_422),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_514),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_512),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_512),
.A2(n_429),
.B1(n_446),
.B2(n_439),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_514),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_488),
.B(n_456),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_492),
.B(n_435),
.Y(n_617)
);

INVx4_ASAP7_75t_L g618 ( 
.A(n_464),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_518),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_464),
.B(n_429),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_518),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_512),
.B(n_439),
.Y(n_622)
);

NAND3xp33_ASAP7_75t_L g623 ( 
.A(n_531),
.B(n_406),
.C(n_439),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_494),
.B(n_444),
.Y(n_624)
);

OR2x6_ASAP7_75t_L g625 ( 
.A(n_462),
.B(n_446),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_490),
.B(n_446),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_505),
.B(n_421),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_486),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_495),
.A2(n_421),
.B1(n_406),
.B2(n_251),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_511),
.B(n_195),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_584),
.B(n_496),
.Y(n_631)
);

O2A1O1Ixp33_ASAP7_75t_L g632 ( 
.A1(n_547),
.A2(n_500),
.B(n_499),
.C(n_483),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_538),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_538),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_541),
.Y(n_635)
);

AO21x1_ASAP7_75t_L g636 ( 
.A1(n_577),
.A2(n_516),
.B(n_511),
.Y(n_636)
);

AOI21x1_ASAP7_75t_L g637 ( 
.A1(n_602),
.A2(n_486),
.B(n_287),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_533),
.A2(n_571),
.B(n_577),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_592),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_571),
.A2(n_499),
.B(n_505),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_548),
.A2(n_521),
.B(n_505),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_541),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_548),
.A2(n_485),
.B(n_466),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_555),
.A2(n_485),
.B(n_466),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_542),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_550),
.B(n_502),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_584),
.B(n_406),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_L g648 ( 
.A1(n_602),
.A2(n_521),
.B(n_485),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_535),
.A2(n_558),
.B1(n_608),
.B2(n_568),
.Y(n_649)
);

NAND2x2_ASAP7_75t_L g650 ( 
.A(n_599),
.B(n_502),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_579),
.B(n_521),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_556),
.B(n_302),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_545),
.B(n_398),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_552),
.B(n_511),
.Y(n_654)
);

NOR2x1p5_ASAP7_75t_SL g655 ( 
.A(n_551),
.B(n_246),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_537),
.B(n_516),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_555),
.A2(n_466),
.B(n_516),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_551),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_572),
.A2(n_575),
.B(n_540),
.Y(n_659)
);

OAI21xp5_ASAP7_75t_L g660 ( 
.A1(n_611),
.A2(n_497),
.B(n_495),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_540),
.A2(n_578),
.B(n_626),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g662 ( 
.A(n_594),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_588),
.B(n_497),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_L g664 ( 
.A1(n_539),
.A2(n_481),
.B1(n_215),
.B2(n_489),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_550),
.B(n_501),
.Y(n_665)
);

OAI21xp5_ASAP7_75t_L g666 ( 
.A1(n_564),
.A2(n_481),
.B(n_421),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_542),
.B(n_467),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_616),
.B(n_599),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_620),
.A2(n_489),
.B(n_467),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_597),
.B(n_503),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_536),
.B(n_467),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_545),
.B(n_314),
.Y(n_672)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_620),
.A2(n_489),
.B(n_467),
.Y(n_673)
);

AND2x6_ASAP7_75t_L g674 ( 
.A(n_536),
.B(n_489),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_570),
.A2(n_489),
.B(n_467),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_565),
.A2(n_291),
.B(n_289),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_536),
.B(n_591),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_617),
.Y(n_678)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_591),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_591),
.B(n_404),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_534),
.B(n_613),
.Y(n_681)
);

NAND2xp33_ASAP7_75t_L g682 ( 
.A(n_598),
.B(n_421),
.Y(n_682)
);

OAI321xp33_ASAP7_75t_L g683 ( 
.A1(n_589),
.A2(n_593),
.A3(n_623),
.B1(n_624),
.B2(n_629),
.C(n_614),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_549),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_613),
.B(n_421),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_553),
.Y(n_686)
);

AOI21xp5_ASAP7_75t_L g687 ( 
.A1(n_566),
.A2(n_291),
.B(n_289),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_587),
.B(n_314),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_546),
.A2(n_207),
.B(n_203),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_598),
.A2(n_210),
.B(n_208),
.Y(n_690)
);

OAI21xp5_ASAP7_75t_L g691 ( 
.A1(n_627),
.A2(n_421),
.B(n_278),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_622),
.B(n_561),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_561),
.B(n_421),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_573),
.B(n_421),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_598),
.A2(n_255),
.B(n_297),
.Y(n_695)
);

OAI21xp5_ASAP7_75t_L g696 ( 
.A1(n_569),
.A2(n_287),
.B(n_290),
.Y(n_696)
);

OAI22xp5_ASAP7_75t_L g697 ( 
.A1(n_570),
.A2(n_608),
.B1(n_560),
.B2(n_557),
.Y(n_697)
);

NAND3xp33_ASAP7_75t_L g698 ( 
.A(n_559),
.B(n_316),
.C(n_315),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_573),
.B(n_212),
.Y(n_699)
);

OAI21xp5_ASAP7_75t_L g700 ( 
.A1(n_574),
.A2(n_576),
.B(n_563),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_581),
.A2(n_290),
.B(n_213),
.Y(n_701)
);

O2A1O1Ixp33_ASAP7_75t_SL g702 ( 
.A1(n_630),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_562),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_560),
.B(n_216),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_590),
.A2(n_252),
.B(n_284),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_543),
.Y(n_706)
);

O2A1O1Ixp5_ASAP7_75t_L g707 ( 
.A1(n_630),
.A2(n_6),
.B(n_8),
.C(n_9),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_567),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_574),
.B(n_217),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_554),
.Y(n_710)
);

INVx1_ASAP7_75t_SL g711 ( 
.A(n_625),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_576),
.A2(n_250),
.B(n_220),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_618),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_610),
.A2(n_262),
.B(n_221),
.Y(n_714)
);

OAI22xp5_ASAP7_75t_L g715 ( 
.A1(n_554),
.A2(n_316),
.B1(n_315),
.B2(n_282),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_628),
.A2(n_605),
.B(n_621),
.Y(n_716)
);

AND2x2_ASAP7_75t_SL g717 ( 
.A(n_607),
.B(n_183),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_582),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_625),
.B(n_618),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_585),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_625),
.B(n_224),
.Y(n_721)
);

NOR2x1_ASAP7_75t_L g722 ( 
.A(n_625),
.B(n_183),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_595),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_595),
.Y(n_724)
);

NOR3xp33_ASAP7_75t_L g725 ( 
.A(n_618),
.B(n_580),
.C(n_554),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_580),
.B(n_231),
.Y(n_726)
);

OAI21x1_ASAP7_75t_L g727 ( 
.A1(n_638),
.A2(n_628),
.B(n_596),
.Y(n_727)
);

AOI21x1_ASAP7_75t_SL g728 ( 
.A1(n_656),
.A2(n_600),
.B(n_601),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_684),
.Y(n_729)
);

AO21x1_ASAP7_75t_L g730 ( 
.A1(n_697),
.A2(n_604),
.B(n_609),
.Y(n_730)
);

OAI21x1_ASAP7_75t_L g731 ( 
.A1(n_638),
.A2(n_621),
.B(n_619),
.Y(n_731)
);

A2O1A1Ixp33_ASAP7_75t_L g732 ( 
.A1(n_649),
.A2(n_586),
.B(n_580),
.C(n_612),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_661),
.A2(n_619),
.B(n_615),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_674),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_659),
.A2(n_615),
.B(n_612),
.Y(n_735)
);

OAI21x1_ASAP7_75t_L g736 ( 
.A1(n_675),
.A2(n_637),
.B(n_659),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_678),
.Y(n_737)
);

OAI21x1_ASAP7_75t_L g738 ( 
.A1(n_675),
.A2(n_606),
.B(n_605),
.Y(n_738)
);

OAI21x1_ASAP7_75t_L g739 ( 
.A1(n_669),
.A2(n_606),
.B(n_603),
.Y(n_739)
);

NAND3xp33_ASAP7_75t_L g740 ( 
.A(n_662),
.B(n_603),
.C(n_270),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_635),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_674),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_674),
.Y(n_743)
);

AO21x1_ASAP7_75t_L g744 ( 
.A1(n_701),
.A2(n_246),
.B(n_229),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_651),
.A2(n_268),
.B(n_280),
.Y(n_745)
);

BUFx2_ASAP7_75t_L g746 ( 
.A(n_639),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_668),
.B(n_544),
.Y(n_747)
);

OAI21x1_ASAP7_75t_L g748 ( 
.A1(n_669),
.A2(n_246),
.B(n_583),
.Y(n_748)
);

AND3x2_ASAP7_75t_L g749 ( 
.A(n_652),
.B(n_583),
.C(n_11),
.Y(n_749)
);

AO21x1_ASAP7_75t_L g750 ( 
.A1(n_701),
.A2(n_246),
.B(n_229),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_688),
.A2(n_583),
.B1(n_279),
.B2(n_277),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_653),
.A2(n_271),
.B1(n_267),
.B2(n_238),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_633),
.B(n_10),
.Y(n_753)
);

OAI21x1_ASAP7_75t_L g754 ( 
.A1(n_673),
.A2(n_246),
.B(n_229),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_647),
.B(n_12),
.Y(n_755)
);

OAI21x1_ASAP7_75t_L g756 ( 
.A1(n_673),
.A2(n_183),
.B(n_229),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_634),
.B(n_14),
.Y(n_757)
);

OAI21x1_ASAP7_75t_L g758 ( 
.A1(n_716),
.A2(n_92),
.B(n_129),
.Y(n_758)
);

OAI22x1_ASAP7_75t_L g759 ( 
.A1(n_698),
.A2(n_232),
.B1(n_15),
.B2(n_16),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_686),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_703),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_708),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_642),
.Y(n_763)
);

OAI21x1_ASAP7_75t_L g764 ( 
.A1(n_716),
.A2(n_183),
.B(n_93),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_682),
.A2(n_91),
.B(n_177),
.Y(n_765)
);

A2O1A1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_632),
.A2(n_14),
.B(n_17),
.C(n_18),
.Y(n_766)
);

OAI21x1_ASAP7_75t_L g767 ( 
.A1(n_640),
.A2(n_722),
.B(n_666),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_717),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_631),
.B(n_19),
.Y(n_769)
);

OAI21xp5_ASAP7_75t_L g770 ( 
.A1(n_654),
.A2(n_20),
.B(n_21),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_718),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_640),
.A2(n_98),
.B(n_176),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_700),
.A2(n_94),
.B(n_175),
.Y(n_773)
);

OAI21xp5_ASAP7_75t_L g774 ( 
.A1(n_648),
.A2(n_20),
.B(n_22),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_643),
.A2(n_100),
.B(n_173),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_720),
.Y(n_776)
);

OAI21x1_ASAP7_75t_SL g777 ( 
.A1(n_636),
.A2(n_24),
.B(n_25),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_658),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_667),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_674),
.Y(n_780)
);

NOR2x1_ASAP7_75t_R g781 ( 
.A(n_672),
.B(n_26),
.Y(n_781)
);

AOI21x1_ASAP7_75t_SL g782 ( 
.A1(n_671),
.A2(n_29),
.B(n_30),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_645),
.B(n_32),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_674),
.Y(n_784)
);

OAI21x1_ASAP7_75t_L g785 ( 
.A1(n_660),
.A2(n_105),
.B(n_168),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_723),
.Y(n_786)
);

OAI21x1_ASAP7_75t_L g787 ( 
.A1(n_691),
.A2(n_104),
.B(n_166),
.Y(n_787)
);

OR2x6_ASAP7_75t_L g788 ( 
.A(n_677),
.B(n_32),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_679),
.B(n_33),
.Y(n_789)
);

OAI21x1_ASAP7_75t_L g790 ( 
.A1(n_641),
.A2(n_106),
.B(n_164),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_644),
.A2(n_101),
.B(n_159),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_741),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_769),
.B(n_706),
.Y(n_793)
);

OAI21xp33_ASAP7_75t_SL g794 ( 
.A1(n_768),
.A2(n_665),
.B(n_681),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_741),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_769),
.B(n_715),
.Y(n_796)
);

OA21x2_ASAP7_75t_L g797 ( 
.A1(n_736),
.A2(n_696),
.B(n_641),
.Y(n_797)
);

O2A1O1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_766),
.A2(n_702),
.B(n_646),
.C(n_683),
.Y(n_798)
);

AND2x4_ASAP7_75t_L g799 ( 
.A(n_734),
.B(n_719),
.Y(n_799)
);

NAND2x1p5_ASAP7_75t_L g800 ( 
.A(n_734),
.B(n_719),
.Y(n_800)
);

INVx4_ASAP7_75t_L g801 ( 
.A(n_743),
.Y(n_801)
);

CKINVDCx8_ASAP7_75t_R g802 ( 
.A(n_737),
.Y(n_802)
);

OAI33xp33_ASAP7_75t_L g803 ( 
.A1(n_779),
.A2(n_670),
.A3(n_721),
.B1(n_680),
.B2(n_704),
.B3(n_709),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_755),
.B(n_711),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_755),
.B(n_747),
.Y(n_805)
);

AOI21xp33_ASAP7_75t_SL g806 ( 
.A1(n_737),
.A2(n_726),
.B(n_650),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_729),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_763),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_760),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_743),
.Y(n_810)
);

OR2x6_ASAP7_75t_L g811 ( 
.A(n_780),
.B(n_692),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_746),
.B(n_699),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_768),
.A2(n_664),
.B1(n_713),
.B2(n_663),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_759),
.A2(n_724),
.B1(n_712),
.B2(n_714),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_774),
.B(n_710),
.Y(n_815)
);

OR2x2_ASAP7_75t_L g816 ( 
.A(n_761),
.B(n_710),
.Y(n_816)
);

BUFx2_ASAP7_75t_L g817 ( 
.A(n_780),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_762),
.B(n_710),
.Y(n_818)
);

NAND2x1p5_ASAP7_75t_L g819 ( 
.A(n_742),
.B(n_713),
.Y(n_819)
);

INVx5_ASAP7_75t_L g820 ( 
.A(n_742),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_751),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_771),
.Y(n_822)
);

BUFx2_ASAP7_75t_L g823 ( 
.A(n_788),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_776),
.B(n_712),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_786),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_763),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_752),
.B(n_689),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_788),
.B(n_35),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_L g829 ( 
.A1(n_788),
.A2(n_714),
.B1(n_687),
.B2(n_676),
.Y(n_829)
);

INVxp67_ASAP7_75t_SL g830 ( 
.A(n_784),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_735),
.A2(n_657),
.B(n_725),
.Y(n_831)
);

AO21x2_ASAP7_75t_L g832 ( 
.A1(n_744),
.A2(n_693),
.B(n_694),
.Y(n_832)
);

A2O1A1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_766),
.A2(n_707),
.B(n_657),
.C(n_655),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_778),
.Y(n_834)
);

INVx8_ASAP7_75t_L g835 ( 
.A(n_784),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_778),
.B(n_685),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_738),
.Y(n_837)
);

O2A1O1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_770),
.A2(n_705),
.B(n_695),
.C(n_690),
.Y(n_838)
);

CKINVDCx6p67_ASAP7_75t_R g839 ( 
.A(n_789),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_767),
.Y(n_840)
);

INVxp67_ASAP7_75t_L g841 ( 
.A(n_781),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_738),
.Y(n_842)
);

OAI21xp5_ASAP7_75t_L g843 ( 
.A1(n_732),
.A2(n_35),
.B(n_36),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_753),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_757),
.B(n_39),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_749),
.B(n_40),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_821),
.A2(n_783),
.B1(n_740),
.B2(n_730),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_799),
.B(n_748),
.Y(n_848)
);

BUFx4f_ASAP7_75t_L g849 ( 
.A(n_800),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_817),
.Y(n_850)
);

AO21x1_ASAP7_75t_L g851 ( 
.A1(n_843),
.A2(n_773),
.B(n_785),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_792),
.Y(n_852)
);

AO21x1_ASAP7_75t_L g853 ( 
.A1(n_815),
.A2(n_785),
.B(n_733),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_807),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_799),
.B(n_748),
.Y(n_855)
);

OAI22xp33_ASAP7_75t_L g856 ( 
.A1(n_796),
.A2(n_765),
.B1(n_772),
.B2(n_791),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_812),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_809),
.Y(n_858)
);

OAI21x1_ASAP7_75t_L g859 ( 
.A1(n_831),
.A2(n_756),
.B(n_736),
.Y(n_859)
);

INVx3_ASAP7_75t_L g860 ( 
.A(n_835),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_816),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_822),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_825),
.Y(n_863)
);

OAI21x1_ASAP7_75t_L g864 ( 
.A1(n_837),
.A2(n_756),
.B(n_754),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_824),
.B(n_732),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_792),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_834),
.Y(n_867)
);

OAI21x1_ASAP7_75t_L g868 ( 
.A1(n_837),
.A2(n_754),
.B(n_764),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_SL g869 ( 
.A1(n_821),
.A2(n_793),
.B1(n_828),
.B2(n_794),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_795),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_795),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_805),
.B(n_804),
.Y(n_872)
);

NAND2x1p5_ASAP7_75t_L g873 ( 
.A(n_820),
.B(n_767),
.Y(n_873)
);

CKINVDCx11_ASAP7_75t_R g874 ( 
.A(n_802),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_835),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_808),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_808),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_823),
.B(n_811),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_826),
.Y(n_879)
);

HB1xp67_ASAP7_75t_SL g880 ( 
.A(n_802),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_803),
.A2(n_750),
.B1(n_777),
.B2(n_745),
.Y(n_881)
);

CKINVDCx6p67_ASAP7_75t_R g882 ( 
.A(n_839),
.Y(n_882)
);

OAI22xp33_ASAP7_75t_L g883 ( 
.A1(n_844),
.A2(n_775),
.B1(n_782),
.B2(n_728),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_810),
.B(n_826),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_SL g885 ( 
.A1(n_846),
.A2(n_787),
.B1(n_790),
.B2(n_764),
.Y(n_885)
);

AO21x2_ASAP7_75t_L g886 ( 
.A1(n_815),
.A2(n_739),
.B(n_731),
.Y(n_886)
);

OAI21x1_ASAP7_75t_L g887 ( 
.A1(n_840),
.A2(n_739),
.B(n_731),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_818),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_841),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_811),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_810),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_835),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_836),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_811),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_799),
.B(n_790),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_839),
.A2(n_787),
.B1(n_727),
.B2(n_758),
.Y(n_896)
);

CKINVDCx20_ASAP7_75t_R g897 ( 
.A(n_801),
.Y(n_897)
);

OAI22xp33_ASAP7_75t_L g898 ( 
.A1(n_845),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_898)
);

INVx4_ASAP7_75t_SL g899 ( 
.A(n_811),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_835),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_814),
.A2(n_727),
.B1(n_45),
.B2(n_44),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_L g902 ( 
.A1(n_814),
.A2(n_47),
.B1(n_49),
.B2(n_52),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_842),
.Y(n_903)
);

BUFx2_ASAP7_75t_L g904 ( 
.A(n_840),
.Y(n_904)
);

OR2x6_ASAP7_75t_L g905 ( 
.A(n_895),
.B(n_801),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_887),
.Y(n_906)
);

OAI21x1_ASAP7_75t_L g907 ( 
.A1(n_859),
.A2(n_840),
.B(n_797),
.Y(n_907)
);

HB1xp67_ASAP7_75t_L g908 ( 
.A(n_903),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_867),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_903),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_887),
.Y(n_911)
);

BUFx12f_ASAP7_75t_L g912 ( 
.A(n_874),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_870),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_871),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_865),
.B(n_798),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_886),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_865),
.B(n_842),
.Y(n_917)
);

OA21x2_ASAP7_75t_L g918 ( 
.A1(n_859),
.A2(n_868),
.B(n_864),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_876),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_886),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_886),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_879),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_852),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_852),
.Y(n_924)
);

NAND2x1p5_ASAP7_75t_L g925 ( 
.A(n_895),
.B(n_797),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_904),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_866),
.Y(n_927)
);

BUFx12f_ASAP7_75t_L g928 ( 
.A(n_874),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_872),
.B(n_810),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_897),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_904),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_877),
.Y(n_932)
);

OR2x6_ASAP7_75t_L g933 ( 
.A(n_895),
.B(n_848),
.Y(n_933)
);

AND2x4_ASAP7_75t_SL g934 ( 
.A(n_848),
.B(n_801),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_897),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_848),
.B(n_820),
.Y(n_936)
);

BUFx4f_ASAP7_75t_SL g937 ( 
.A(n_882),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_873),
.Y(n_938)
);

AO21x2_ASAP7_75t_L g939 ( 
.A1(n_851),
.A2(n_833),
.B(n_832),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_864),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_917),
.B(n_854),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_927),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_938),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_925),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_909),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_916),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_909),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_913),
.Y(n_948)
);

AOI22xp33_ASAP7_75t_L g949 ( 
.A1(n_915),
.A2(n_869),
.B1(n_847),
.B2(n_898),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_933),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_925),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_913),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_912),
.Y(n_953)
);

OR2x2_ASAP7_75t_L g954 ( 
.A(n_917),
.B(n_858),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_917),
.B(n_862),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_915),
.B(n_863),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_916),
.Y(n_957)
);

NOR2x1_ASAP7_75t_L g958 ( 
.A(n_929),
.B(n_878),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_927),
.Y(n_959)
);

AOI21xp33_ASAP7_75t_L g960 ( 
.A1(n_939),
.A2(n_883),
.B(n_902),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_926),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_926),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_914),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_912),
.A2(n_857),
.B1(n_851),
.B2(n_827),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_908),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_914),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_927),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_929),
.B(n_850),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_933),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_933),
.B(n_868),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_933),
.B(n_855),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_919),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_919),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_927),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_908),
.B(n_850),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_916),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_916),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_922),
.Y(n_978)
);

OR2x2_ASAP7_75t_L g979 ( 
.A(n_933),
.B(n_910),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_933),
.B(n_855),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_949),
.A2(n_882),
.B1(n_930),
.B2(n_935),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_956),
.B(n_930),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_971),
.B(n_930),
.Y(n_983)
);

NAND4xp25_ASAP7_75t_L g984 ( 
.A(n_949),
.B(n_935),
.C(n_930),
.D(n_806),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_971),
.B(n_935),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_958),
.B(n_935),
.Y(n_986)
);

NAND3xp33_ASAP7_75t_L g987 ( 
.A(n_964),
.B(n_910),
.C(n_881),
.Y(n_987)
);

NOR3xp33_ASAP7_75t_L g988 ( 
.A(n_960),
.B(n_856),
.C(n_829),
.Y(n_988)
);

AND2x2_ASAP7_75t_SL g989 ( 
.A(n_950),
.B(n_934),
.Y(n_989)
);

NAND4xp25_ASAP7_75t_L g990 ( 
.A(n_964),
.B(n_901),
.C(n_911),
.D(n_906),
.Y(n_990)
);

NAND3xp33_ASAP7_75t_L g991 ( 
.A(n_960),
.B(n_931),
.C(n_885),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_971),
.B(n_933),
.Y(n_992)
);

AND2x2_ASAP7_75t_SL g993 ( 
.A(n_950),
.B(n_934),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_SL g994 ( 
.A1(n_950),
.A2(n_934),
.B(n_925),
.Y(n_994)
);

NAND4xp25_ASAP7_75t_L g995 ( 
.A(n_968),
.B(n_956),
.C(n_975),
.D(n_955),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_980),
.B(n_905),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_980),
.B(n_905),
.Y(n_997)
);

NAND4xp25_ASAP7_75t_L g998 ( 
.A(n_968),
.B(n_975),
.C(n_955),
.D(n_941),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_SL g999 ( 
.A1(n_980),
.A2(n_934),
.B(n_925),
.Y(n_999)
);

NAND3xp33_ASAP7_75t_L g1000 ( 
.A(n_958),
.B(n_931),
.C(n_921),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_SL g1001 ( 
.A1(n_969),
.A2(n_939),
.B1(n_928),
.B2(n_912),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_954),
.A2(n_905),
.B1(n_880),
.B2(n_937),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_941),
.B(n_931),
.Y(n_1003)
);

OAI221xp5_ASAP7_75t_SL g1004 ( 
.A1(n_954),
.A2(n_979),
.B1(n_970),
.B2(n_905),
.C(n_969),
.Y(n_1004)
);

OA21x2_ASAP7_75t_L g1005 ( 
.A1(n_946),
.A2(n_920),
.B(n_921),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_995),
.B(n_965),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_996),
.B(n_970),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_998),
.B(n_965),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_1003),
.B(n_961),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_984),
.B(n_953),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_997),
.B(n_970),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_1005),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_982),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_1005),
.Y(n_1014)
);

AND2x2_ASAP7_75t_SL g1015 ( 
.A(n_989),
.B(n_979),
.Y(n_1015)
);

HB1xp67_ASAP7_75t_L g1016 ( 
.A(n_986),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_992),
.B(n_969),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_989),
.Y(n_1018)
);

INVx4_ASAP7_75t_L g1019 ( 
.A(n_993),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_993),
.B(n_969),
.Y(n_1020)
);

INVx2_ASAP7_75t_SL g1021 ( 
.A(n_986),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_1000),
.B(n_961),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_983),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_985),
.B(n_944),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_987),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_991),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_1026),
.B(n_945),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1006),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_1026),
.B(n_962),
.Y(n_1029)
);

OR2x2_ASAP7_75t_L g1030 ( 
.A(n_1009),
.B(n_1008),
.Y(n_1030)
);

OR2x6_ASAP7_75t_L g1031 ( 
.A(n_1019),
.B(n_912),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1006),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_1019),
.B(n_999),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_1019),
.B(n_994),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_1019),
.B(n_1001),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_1008),
.B(n_945),
.Y(n_1036)
);

NAND2xp33_ASAP7_75t_L g1037 ( 
.A(n_1021),
.B(n_1002),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_1027),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_1033),
.B(n_1016),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1027),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_1034),
.B(n_1031),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_L g1042 ( 
.A(n_1029),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_1031),
.B(n_1016),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_1031),
.B(n_1018),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1038),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1040),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_1042),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_1041),
.B(n_1028),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_1048),
.A2(n_1025),
.B1(n_1032),
.B2(n_1035),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_1047),
.B(n_1039),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_1048),
.B(n_1039),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_1045),
.A2(n_1025),
.B(n_1030),
.C(n_1010),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_1045),
.B(n_1040),
.Y(n_1053)
);

OAI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_1046),
.A2(n_1018),
.B1(n_1036),
.B2(n_1021),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1047),
.Y(n_1055)
);

OR2x2_ASAP7_75t_L g1056 ( 
.A(n_1047),
.B(n_1036),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1047),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1047),
.Y(n_1058)
);

INVxp67_ASAP7_75t_SL g1059 ( 
.A(n_1047),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_1059),
.B(n_1041),
.Y(n_1060)
);

INVx1_ASAP7_75t_SL g1061 ( 
.A(n_1050),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_1051),
.B(n_1043),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_1055),
.B(n_1043),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_1057),
.B(n_1044),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_1052),
.A2(n_1021),
.B1(n_981),
.B2(n_1044),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_1058),
.Y(n_1066)
);

OR2x2_ASAP7_75t_L g1067 ( 
.A(n_1056),
.B(n_1053),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1049),
.B(n_1013),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_1054),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_SL g1070 ( 
.A(n_1059),
.B(n_928),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1059),
.Y(n_1071)
);

INVx2_ASAP7_75t_SL g1072 ( 
.A(n_1055),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_1049),
.A2(n_1044),
.B1(n_1037),
.B2(n_1001),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1059),
.B(n_1013),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1059),
.Y(n_1075)
);

AOI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_1069),
.A2(n_988),
.B1(n_1018),
.B2(n_889),
.Y(n_1076)
);

AOI221xp5_ASAP7_75t_L g1077 ( 
.A1(n_1065),
.A2(n_1022),
.B1(n_990),
.B2(n_1014),
.C(n_1012),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_1062),
.B(n_1023),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_1070),
.B(n_928),
.Y(n_1079)
);

AOI322xp5_ASAP7_75t_L g1080 ( 
.A1(n_1061),
.A2(n_1012),
.A3(n_1014),
.B1(n_1022),
.B2(n_1015),
.C1(n_988),
.C2(n_928),
.Y(n_1080)
);

NOR3xp33_ASAP7_75t_L g1081 ( 
.A(n_1071),
.B(n_1004),
.C(n_1020),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_1065),
.A2(n_889),
.B(n_1009),
.Y(n_1082)
);

NAND3xp33_ASAP7_75t_L g1083 ( 
.A(n_1075),
.B(n_1004),
.C(n_1015),
.Y(n_1083)
);

OAI211xp5_ASAP7_75t_L g1084 ( 
.A1(n_1060),
.A2(n_937),
.B(n_1023),
.C(n_962),
.Y(n_1084)
);

OAI221xp5_ASAP7_75t_L g1085 ( 
.A1(n_1073),
.A2(n_1014),
.B1(n_1012),
.B2(n_1020),
.C(n_1007),
.Y(n_1085)
);

AOI222xp33_ASAP7_75t_L g1086 ( 
.A1(n_1068),
.A2(n_1015),
.B1(n_1020),
.B2(n_888),
.C1(n_1007),
.C2(n_1011),
.Y(n_1086)
);

OAI221xp5_ASAP7_75t_L g1087 ( 
.A1(n_1068),
.A2(n_1007),
.B1(n_1011),
.B2(n_1023),
.C(n_1017),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_SL g1088 ( 
.A1(n_1072),
.A2(n_838),
.B(n_1011),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1074),
.Y(n_1089)
);

AOI221xp5_ASAP7_75t_L g1090 ( 
.A1(n_1066),
.A2(n_939),
.B1(n_963),
.B2(n_972),
.C(n_948),
.Y(n_1090)
);

O2A1O1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_1067),
.A2(n_833),
.B(n_939),
.C(n_1023),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1064),
.A2(n_1024),
.B(n_1017),
.Y(n_1092)
);

AOI21xp33_ASAP7_75t_SL g1093 ( 
.A1(n_1063),
.A2(n_1024),
.B(n_1017),
.Y(n_1093)
);

AOI21x1_ASAP7_75t_L g1094 ( 
.A1(n_1074),
.A2(n_1024),
.B(n_947),
.Y(n_1094)
);

OAI22x1_ASAP7_75t_L g1095 ( 
.A1(n_1076),
.A2(n_860),
.B1(n_892),
.B2(n_900),
.Y(n_1095)
);

NOR3xp33_ASAP7_75t_L g1096 ( 
.A(n_1079),
.B(n_948),
.C(n_978),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_1078),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1088),
.A2(n_954),
.B(n_947),
.Y(n_1098)
);

AOI211x1_ASAP7_75t_L g1099 ( 
.A1(n_1082),
.A2(n_978),
.B(n_973),
.C(n_972),
.Y(n_1099)
);

INVx2_ASAP7_75t_SL g1100 ( 
.A(n_1089),
.Y(n_1100)
);

INVxp67_ASAP7_75t_L g1101 ( 
.A(n_1085),
.Y(n_1101)
);

OA22x2_ASAP7_75t_L g1102 ( 
.A1(n_1084),
.A2(n_905),
.B1(n_963),
.B2(n_973),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1094),
.Y(n_1103)
);

NAND3xp33_ASAP7_75t_L g1104 ( 
.A(n_1077),
.B(n_966),
.C(n_952),
.Y(n_1104)
);

NOR4xp75_ASAP7_75t_L g1105 ( 
.A(n_1092),
.B(n_951),
.C(n_944),
.D(n_892),
.Y(n_1105)
);

NAND3xp33_ASAP7_75t_L g1106 ( 
.A(n_1080),
.B(n_966),
.C(n_952),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_SL g1107 ( 
.A1(n_1093),
.A2(n_853),
.B(n_891),
.Y(n_1107)
);

NOR2x1_ASAP7_75t_L g1108 ( 
.A(n_1083),
.B(n_860),
.Y(n_1108)
);

NAND4xp75_ASAP7_75t_L g1109 ( 
.A(n_1090),
.B(n_813),
.C(n_853),
.D(n_891),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1086),
.B(n_944),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_1087),
.B(n_944),
.Y(n_1111)
);

OAI221xp5_ASAP7_75t_L g1112 ( 
.A1(n_1101),
.A2(n_1081),
.B1(n_1091),
.B2(n_896),
.C(n_951),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_1097),
.Y(n_1113)
);

NAND3xp33_ASAP7_75t_SL g1114 ( 
.A(n_1105),
.B(n_800),
.C(n_819),
.Y(n_1114)
);

NOR3xp33_ASAP7_75t_L g1115 ( 
.A(n_1100),
.B(n_944),
.C(n_951),
.Y(n_1115)
);

AOI211xp5_ASAP7_75t_SL g1116 ( 
.A1(n_1097),
.A2(n_892),
.B(n_900),
.C(n_860),
.Y(n_1116)
);

OAI221xp5_ASAP7_75t_L g1117 ( 
.A1(n_1098),
.A2(n_1108),
.B1(n_1103),
.B2(n_1104),
.C(n_1106),
.Y(n_1117)
);

NOR2x1_ASAP7_75t_L g1118 ( 
.A(n_1109),
.B(n_900),
.Y(n_1118)
);

AOI211xp5_ASAP7_75t_L g1119 ( 
.A1(n_1096),
.A2(n_951),
.B(n_875),
.C(n_943),
.Y(n_1119)
);

NAND3xp33_ASAP7_75t_SL g1120 ( 
.A(n_1110),
.B(n_819),
.C(n_878),
.Y(n_1120)
);

NAND4xp75_ASAP7_75t_L g1121 ( 
.A(n_1099),
.B(n_797),
.C(n_918),
.D(n_922),
.Y(n_1121)
);

NAND3xp33_ASAP7_75t_L g1122 ( 
.A(n_1111),
.B(n_943),
.C(n_820),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1095),
.A2(n_939),
.B(n_905),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_1102),
.Y(n_1124)
);

NOR3xp33_ASAP7_75t_L g1125 ( 
.A(n_1107),
.B(n_951),
.C(n_861),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1100),
.Y(n_1126)
);

OAI21xp33_ASAP7_75t_L g1127 ( 
.A1(n_1108),
.A2(n_925),
.B(n_905),
.Y(n_1127)
);

AOI221xp5_ASAP7_75t_L g1128 ( 
.A1(n_1101),
.A2(n_921),
.B1(n_920),
.B2(n_943),
.C(n_957),
.Y(n_1128)
);

NOR4xp25_ASAP7_75t_L g1129 ( 
.A(n_1100),
.B(n_911),
.C(n_906),
.D(n_920),
.Y(n_1129)
);

NAND4xp25_ASAP7_75t_SL g1130 ( 
.A(n_1098),
.B(n_979),
.C(n_911),
.D(n_906),
.Y(n_1130)
);

NOR3xp33_ASAP7_75t_L g1131 ( 
.A(n_1100),
.B(n_920),
.C(n_921),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_1097),
.B(n_875),
.Y(n_1132)
);

NOR4xp25_ASAP7_75t_L g1133 ( 
.A(n_1100),
.B(n_906),
.C(n_911),
.D(n_940),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1100),
.Y(n_1134)
);

NOR5xp2_ASAP7_75t_L g1135 ( 
.A(n_1101),
.B(n_830),
.C(n_890),
.D(n_894),
.E(n_893),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1113),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1126),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1124),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1134),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1117),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1132),
.B(n_943),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1112),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1121),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_1118),
.B(n_875),
.Y(n_1144)
);

NOR2x1_ASAP7_75t_L g1145 ( 
.A(n_1122),
.B(n_875),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1120),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1133),
.B(n_943),
.Y(n_1147)
);

AOI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_1127),
.A2(n_943),
.B1(n_875),
.B2(n_936),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1131),
.Y(n_1149)
);

AOI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1125),
.A2(n_943),
.B1(n_936),
.B2(n_836),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1135),
.Y(n_1151)
);

OR2x2_ASAP7_75t_L g1152 ( 
.A(n_1115),
.B(n_1129),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1114),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1128),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1116),
.B(n_943),
.Y(n_1155)
);

INVxp67_ASAP7_75t_L g1156 ( 
.A(n_1130),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_1119),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1123),
.B(n_940),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1113),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_1136),
.Y(n_1160)
);

OR2x2_ASAP7_75t_L g1161 ( 
.A(n_1159),
.B(n_918),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1138),
.A2(n_849),
.B(n_918),
.Y(n_1162)
);

OAI21xp33_ASAP7_75t_L g1163 ( 
.A1(n_1140),
.A2(n_936),
.B(n_940),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1152),
.Y(n_1164)
);

INVx2_ASAP7_75t_SL g1165 ( 
.A(n_1137),
.Y(n_1165)
);

NAND3xp33_ASAP7_75t_L g1166 ( 
.A(n_1139),
.B(n_820),
.C(n_938),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1151),
.B(n_946),
.Y(n_1167)
);

AOI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1143),
.A2(n_936),
.B1(n_849),
.B2(n_855),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1153),
.B(n_54),
.Y(n_1169)
);

AOI22xp5_ASAP7_75t_SL g1170 ( 
.A1(n_1157),
.A2(n_936),
.B1(n_918),
.B2(n_938),
.Y(n_1170)
);

AOI221xp5_ASAP7_75t_L g1171 ( 
.A1(n_1156),
.A2(n_836),
.B1(n_976),
.B2(n_977),
.C(n_946),
.Y(n_1171)
);

AOI221xp5_ASAP7_75t_L g1172 ( 
.A1(n_1154),
.A2(n_977),
.B1(n_976),
.B2(n_946),
.C(n_957),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1142),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1146),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1155),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_1144),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_1149),
.Y(n_1177)
);

OAI21xp33_ASAP7_75t_L g1178 ( 
.A1(n_1145),
.A2(n_936),
.B(n_940),
.Y(n_1178)
);

NAND4xp75_ASAP7_75t_L g1179 ( 
.A(n_1150),
.B(n_918),
.C(n_884),
.D(n_957),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1150),
.B(n_977),
.Y(n_1180)
);

NOR2x1_ASAP7_75t_L g1181 ( 
.A(n_1147),
.B(n_918),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1160),
.Y(n_1182)
);

AO22x2_ASAP7_75t_L g1183 ( 
.A1(n_1164),
.A2(n_1141),
.B1(n_1158),
.B2(n_1148),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1165),
.Y(n_1184)
);

NAND2xp33_ASAP7_75t_L g1185 ( 
.A(n_1176),
.B(n_1148),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1173),
.Y(n_1186)
);

INVxp67_ASAP7_75t_SL g1187 ( 
.A(n_1176),
.Y(n_1187)
);

OR2x2_ASAP7_75t_L g1188 ( 
.A(n_1174),
.B(n_907),
.Y(n_1188)
);

NAND3xp33_ASAP7_75t_SL g1189 ( 
.A(n_1177),
.B(n_1169),
.C(n_1175),
.Y(n_1189)
);

AOI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1167),
.A2(n_1168),
.B1(n_1163),
.B2(n_1162),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1176),
.B(n_907),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1161),
.B(n_907),
.Y(n_1192)
);

OR2x2_ASAP7_75t_L g1193 ( 
.A(n_1178),
.B(n_977),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1179),
.Y(n_1194)
);

OA22x2_ASAP7_75t_L g1195 ( 
.A1(n_1180),
.A2(n_1166),
.B1(n_1171),
.B2(n_1170),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1181),
.B(n_1172),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1187),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1184),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1189),
.B(n_55),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1182),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1186),
.Y(n_1201)
);

XOR2x1_ASAP7_75t_L g1202 ( 
.A(n_1194),
.B(n_58),
.Y(n_1202)
);

AOI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1183),
.A2(n_849),
.B1(n_938),
.B2(n_976),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1183),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1185),
.Y(n_1205)
);

AO22x2_ASAP7_75t_L g1206 ( 
.A1(n_1188),
.A2(n_957),
.B1(n_976),
.B2(n_899),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1196),
.B(n_59),
.Y(n_1207)
);

AO22x2_ASAP7_75t_L g1208 ( 
.A1(n_1191),
.A2(n_899),
.B1(n_967),
.B2(n_959),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1195),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1190),
.Y(n_1210)
);

XNOR2xp5_ASAP7_75t_L g1211 ( 
.A(n_1193),
.B(n_62),
.Y(n_1211)
);

OR3x1_ASAP7_75t_L g1212 ( 
.A(n_1197),
.B(n_1192),
.C(n_64),
.Y(n_1212)
);

AOI221xp5_ASAP7_75t_L g1213 ( 
.A1(n_1201),
.A2(n_832),
.B1(n_967),
.B2(n_959),
.C(n_942),
.Y(n_1213)
);

NOR4xp25_ASAP7_75t_L g1214 ( 
.A(n_1209),
.B(n_63),
.C(n_67),
.D(n_71),
.Y(n_1214)
);

NOR3xp33_ASAP7_75t_SL g1215 ( 
.A(n_1205),
.B(n_74),
.C(n_78),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_SL g1216 ( 
.A1(n_1204),
.A2(n_1207),
.B1(n_1200),
.B2(n_1210),
.Y(n_1216)
);

NOR3x2_ASAP7_75t_L g1217 ( 
.A(n_1198),
.B(n_79),
.C(n_82),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1202),
.Y(n_1218)
);

NAND5xp2_ASAP7_75t_L g1219 ( 
.A(n_1199),
.B(n_873),
.C(n_88),
.D(n_109),
.E(n_110),
.Y(n_1219)
);

XOR2xp5_ASAP7_75t_L g1220 ( 
.A(n_1211),
.B(n_86),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1203),
.A2(n_1206),
.B1(n_1208),
.B2(n_938),
.Y(n_1221)
);

AO21x2_ASAP7_75t_L g1222 ( 
.A1(n_1218),
.A2(n_1206),
.B(n_113),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1216),
.A2(n_938),
.B1(n_967),
.B2(n_959),
.Y(n_1223)
);

OA21x2_ASAP7_75t_L g1224 ( 
.A1(n_1215),
.A2(n_111),
.B(n_114),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1214),
.A2(n_942),
.B(n_974),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1212),
.A2(n_1220),
.B1(n_1221),
.B2(n_1213),
.Y(n_1226)
);

AOI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1219),
.A2(n_938),
.B1(n_942),
.B2(n_974),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1222),
.A2(n_1217),
.B1(n_938),
.B2(n_974),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1226),
.A2(n_873),
.B(n_932),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1224),
.A2(n_932),
.B1(n_924),
.B2(n_923),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1223),
.A2(n_116),
.B(n_122),
.Y(n_1231)
);

OAI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1231),
.A2(n_1227),
.B(n_1225),
.Y(n_1232)
);

XNOR2xp5_ASAP7_75t_L g1233 ( 
.A(n_1232),
.B(n_1228),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1233),
.A2(n_1230),
.B1(n_1229),
.B2(n_924),
.Y(n_1234)
);

OAI221xp5_ASAP7_75t_R g1235 ( 
.A1(n_1234),
.A2(n_126),
.B1(n_127),
.B2(n_130),
.C(n_131),
.Y(n_1235)
);

AOI211xp5_ASAP7_75t_L g1236 ( 
.A1(n_1235),
.A2(n_134),
.B(n_136),
.C(n_137),
.Y(n_1236)
);


endmodule