module real_jpeg_33816_n_27 (n_17, n_199, n_8, n_0, n_21, n_2, n_196, n_201, n_10, n_9, n_12, n_24, n_6, n_194, n_202, n_198, n_203, n_23, n_11, n_14, n_25, n_195, n_7, n_22, n_18, n_3, n_193, n_197, n_5, n_4, n_1, n_26, n_200, n_20, n_19, n_16, n_15, n_13, n_27);

input n_17;
input n_199;
input n_8;
input n_0;
input n_21;
input n_2;
input n_196;
input n_201;
input n_10;
input n_9;
input n_12;
input n_24;
input n_6;
input n_194;
input n_202;
input n_198;
input n_203;
input n_23;
input n_11;
input n_14;
input n_25;
input n_195;
input n_7;
input n_22;
input n_18;
input n_3;
input n_193;
input n_197;
input n_5;
input n_4;
input n_1;
input n_26;
input n_200;
input n_20;
input n_19;
input n_16;
input n_15;
input n_13;

output n_27;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_174;
wire n_87;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_0),
.B(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_0),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_1),
.B(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_1),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_2),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_2),
.B(n_77),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_3),
.B(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

AOI221xp5_ASAP7_75t_L g124 ( 
.A1(n_5),
.A2(n_6),
.B1(n_125),
.B2(n_130),
.C(n_132),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_5),
.B(n_125),
.C(n_130),
.Y(n_135)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_6),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_7),
.B(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_7),
.Y(n_167)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_8),
.Y(n_104)
);

AOI322xp5_ASAP7_75t_L g163 ( 
.A1(n_8),
.A2(n_98),
.A3(n_100),
.B1(n_106),
.B2(n_164),
.C1(n_166),
.C2(n_203),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_9),
.B(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_10),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_10),
.B(n_84),
.Y(n_186)
);

FAx1_ASAP7_75t_SL g27 ( 
.A(n_11),
.B(n_28),
.CI(n_35),
.CON(n_27),
.SN(n_27)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_12),
.Y(n_142)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_13),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_13),
.B(n_155),
.Y(n_165)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_14),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_14),
.B(n_108),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_15),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_16),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_17),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_18),
.B(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_20),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_20),
.B(n_114),
.Y(n_161)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_24),
.A2(n_38),
.B1(n_40),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_25),
.Y(n_144)
);

NOR2x1_ASAP7_75t_L g71 ( 
.A(n_26),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_26),
.B(n_72),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_34),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_34),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_89),
.B(n_169),
.Y(n_36)
);

NAND4xp25_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_51),
.C(n_75),
.D(n_82),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_50),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_47),
.Y(n_152)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

NOR3xp33_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_60),
.C(n_65),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND3xp33_ASAP7_75t_L g184 ( 
.A(n_53),
.B(n_185),
.C(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_59),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_54),
.B(n_59),
.Y(n_178)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_60),
.B(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_60),
.A2(n_184),
.B(n_187),
.Y(n_183)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_61),
.Y(n_176)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

AOI21xp33_ASAP7_75t_L g177 ( 
.A1(n_65),
.A2(n_173),
.B(n_178),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_71),
.Y(n_65)
);

INVxp67_ASAP7_75t_SL g188 ( 
.A(n_66),
.Y(n_188)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_67),
.Y(n_181)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_71),
.Y(n_185)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI31xp33_ASAP7_75t_L g182 ( 
.A1(n_75),
.A2(n_183),
.A3(n_188),
.B(n_189),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_76),
.A2(n_171),
.B(n_182),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

NOR2x1_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_115),
.Y(n_114)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_88),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_86),
.Y(n_85)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI31xp67_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_116),
.A3(n_153),
.B(n_159),
.Y(n_89)
);

NOR3xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_105),
.C(n_113),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_91),
.A2(n_160),
.B(n_163),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_98),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR3xp33_ASAP7_75t_L g164 ( 
.A(n_93),
.B(n_113),
.C(n_165),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_94),
.Y(n_168)
);

NOR2x1_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_104),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_194),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

OA21x2_ASAP7_75t_SL g160 ( 
.A1(n_105),
.A2(n_161),
.B(n_162),
.Y(n_160)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_112),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_144),
.C(n_145),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_136),
.B(n_143),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_124),
.B1(n_134),
.B2(n_135),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_126),
.B(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_199),
.Y(n_130)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_142),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_142),
.Y(n_143)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_158),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_177),
.B(n_179),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_193),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_195),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_196),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_197),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_198),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_200),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_201),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_202),
.Y(n_156)
);


endmodule