module real_aes_7518_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_0), .B(n_85), .C(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g124 ( .A(n_0), .Y(n_124) );
A2O1A1Ixp33_ASAP7_75t_L g456 ( .A1(n_1), .A2(n_145), .B(n_157), .C(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g264 ( .A(n_2), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_3), .A2(n_172), .B(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_4), .B(n_168), .Y(n_501) );
AOI21xp33_ASAP7_75t_L g171 ( .A1(n_5), .A2(n_172), .B(n_173), .Y(n_171) );
AND2x6_ASAP7_75t_L g145 ( .A(n_6), .B(n_146), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_7), .A2(n_240), .B(n_241), .Y(n_239) );
INVx1_ASAP7_75t_L g106 ( .A(n_8), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_8), .B(n_39), .Y(n_125) );
INVx1_ASAP7_75t_L g472 ( .A(n_9), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_10), .B(n_178), .Y(n_460) );
INVx1_ASAP7_75t_L g180 ( .A(n_11), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_12), .B(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g142 ( .A(n_13), .Y(n_142) );
INVx1_ASAP7_75t_L g246 ( .A(n_14), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_15), .A2(n_181), .B(n_247), .C(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_16), .B(n_168), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_17), .B(n_191), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_18), .B(n_172), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_19), .B(n_514), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_20), .A2(n_148), .B(n_232), .C(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_21), .B(n_168), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_22), .B(n_178), .Y(n_535) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_23), .A2(n_244), .B(n_245), .C(n_247), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_24), .B(n_178), .Y(n_522) );
CKINVDCx16_ASAP7_75t_R g531 ( .A(n_25), .Y(n_531) );
INVx1_ASAP7_75t_L g521 ( .A(n_26), .Y(n_521) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_27), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_28), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_29), .B(n_178), .Y(n_265) );
INVx1_ASAP7_75t_L g510 ( .A(n_30), .Y(n_510) );
INVx1_ASAP7_75t_L g156 ( .A(n_31), .Y(n_156) );
INVx2_ASAP7_75t_L g150 ( .A(n_32), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_33), .Y(n_462) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_34), .A2(n_182), .B(n_232), .C(n_499), .Y(n_498) );
INVxp67_ASAP7_75t_L g511 ( .A(n_35), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_36), .A2(n_145), .B(n_157), .C(n_202), .Y(n_201) );
CKINVDCx14_ASAP7_75t_R g497 ( .A(n_37), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_38), .A2(n_157), .B(n_520), .C(n_524), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_39), .B(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g154 ( .A(n_40), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_41), .A2(n_177), .B(n_207), .C(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_42), .B(n_178), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_43), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_44), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_45), .Y(n_126) );
INVx1_ASAP7_75t_L g487 ( .A(n_46), .Y(n_487) );
CKINVDCx16_ASAP7_75t_R g160 ( .A(n_47), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_48), .B(n_172), .Y(n_234) );
AOI222xp33_ASAP7_75t_SL g127 ( .A1(n_49), .A2(n_58), .B1(n_128), .B2(n_714), .C1(n_715), .C2(n_719), .Y(n_127) );
AOI22xp5_ASAP7_75t_L g147 ( .A1(n_50), .A2(n_148), .B1(n_151), .B2(n_157), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_51), .Y(n_211) );
CKINVDCx16_ASAP7_75t_R g261 ( .A(n_52), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g176 ( .A1(n_53), .A2(n_177), .B(n_179), .C(n_182), .Y(n_176) );
CKINVDCx14_ASAP7_75t_R g469 ( .A(n_54), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_55), .Y(n_221) );
INVx1_ASAP7_75t_L g174 ( .A(n_56), .Y(n_174) );
INVx1_ASAP7_75t_L g146 ( .A(n_57), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_58), .Y(n_714) );
INVx1_ASAP7_75t_L g141 ( .A(n_59), .Y(n_141) );
INVx1_ASAP7_75t_SL g500 ( .A(n_60), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_61), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_62), .B(n_168), .Y(n_491) );
OAI22xp5_ASAP7_75t_SL g724 ( .A1(n_63), .A2(n_446), .B1(n_716), .B2(n_725), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_63), .Y(n_725) );
INVx1_ASAP7_75t_L g534 ( .A(n_64), .Y(n_534) );
A2O1A1Ixp33_ASAP7_75t_SL g190 ( .A1(n_65), .A2(n_182), .B(n_191), .C(n_192), .Y(n_190) );
INVxp67_ASAP7_75t_L g193 ( .A(n_66), .Y(n_193) );
INVx1_ASAP7_75t_L g110 ( .A(n_67), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_68), .A2(n_172), .B(n_468), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_69), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_70), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_71), .A2(n_172), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g214 ( .A(n_72), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_73), .A2(n_240), .B(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g479 ( .A(n_74), .Y(n_479) );
CKINVDCx16_ASAP7_75t_R g518 ( .A(n_75), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_76), .A2(n_145), .B(n_157), .C(n_216), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_77), .A2(n_172), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g482 ( .A(n_78), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_79), .A2(n_100), .B1(n_111), .B2(n_728), .Y(n_99) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_80), .B(n_204), .Y(n_203) );
INVx2_ASAP7_75t_L g139 ( .A(n_81), .Y(n_139) );
INVx1_ASAP7_75t_L g458 ( .A(n_82), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_83), .B(n_191), .Y(n_205) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_84), .A2(n_145), .B(n_157), .C(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g121 ( .A(n_85), .B(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g445 ( .A(n_85), .Y(n_445) );
OR2x2_ASAP7_75t_L g713 ( .A(n_85), .B(n_123), .Y(n_713) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_86), .A2(n_157), .B(n_533), .C(n_536), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_87), .B(n_185), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g268 ( .A(n_88), .Y(n_268) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_89), .A2(n_145), .B(n_157), .C(n_229), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_90), .Y(n_236) );
INVx1_ASAP7_75t_L g189 ( .A(n_91), .Y(n_189) );
CKINVDCx16_ASAP7_75t_R g242 ( .A(n_92), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_93), .B(n_204), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_94), .B(n_170), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_95), .B(n_170), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_96), .B(n_110), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_97), .A2(n_172), .B(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g490 ( .A(n_98), .Y(n_490) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_102), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_103), .Y(n_729) );
CKINVDCx9p33_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_105), .B(n_107), .Y(n_104) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AOI22xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_127), .B1(n_722), .B2(n_723), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_114), .B(n_118), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_SL g722 ( .A(n_115), .Y(n_722) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g723 ( .A1(n_118), .A2(n_724), .B(n_726), .Y(n_723) );
NOR2xp33_ASAP7_75t_SL g118 ( .A(n_119), .B(n_126), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_SL g727 ( .A(n_121), .Y(n_727) );
NOR2x2_ASAP7_75t_L g721 ( .A(n_122), .B(n_445), .Y(n_721) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g444 ( .A(n_123), .B(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
OAI22xp5_ASAP7_75t_SL g128 ( .A1(n_129), .A2(n_442), .B1(n_446), .B2(n_713), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OAI22xp5_ASAP7_75t_SL g715 ( .A1(n_130), .A2(n_442), .B1(n_716), .B2(n_717), .Y(n_715) );
AND3x1_ASAP7_75t_L g130 ( .A(n_131), .B(n_367), .C(n_416), .Y(n_130) );
NOR3xp33_ASAP7_75t_SL g131 ( .A(n_132), .B(n_274), .C(n_312), .Y(n_131) );
OAI222xp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_195), .B1(n_249), .B2(n_255), .C1(n_269), .C2(n_272), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_166), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_134), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_134), .B(n_317), .Y(n_408) );
BUFx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OR2x2_ASAP7_75t_L g285 ( .A(n_135), .B(n_186), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_135), .B(n_167), .Y(n_293) );
AND2x2_ASAP7_75t_L g328 ( .A(n_135), .B(n_305), .Y(n_328) );
OR2x2_ASAP7_75t_L g352 ( .A(n_135), .B(n_167), .Y(n_352) );
OR2x2_ASAP7_75t_L g360 ( .A(n_135), .B(n_259), .Y(n_360) );
AND2x2_ASAP7_75t_L g363 ( .A(n_135), .B(n_186), .Y(n_363) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
OR2x2_ASAP7_75t_L g257 ( .A(n_136), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g271 ( .A(n_136), .B(n_186), .Y(n_271) );
AND2x2_ASAP7_75t_L g321 ( .A(n_136), .B(n_259), .Y(n_321) );
AND2x2_ASAP7_75t_L g334 ( .A(n_136), .B(n_167), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_136), .B(n_420), .Y(n_441) );
AO21x2_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_143), .B(n_164), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_137), .B(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g209 ( .A(n_137), .Y(n_209) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_137), .A2(n_260), .B(n_267), .Y(n_259) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_138), .Y(n_170) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x2_ASAP7_75t_SL g185 ( .A(n_139), .B(n_140), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
OAI22xp33_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_147), .B1(n_160), .B2(n_161), .Y(n_143) );
O2A1O1Ixp33_ASAP7_75t_L g173 ( .A1(n_144), .A2(n_174), .B(n_175), .C(n_176), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_L g188 ( .A1(n_144), .A2(n_175), .B(n_189), .C(n_190), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g241 ( .A1(n_144), .A2(n_175), .B(n_242), .C(n_243), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_SL g468 ( .A1(n_144), .A2(n_175), .B(n_469), .C(n_470), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_SL g478 ( .A1(n_144), .A2(n_175), .B(n_479), .C(n_480), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_SL g486 ( .A1(n_144), .A2(n_175), .B(n_487), .C(n_488), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_L g496 ( .A1(n_144), .A2(n_175), .B(n_497), .C(n_498), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_SL g506 ( .A1(n_144), .A2(n_175), .B(n_507), .C(n_508), .Y(n_506) );
INVx1_ASAP7_75t_L g536 ( .A(n_144), .Y(n_536) );
INVx4_ASAP7_75t_SL g144 ( .A(n_145), .Y(n_144) );
NAND2x1p5_ASAP7_75t_L g161 ( .A(n_145), .B(n_162), .Y(n_161) );
AND2x4_ASAP7_75t_L g172 ( .A(n_145), .B(n_162), .Y(n_172) );
BUFx3_ASAP7_75t_L g524 ( .A(n_145), .Y(n_524) );
INVx2_ASAP7_75t_L g266 ( .A(n_148), .Y(n_266) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g158 ( .A(n_150), .Y(n_158) );
INVx1_ASAP7_75t_L g163 ( .A(n_150), .Y(n_163) );
OAI22xp5_ASAP7_75t_SL g151 ( .A1(n_152), .A2(n_154), .B1(n_155), .B2(n_156), .Y(n_151) );
INVx2_ASAP7_75t_L g155 ( .A(n_152), .Y(n_155) );
INVx4_ASAP7_75t_L g244 ( .A(n_152), .Y(n_244) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g159 ( .A(n_153), .Y(n_159) );
AND2x2_ASAP7_75t_L g162 ( .A(n_153), .B(n_163), .Y(n_162) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_153), .Y(n_178) );
INVx3_ASAP7_75t_L g181 ( .A(n_153), .Y(n_181) );
INVx1_ASAP7_75t_L g191 ( .A(n_153), .Y(n_191) );
INVx2_ASAP7_75t_L g459 ( .A(n_155), .Y(n_459) );
INVx5_ASAP7_75t_L g175 ( .A(n_157), .Y(n_175) );
AND2x6_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_158), .Y(n_183) );
BUFx3_ASAP7_75t_L g208 ( .A(n_158), .Y(n_208) );
OAI21xp5_ASAP7_75t_L g213 ( .A1(n_161), .A2(n_214), .B(n_215), .Y(n_213) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_161), .A2(n_261), .B(n_262), .Y(n_260) );
OAI21xp5_ASAP7_75t_L g454 ( .A1(n_161), .A2(n_455), .B(n_456), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_L g517 ( .A1(n_161), .A2(n_185), .B(n_518), .C(n_519), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g530 ( .A1(n_161), .A2(n_531), .B(n_532), .Y(n_530) );
INVx1_ASAP7_75t_L g512 ( .A(n_163), .Y(n_512) );
O2A1O1Ixp33_ASAP7_75t_L g359 ( .A1(n_166), .A2(n_360), .B(n_361), .C(n_364), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_166), .B(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_166), .B(n_304), .Y(n_426) );
AND2x2_ASAP7_75t_L g166 ( .A(n_167), .B(n_186), .Y(n_166) );
AND2x2_ASAP7_75t_SL g270 ( .A(n_167), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g284 ( .A(n_167), .Y(n_284) );
AND2x2_ASAP7_75t_L g311 ( .A(n_167), .B(n_305), .Y(n_311) );
INVx1_ASAP7_75t_SL g319 ( .A(n_167), .Y(n_319) );
AND2x2_ASAP7_75t_L g342 ( .A(n_167), .B(n_343), .Y(n_342) );
BUFx2_ASAP7_75t_L g420 ( .A(n_167), .Y(n_420) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_171), .B(n_184), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_SL g210 ( .A(n_169), .B(n_211), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_169), .B(n_462), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_169), .B(n_526), .Y(n_525) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_169), .A2(n_530), .B(n_537), .Y(n_529) );
INVx4_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_170), .A2(n_187), .B(n_194), .Y(n_186) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_170), .Y(n_476) );
BUFx2_ASAP7_75t_L g240 ( .A(n_172), .Y(n_240) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx4_ASAP7_75t_L g232 ( .A(n_178), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_181), .B(n_193), .Y(n_192) );
INVx5_ASAP7_75t_L g204 ( .A(n_181), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_181), .B(n_472), .Y(n_471) );
INVx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_183), .Y(n_233) );
INVx1_ASAP7_75t_L g222 ( .A(n_185), .Y(n_222) );
INVx2_ASAP7_75t_L g226 ( .A(n_185), .Y(n_226) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_185), .A2(n_239), .B(n_248), .Y(n_238) );
OA21x2_ASAP7_75t_L g466 ( .A1(n_185), .A2(n_467), .B(n_473), .Y(n_466) );
BUFx2_ASAP7_75t_L g256 ( .A(n_186), .Y(n_256) );
INVx1_ASAP7_75t_L g318 ( .A(n_186), .Y(n_318) );
INVx3_ASAP7_75t_L g343 ( .A(n_186), .Y(n_343) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_195), .B(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_223), .Y(n_195) );
INVx1_ASAP7_75t_L g339 ( .A(n_196), .Y(n_339) );
OAI32xp33_ASAP7_75t_L g345 ( .A1(n_196), .A2(n_284), .A3(n_346), .B1(n_347), .B2(n_348), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_196), .A2(n_350), .B1(n_353), .B2(n_358), .Y(n_349) );
INVx4_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g287 ( .A(n_197), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g365 ( .A(n_197), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g435 ( .A(n_197), .B(n_381), .Y(n_435) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_212), .Y(n_197) );
AND2x2_ASAP7_75t_L g250 ( .A(n_198), .B(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g280 ( .A(n_198), .Y(n_280) );
INVx1_ASAP7_75t_L g299 ( .A(n_198), .Y(n_299) );
OR2x2_ASAP7_75t_L g307 ( .A(n_198), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g314 ( .A(n_198), .B(n_288), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_198), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g335 ( .A(n_198), .B(n_253), .Y(n_335) );
INVx3_ASAP7_75t_L g357 ( .A(n_198), .Y(n_357) );
AND2x2_ASAP7_75t_L g382 ( .A(n_198), .B(n_254), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_198), .B(n_347), .Y(n_430) );
OR2x6_ASAP7_75t_L g198 ( .A(n_199), .B(n_210), .Y(n_198) );
AOI21xp5_ASAP7_75t_SL g199 ( .A1(n_200), .A2(n_201), .B(n_209), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_205), .B(n_206), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_204), .A2(n_264), .B(n_265), .C(n_266), .Y(n_263) );
OAI22xp33_ASAP7_75t_L g509 ( .A1(n_204), .A2(n_244), .B1(n_510), .B2(n_511), .Y(n_509) );
O2A1O1Ixp33_ASAP7_75t_L g520 ( .A1(n_204), .A2(n_521), .B(n_522), .C(n_523), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_206), .A2(n_217), .B(n_218), .Y(n_216) );
O2A1O1Ixp5_ASAP7_75t_L g457 ( .A1(n_206), .A2(n_458), .B(n_459), .C(n_460), .Y(n_457) );
O2A1O1Ixp33_ASAP7_75t_L g533 ( .A1(n_206), .A2(n_459), .B(n_534), .C(n_535), .Y(n_533) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g247 ( .A(n_208), .Y(n_247) );
INVx1_ASAP7_75t_L g219 ( .A(n_209), .Y(n_219) );
INVx2_ASAP7_75t_L g254 ( .A(n_212), .Y(n_254) );
AND2x2_ASAP7_75t_L g386 ( .A(n_212), .B(n_224), .Y(n_386) );
AO21x2_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_219), .B(n_220), .Y(n_212) );
INVx1_ASAP7_75t_L g504 ( .A(n_219), .Y(n_504) );
AO21x2_ASAP7_75t_L g556 ( .A1(n_219), .A2(n_557), .B(n_558), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_222), .B(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_222), .B(n_268), .Y(n_267) );
AO21x2_ASAP7_75t_L g453 ( .A1(n_222), .A2(n_454), .B(n_461), .Y(n_453) );
INVx2_ASAP7_75t_L g428 ( .A(n_223), .Y(n_428) );
OR2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_237), .Y(n_223) );
INVx1_ASAP7_75t_L g273 ( .A(n_224), .Y(n_273) );
AND2x2_ASAP7_75t_L g300 ( .A(n_224), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_224), .B(n_254), .Y(n_308) );
AND2x2_ASAP7_75t_L g366 ( .A(n_224), .B(n_289), .Y(n_366) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g252 ( .A(n_225), .Y(n_252) );
AND2x2_ASAP7_75t_L g279 ( .A(n_225), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g288 ( .A(n_225), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_225), .B(n_254), .Y(n_354) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_235), .Y(n_225) );
INVx1_ASAP7_75t_L g514 ( .A(n_226), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_226), .B(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_228), .B(n_234), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_233), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_232), .B(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_237), .B(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g301 ( .A(n_237), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_237), .B(n_254), .Y(n_347) );
AND2x2_ASAP7_75t_L g356 ( .A(n_237), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g381 ( .A(n_237), .Y(n_381) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g253 ( .A(n_238), .B(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g289 ( .A(n_238), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_244), .B(n_246), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_244), .B(n_482), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_244), .B(n_490), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_249), .A2(n_259), .B1(n_418), .B2(n_421), .Y(n_417) );
INVx1_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
OAI21xp5_ASAP7_75t_SL g440 ( .A1(n_251), .A2(n_362), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_252), .B(n_357), .Y(n_374) );
INVx1_ASAP7_75t_L g399 ( .A(n_252), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_253), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g326 ( .A(n_253), .B(n_279), .Y(n_326) );
INVx2_ASAP7_75t_L g282 ( .A(n_254), .Y(n_282) );
INVx1_ASAP7_75t_L g332 ( .A(n_254), .Y(n_332) );
OAI221xp5_ASAP7_75t_L g423 ( .A1(n_255), .A2(n_407), .B1(n_424), .B2(n_427), .C(n_429), .Y(n_423) );
OR2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
INVx1_ASAP7_75t_L g294 ( .A(n_256), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_256), .B(n_305), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_257), .B(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g348 ( .A(n_257), .B(n_294), .Y(n_348) );
INVx3_ASAP7_75t_SL g389 ( .A(n_257), .Y(n_389) );
AND2x2_ASAP7_75t_L g333 ( .A(n_258), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g362 ( .A(n_258), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_258), .B(n_271), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_258), .B(n_317), .Y(n_403) );
INVx3_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx3_ASAP7_75t_L g305 ( .A(n_259), .Y(n_305) );
OAI322xp33_ASAP7_75t_L g400 ( .A1(n_259), .A2(n_331), .A3(n_353), .B1(n_401), .B2(n_403), .C1(n_404), .C2(n_405), .Y(n_400) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AOI21xp33_ASAP7_75t_L g424 ( .A1(n_270), .A2(n_273), .B(n_425), .Y(n_424) );
NOR2xp33_ASAP7_75t_SL g350 ( .A(n_271), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g372 ( .A(n_271), .B(n_284), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_271), .B(n_311), .Y(n_387) );
INVxp67_ASAP7_75t_L g338 ( .A(n_273), .Y(n_338) );
AOI211xp5_ASAP7_75t_L g344 ( .A1(n_273), .A2(n_345), .B(n_349), .C(n_359), .Y(n_344) );
OAI221xp5_ASAP7_75t_SL g274 ( .A1(n_275), .A2(n_283), .B1(n_286), .B2(n_290), .C(n_295), .Y(n_274) );
INVxp67_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_281), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g298 ( .A(n_282), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g415 ( .A(n_282), .Y(n_415) );
OAI221xp5_ASAP7_75t_L g431 ( .A1(n_283), .A2(n_432), .B1(n_437), .B2(n_438), .C(n_440), .Y(n_431) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_284), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_SL g331 ( .A(n_284), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_284), .B(n_362), .Y(n_369) );
AND2x2_ASAP7_75t_L g411 ( .A(n_284), .B(n_389), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_285), .B(n_310), .Y(n_309) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_285), .A2(n_297), .B1(n_407), .B2(n_408), .Y(n_406) );
OR2x2_ASAP7_75t_L g437 ( .A(n_285), .B(n_305), .Y(n_437) );
CKINVDCx16_ASAP7_75t_R g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g414 ( .A(n_288), .Y(n_414) );
AND2x2_ASAP7_75t_L g439 ( .A(n_288), .B(n_382), .Y(n_439) );
INVxp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_SL g291 ( .A(n_292), .B(n_294), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g303 ( .A(n_293), .B(n_304), .Y(n_303) );
AOI22xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_302), .B1(n_306), .B2(n_309), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_300), .Y(n_297) );
INVx1_ASAP7_75t_L g370 ( .A(n_298), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_298), .B(n_338), .Y(n_405) );
AOI322xp5_ASAP7_75t_L g329 ( .A1(n_300), .A2(n_330), .A3(n_332), .B1(n_333), .B2(n_335), .C1(n_336), .C2(n_340), .Y(n_329) );
INVxp67_ASAP7_75t_L g323 ( .A(n_301), .Y(n_323) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g324 ( .A1(n_303), .A2(n_308), .B1(n_325), .B2(n_327), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_304), .B(n_317), .Y(n_404) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_305), .B(n_343), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_305), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g401 ( .A(n_307), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
NAND3xp33_ASAP7_75t_SL g312 ( .A(n_313), .B(n_329), .C(n_344), .Y(n_312) );
AOI221xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_315), .B1(n_320), .B2(n_322), .C(n_324), .Y(n_313) );
AND2x2_ASAP7_75t_L g320 ( .A(n_316), .B(n_321), .Y(n_320) );
INVx3_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
AND2x2_ASAP7_75t_L g330 ( .A(n_321), .B(n_331), .Y(n_330) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_323), .Y(n_402) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_328), .B(n_342), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_331), .B(n_389), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_332), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_SL g407 ( .A(n_335), .Y(n_407) );
AND2x2_ASAP7_75t_L g422 ( .A(n_335), .B(n_399), .Y(n_422) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AOI211xp5_ASAP7_75t_L g416 ( .A1(n_346), .A2(n_417), .B(n_423), .C(n_431), .Y(n_416) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g385 ( .A(n_356), .B(n_386), .Y(n_385) );
NAND2x1_ASAP7_75t_SL g427 ( .A(n_357), .B(n_428), .Y(n_427) );
CKINVDCx16_ASAP7_75t_R g397 ( .A(n_360), .Y(n_397) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g392 ( .A(n_366), .Y(n_392) );
AND2x2_ASAP7_75t_L g396 ( .A(n_366), .B(n_382), .Y(n_396) );
NOR5xp2_ASAP7_75t_L g367 ( .A(n_368), .B(n_383), .C(n_400), .D(n_406), .E(n_409), .Y(n_367) );
OAI221xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_370), .B1(n_371), .B2(n_373), .C(n_375), .Y(n_368) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_372), .B(n_430), .Y(n_429) );
INVxp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_376), .B(n_378), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g398 ( .A(n_382), .B(n_399), .Y(n_398) );
OAI221xp5_ASAP7_75t_SL g383 ( .A1(n_384), .A2(n_387), .B1(n_388), .B2(n_390), .C(n_393), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_396), .B1(n_397), .B2(n_398), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g436 ( .A(n_396), .Y(n_436) );
AOI211xp5_ASAP7_75t_SL g409 ( .A1(n_410), .A2(n_412), .B(n_414), .C(n_415), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVxp67_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_434), .B(n_436), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
CKINVDCx14_ASAP7_75t_R g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g716 ( .A(n_446), .Y(n_716) );
OR2x2_ASAP7_75t_SL g446 ( .A(n_447), .B(n_668), .Y(n_446) );
NAND5xp2_ASAP7_75t_L g447 ( .A(n_448), .B(n_580), .C(n_618), .D(n_639), .E(n_656), .Y(n_447) );
NOR3xp33_ASAP7_75t_L g448 ( .A(n_449), .B(n_552), .C(n_573), .Y(n_448) );
OAI221xp5_ASAP7_75t_SL g449 ( .A1(n_450), .A2(n_492), .B1(n_515), .B2(n_539), .C(n_543), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_463), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_452), .B(n_541), .Y(n_560) );
OR2x2_ASAP7_75t_L g587 ( .A(n_452), .B(n_475), .Y(n_587) );
AND2x2_ASAP7_75t_L g601 ( .A(n_452), .B(n_475), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_452), .B(n_466), .Y(n_615) );
AND2x2_ASAP7_75t_L g653 ( .A(n_452), .B(n_617), .Y(n_653) );
AND2x2_ASAP7_75t_L g682 ( .A(n_452), .B(n_592), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_452), .B(n_564), .Y(n_699) );
INVx4_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g579 ( .A(n_453), .B(n_474), .Y(n_579) );
BUFx3_ASAP7_75t_L g604 ( .A(n_453), .Y(n_604) );
AND2x2_ASAP7_75t_L g633 ( .A(n_453), .B(n_475), .Y(n_633) );
AND3x2_ASAP7_75t_L g646 ( .A(n_453), .B(n_647), .C(n_648), .Y(n_646) );
INVx1_ASAP7_75t_L g569 ( .A(n_463), .Y(n_569) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_474), .Y(n_463) );
AOI32xp33_ASAP7_75t_L g624 ( .A1(n_464), .A2(n_576), .A3(n_625), .B1(n_628), .B2(n_629), .Y(n_624) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g551 ( .A(n_465), .B(n_474), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_465), .B(n_579), .Y(n_622) );
AND2x2_ASAP7_75t_L g629 ( .A(n_465), .B(n_601), .Y(n_629) );
OR2x2_ASAP7_75t_L g635 ( .A(n_465), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_465), .B(n_590), .Y(n_660) );
OR2x2_ASAP7_75t_L g678 ( .A(n_465), .B(n_503), .Y(n_678) );
BUFx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g542 ( .A(n_466), .B(n_484), .Y(n_542) );
INVx2_ASAP7_75t_L g564 ( .A(n_466), .Y(n_564) );
OR2x2_ASAP7_75t_L g586 ( .A(n_466), .B(n_484), .Y(n_586) );
AND2x2_ASAP7_75t_L g591 ( .A(n_466), .B(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_466), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g647 ( .A(n_466), .B(n_541), .Y(n_647) );
INVx1_ASAP7_75t_SL g698 ( .A(n_474), .Y(n_698) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_484), .Y(n_474) );
INVx1_ASAP7_75t_SL g541 ( .A(n_475), .Y(n_541) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_475), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_475), .B(n_627), .Y(n_626) );
NAND3xp33_ASAP7_75t_L g693 ( .A(n_475), .B(n_564), .C(n_682), .Y(n_693) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B(n_483), .Y(n_475) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_476), .A2(n_485), .B(n_491), .Y(n_484) );
OA21x2_ASAP7_75t_L g494 ( .A1(n_476), .A2(n_495), .B(n_501), .Y(n_494) );
INVx2_ASAP7_75t_L g592 ( .A(n_484), .Y(n_592) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_484), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_502), .Y(n_492) );
INVx1_ASAP7_75t_L g628 ( .A(n_493), .Y(n_628) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g546 ( .A(n_494), .B(n_528), .Y(n_546) );
INVx2_ASAP7_75t_L g563 ( .A(n_494), .Y(n_563) );
AND2x2_ASAP7_75t_L g568 ( .A(n_494), .B(n_529), .Y(n_568) );
AND2x2_ASAP7_75t_L g583 ( .A(n_494), .B(n_516), .Y(n_583) );
AND2x2_ASAP7_75t_L g595 ( .A(n_494), .B(n_567), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_502), .B(n_611), .Y(n_610) );
NAND2x1p5_ASAP7_75t_L g667 ( .A(n_502), .B(n_568), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_502), .B(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_502), .B(n_562), .Y(n_690) );
BUFx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OR2x2_ASAP7_75t_L g527 ( .A(n_503), .B(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_503), .B(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g572 ( .A(n_503), .B(n_516), .Y(n_572) );
AND2x2_ASAP7_75t_L g598 ( .A(n_503), .B(n_528), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_503), .B(n_638), .Y(n_637) );
OA21x2_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_505), .B(n_513), .Y(n_503) );
INVx1_ASAP7_75t_L g557 ( .A(n_505), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_509), .B(n_512), .Y(n_508) );
INVx2_ASAP7_75t_L g523 ( .A(n_512), .Y(n_523) );
INVx1_ASAP7_75t_L g558 ( .A(n_513), .Y(n_558) );
OR2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_527), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_516), .B(n_549), .Y(n_548) );
AND2x4_ASAP7_75t_L g562 ( .A(n_516), .B(n_563), .Y(n_562) );
INVx3_ASAP7_75t_SL g567 ( .A(n_516), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_516), .B(n_554), .Y(n_620) );
OR2x2_ASAP7_75t_L g630 ( .A(n_516), .B(n_556), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_516), .B(n_598), .Y(n_658) );
OR2x2_ASAP7_75t_L g688 ( .A(n_516), .B(n_528), .Y(n_688) );
AND2x2_ASAP7_75t_L g692 ( .A(n_516), .B(n_529), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_516), .B(n_568), .Y(n_705) );
AND2x2_ASAP7_75t_L g712 ( .A(n_516), .B(n_594), .Y(n_712) );
OR2x6_ASAP7_75t_L g516 ( .A(n_517), .B(n_525), .Y(n_516) );
INVx1_ASAP7_75t_SL g655 ( .A(n_527), .Y(n_655) );
AND2x2_ASAP7_75t_L g594 ( .A(n_528), .B(n_556), .Y(n_594) );
AND2x2_ASAP7_75t_L g608 ( .A(n_528), .B(n_563), .Y(n_608) );
AND2x2_ASAP7_75t_L g611 ( .A(n_528), .B(n_567), .Y(n_611) );
INVx1_ASAP7_75t_L g638 ( .A(n_528), .Y(n_638) );
INVx2_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
BUFx2_ASAP7_75t_L g550 ( .A(n_529), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_542), .Y(n_539) );
A2O1A1Ixp33_ASAP7_75t_L g709 ( .A1(n_540), .A2(n_586), .B(n_710), .C(n_711), .Y(n_709) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g616 ( .A(n_541), .B(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_542), .B(n_559), .Y(n_574) );
AND2x2_ASAP7_75t_L g600 ( .A(n_542), .B(n_601), .Y(n_600) );
OAI21xp5_ASAP7_75t_SL g543 ( .A1(n_544), .A2(n_547), .B(n_551), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_545), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g571 ( .A(n_546), .B(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_546), .B(n_567), .Y(n_612) );
AND2x2_ASAP7_75t_L g703 ( .A(n_546), .B(n_554), .Y(n_703) );
INVxp67_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g576 ( .A(n_550), .B(n_563), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_550), .B(n_561), .Y(n_577) );
OAI322xp33_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_560), .A3(n_561), .B1(n_564), .B2(n_565), .C1(n_569), .C2(n_570), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_559), .Y(n_553) );
AND2x2_ASAP7_75t_L g664 ( .A(n_554), .B(n_576), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_554), .B(n_628), .Y(n_710) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g607 ( .A(n_556), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OR2x2_ASAP7_75t_L g673 ( .A(n_560), .B(n_586), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_561), .B(n_655), .Y(n_654) );
INVx3_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_562), .B(n_594), .Y(n_651) );
AND2x2_ASAP7_75t_L g597 ( .A(n_563), .B(n_567), .Y(n_597) );
AND2x2_ASAP7_75t_L g605 ( .A(n_564), .B(n_606), .Y(n_605) );
A2O1A1Ixp33_ASAP7_75t_L g702 ( .A1(n_564), .A2(n_643), .B(n_703), .C(n_704), .Y(n_702) );
AOI21xp33_ASAP7_75t_L g675 ( .A1(n_565), .A2(n_578), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_567), .B(n_594), .Y(n_634) );
AND2x2_ASAP7_75t_L g640 ( .A(n_567), .B(n_608), .Y(n_640) );
AND2x2_ASAP7_75t_L g674 ( .A(n_567), .B(n_576), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_568), .B(n_583), .Y(n_582) );
INVx2_ASAP7_75t_SL g684 ( .A(n_568), .Y(n_684) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_572), .A2(n_600), .B1(n_602), .B2(n_607), .Y(n_599) );
OAI22xp5_ASAP7_75t_SL g573 ( .A1(n_574), .A2(n_575), .B1(n_577), .B2(n_578), .Y(n_573) );
OAI22xp33_ASAP7_75t_L g609 ( .A1(n_574), .A2(n_610), .B1(n_612), .B2(n_613), .Y(n_609) );
INVxp67_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_579), .A2(n_681), .B1(n_683), .B2(n_685), .C(n_689), .Y(n_680) );
AOI211xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_584), .B(n_588), .C(n_609), .Y(n_580) );
INVxp67_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
OR2x2_ASAP7_75t_L g650 ( .A(n_586), .B(n_603), .Y(n_650) );
INVx1_ASAP7_75t_L g701 ( .A(n_586), .Y(n_701) );
OAI221xp5_ASAP7_75t_L g588 ( .A1(n_587), .A2(n_589), .B1(n_593), .B2(n_596), .C(n_599), .Y(n_588) );
INVx2_ASAP7_75t_SL g643 ( .A(n_587), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
INVx1_ASAP7_75t_L g708 ( .A(n_590), .Y(n_708) );
AND2x2_ASAP7_75t_L g632 ( .A(n_591), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g617 ( .A(n_592), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
INVx1_ASAP7_75t_L g679 ( .A(n_595), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_605), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_603), .B(n_705), .Y(n_704) );
CKINVDCx16_ASAP7_75t_R g603 ( .A(n_604), .Y(n_603) );
INVxp67_ASAP7_75t_L g648 ( .A(n_606), .Y(n_648) );
O2A1O1Ixp33_ASAP7_75t_L g618 ( .A1(n_607), .A2(n_619), .B(n_621), .C(n_623), .Y(n_618) );
INVx1_ASAP7_75t_L g696 ( .A(n_610), .Y(n_696) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_614), .B(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
INVx2_ASAP7_75t_L g627 ( .A(n_617), .Y(n_627) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OAI222xp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_630), .B1(n_631), .B2(n_634), .C1(n_635), .C2(n_637), .Y(n_623) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_SL g663 ( .A(n_627), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_630), .B(n_684), .Y(n_683) );
NAND2xp33_ASAP7_75t_SL g661 ( .A(n_631), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_SL g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_SL g636 ( .A(n_633), .Y(n_636) );
AND2x2_ASAP7_75t_L g700 ( .A(n_633), .B(n_701), .Y(n_700) );
OR2x2_ASAP7_75t_L g666 ( .A(n_636), .B(n_663), .Y(n_666) );
INVx1_ASAP7_75t_L g695 ( .A(n_637), .Y(n_695) );
AOI211xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_641), .B(n_644), .C(n_649), .Y(n_639) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_643), .B(n_663), .Y(n_662) );
INVx2_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
AOI322xp5_ASAP7_75t_L g694 ( .A1(n_646), .A2(n_674), .A3(n_679), .B1(n_695), .B2(n_696), .C1(n_697), .C2(n_700), .Y(n_694) );
AND2x2_ASAP7_75t_L g681 ( .A(n_647), .B(n_682), .Y(n_681) );
OAI22xp33_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_651), .B1(n_652), .B2(n_654), .Y(n_649) );
INVxp33_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_659), .B1(n_661), .B2(n_664), .C(n_665), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
NAND5xp2_ASAP7_75t_L g668 ( .A(n_669), .B(n_680), .C(n_694), .D(n_702), .E(n_706), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_674), .B(n_675), .Y(n_669) );
INVxp67_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVxp33_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
A2O1A1Ixp33_ASAP7_75t_L g706 ( .A1(n_682), .A2(n_707), .B(n_708), .C(n_709), .Y(n_706) );
AOI31xp33_ASAP7_75t_L g689 ( .A1(n_684), .A2(n_690), .A3(n_691), .B(n_693), .Y(n_689) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
INVx1_ASAP7_75t_L g707 ( .A(n_705), .Y(n_707) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g718 ( .A(n_713), .Y(n_718) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_729), .Y(n_728) );
endmodule