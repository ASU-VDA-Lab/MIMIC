module fake_aes_7270_n_1359 (n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_292, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_297, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_291, n_170, n_294, n_40, n_111, n_157, n_296, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_295, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_298, n_283, n_299, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_293, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_290, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1359);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_292;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_297;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_291;
input n_170;
input n_294;
input n_40;
input n_111;
input n_157;
input n_296;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_295;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_298;
input n_283;
input n_299;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_293;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1359;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_1328;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1079;
wire n_315;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_994;
wire n_930;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_303;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_1350;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
wire n_1291;
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_213), .Y(n_300) );
INVxp33_ASAP7_75t_SL g301 ( .A(n_154), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_147), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_239), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_233), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_23), .Y(n_305) );
INVxp67_ASAP7_75t_SL g306 ( .A(n_289), .Y(n_306) );
INVxp33_ASAP7_75t_L g307 ( .A(n_193), .Y(n_307) );
BUFx3_ASAP7_75t_L g308 ( .A(n_107), .Y(n_308) );
CKINVDCx16_ASAP7_75t_R g309 ( .A(n_20), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_132), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_272), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_194), .Y(n_312) );
INVxp33_ASAP7_75t_SL g313 ( .A(n_99), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_246), .Y(n_314) );
CKINVDCx20_ASAP7_75t_R g315 ( .A(n_199), .Y(n_315) );
INVxp67_ASAP7_75t_SL g316 ( .A(n_25), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_247), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_42), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_36), .Y(n_319) );
CKINVDCx16_ASAP7_75t_R g320 ( .A(n_80), .Y(n_320) );
INVxp67_ASAP7_75t_SL g321 ( .A(n_222), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_137), .Y(n_322) );
INVxp67_ASAP7_75t_SL g323 ( .A(n_70), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_28), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_291), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_35), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_82), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_17), .Y(n_328) );
CKINVDCx14_ASAP7_75t_R g329 ( .A(n_162), .Y(n_329) );
CKINVDCx20_ASAP7_75t_R g330 ( .A(n_52), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_53), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_261), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_295), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_65), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_293), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_8), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_112), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_174), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_18), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_9), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_270), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_144), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_26), .Y(n_343) );
CKINVDCx20_ASAP7_75t_R g344 ( .A(n_243), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_80), .Y(n_345) );
CKINVDCx20_ASAP7_75t_R g346 ( .A(n_84), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_51), .Y(n_347) );
BUFx3_ASAP7_75t_L g348 ( .A(n_198), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_57), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_12), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_184), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_231), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_71), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_237), .Y(n_354) );
INVxp33_ASAP7_75t_SL g355 ( .A(n_182), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_192), .Y(n_356) );
INVxp67_ASAP7_75t_SL g357 ( .A(n_170), .Y(n_357) );
CKINVDCx20_ASAP7_75t_R g358 ( .A(n_152), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_118), .Y(n_359) );
INVxp33_ASAP7_75t_SL g360 ( .A(n_173), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_73), .Y(n_361) );
INVxp67_ASAP7_75t_SL g362 ( .A(n_101), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_128), .Y(n_363) );
CKINVDCx16_ASAP7_75t_R g364 ( .A(n_191), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_13), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_228), .Y(n_366) );
INVx1_ASAP7_75t_SL g367 ( .A(n_196), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_133), .Y(n_368) );
INVxp67_ASAP7_75t_L g369 ( .A(n_238), .Y(n_369) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_12), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_116), .Y(n_371) );
INVx3_ASAP7_75t_L g372 ( .A(n_103), .Y(n_372) );
BUFx3_ASAP7_75t_L g373 ( .A(n_146), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_236), .Y(n_374) );
INVxp33_ASAP7_75t_SL g375 ( .A(n_29), .Y(n_375) );
INVxp67_ASAP7_75t_SL g376 ( .A(n_176), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_124), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_18), .Y(n_378) );
BUFx5_ASAP7_75t_L g379 ( .A(n_218), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_119), .Y(n_380) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_90), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_47), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_49), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_41), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_298), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_74), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_135), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_102), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_157), .B(n_156), .Y(n_389) );
INVxp67_ASAP7_75t_SL g390 ( .A(n_29), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_2), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_67), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_212), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_105), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_5), .Y(n_395) );
CKINVDCx16_ASAP7_75t_R g396 ( .A(n_19), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_123), .Y(n_397) );
INVxp67_ASAP7_75t_SL g398 ( .A(n_20), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_32), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_39), .Y(n_400) );
CKINVDCx16_ASAP7_75t_R g401 ( .A(n_31), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_296), .Y(n_402) );
CKINVDCx16_ASAP7_75t_R g403 ( .A(n_285), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_83), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_180), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_41), .Y(n_406) );
INVxp67_ASAP7_75t_L g407 ( .A(n_100), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_290), .Y(n_408) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_57), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_226), .Y(n_410) );
CKINVDCx5p33_ASAP7_75t_R g411 ( .A(n_283), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_225), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_276), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_4), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_28), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_210), .Y(n_416) );
INVxp33_ASAP7_75t_L g417 ( .A(n_282), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_110), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_46), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_260), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_227), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_249), .Y(n_422) );
BUFx3_ASAP7_75t_L g423 ( .A(n_19), .Y(n_423) );
INVxp67_ASAP7_75t_L g424 ( .A(n_96), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_26), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_23), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_271), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_148), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_75), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_185), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_109), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_82), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_195), .Y(n_433) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_46), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_83), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_142), .Y(n_436) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_40), .Y(n_437) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_211), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_292), .Y(n_439) );
INVxp33_ASAP7_75t_L g440 ( .A(n_92), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_90), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_172), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_221), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_155), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_65), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_36), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_0), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_181), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_310), .Y(n_449) );
CKINVDCx5p33_ASAP7_75t_R g450 ( .A(n_315), .Y(n_450) );
INVx3_ASAP7_75t_L g451 ( .A(n_372), .Y(n_451) );
BUFx10_ASAP7_75t_L g452 ( .A(n_300), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_344), .Y(n_453) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_345), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_310), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g456 ( .A(n_358), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_436), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_309), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_372), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_320), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_416), .B(n_0), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_364), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_317), .Y(n_463) );
CKINVDCx5p33_ASAP7_75t_R g464 ( .A(n_403), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_317), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_396), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_300), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_332), .Y(n_468) );
CKINVDCx5p33_ASAP7_75t_R g469 ( .A(n_359), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_372), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_440), .B(n_1), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_332), .Y(n_472) );
BUFx2_ASAP7_75t_L g473 ( .A(n_423), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_333), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_333), .Y(n_475) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_308), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_379), .Y(n_477) );
BUFx2_ASAP7_75t_L g478 ( .A(n_423), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_326), .B(n_1), .Y(n_479) );
CKINVDCx5p33_ASAP7_75t_R g480 ( .A(n_359), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_363), .Y(n_481) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_308), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_379), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_473), .B(n_438), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_449), .B(n_304), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_473), .B(n_304), .Y(n_486) );
BUFx3_ASAP7_75t_L g487 ( .A(n_451), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_473), .B(n_312), .Y(n_488) );
INVx3_ASAP7_75t_L g489 ( .A(n_451), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_477), .Y(n_490) );
INVx4_ASAP7_75t_L g491 ( .A(n_451), .Y(n_491) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_476), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_477), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_478), .B(n_451), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_478), .B(n_307), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_478), .B(n_312), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_483), .Y(n_497) );
BUFx3_ASAP7_75t_L g498 ( .A(n_451), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_459), .Y(n_499) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_476), .Y(n_500) );
NAND3xp33_ASAP7_75t_L g501 ( .A(n_449), .B(n_337), .C(n_335), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_479), .B(n_326), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_455), .B(n_417), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_459), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_459), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_455), .B(n_322), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_483), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_477), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_479), .B(n_365), .Y(n_509) );
OAI22xp5_ASAP7_75t_SL g510 ( .A1(n_458), .A2(n_330), .B1(n_346), .B2(n_313), .Y(n_510) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_476), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_463), .B(n_341), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_483), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_470), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_470), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_476), .Y(n_516) );
AND2x4_ASAP7_75t_L g517 ( .A(n_479), .B(n_365), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_467), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_463), .A2(n_318), .B(n_327), .C(n_319), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_470), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_476), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_479), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_479), .Y(n_523) );
AND2x4_ASAP7_75t_L g524 ( .A(n_465), .B(n_384), .Y(n_524) );
INVx3_ASAP7_75t_L g525 ( .A(n_482), .Y(n_525) );
BUFx3_ASAP7_75t_L g526 ( .A(n_476), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_476), .Y(n_527) );
NAND2x1p5_ASAP7_75t_L g528 ( .A(n_465), .B(n_335), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_482), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_450), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_487), .Y(n_531) );
BUFx4f_ASAP7_75t_L g532 ( .A(n_528), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_528), .B(n_452), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_484), .B(n_454), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_487), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_487), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_487), .Y(n_537) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_498), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_528), .B(n_452), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_495), .B(n_452), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_498), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_518), .B(n_471), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_495), .B(n_452), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_503), .B(n_452), .Y(n_544) );
OR2x6_ASAP7_75t_L g545 ( .A(n_510), .B(n_471), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_498), .Y(n_546) );
NOR3xp33_ASAP7_75t_SL g547 ( .A(n_510), .B(n_401), .C(n_453), .Y(n_547) );
BUFx2_ASAP7_75t_L g548 ( .A(n_518), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_484), .B(n_454), .Y(n_549) );
INVxp67_ASAP7_75t_SL g550 ( .A(n_528), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_498), .Y(n_551) );
NOR3xp33_ASAP7_75t_SL g552 ( .A(n_530), .B(n_457), .C(n_456), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_489), .Y(n_553) );
INVxp67_ASAP7_75t_SL g554 ( .A(n_494), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_503), .B(n_494), .Y(n_555) );
INVx4_ASAP7_75t_SL g556 ( .A(n_502), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_486), .B(n_469), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_489), .Y(n_558) );
OR2x6_ASAP7_75t_L g559 ( .A(n_502), .B(n_471), .Y(n_559) );
AND2x4_ASAP7_75t_L g560 ( .A(n_502), .B(n_461), .Y(n_560) );
NOR3xp33_ASAP7_75t_SL g561 ( .A(n_519), .B(n_481), .C(n_480), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_486), .B(n_468), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_502), .B(n_461), .Y(n_563) );
NOR3xp33_ASAP7_75t_SL g564 ( .A(n_519), .B(n_464), .C(n_462), .Y(n_564) );
O2A1O1Ixp33_ASAP7_75t_L g565 ( .A1(n_522), .A2(n_472), .B(n_474), .C(n_468), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_489), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_491), .B(n_472), .Y(n_567) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_491), .Y(n_568) );
INVx6_ASAP7_75t_L g569 ( .A(n_491), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_488), .B(n_474), .Y(n_570) );
INVx2_ASAP7_75t_SL g571 ( .A(n_488), .Y(n_571) );
INVx5_ASAP7_75t_L g572 ( .A(n_491), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_491), .Y(n_573) );
CKINVDCx20_ASAP7_75t_R g574 ( .A(n_496), .Y(n_574) );
AND2x4_ASAP7_75t_L g575 ( .A(n_502), .B(n_381), .Y(n_575) );
INVx5_ASAP7_75t_L g576 ( .A(n_489), .Y(n_576) );
NAND2xp33_ASAP7_75t_SL g577 ( .A(n_522), .B(n_458), .Y(n_577) );
INVx2_ASAP7_75t_SL g578 ( .A(n_496), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_524), .B(n_409), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_512), .B(n_475), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_512), .B(n_475), .Y(n_581) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_492), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_489), .Y(n_583) );
AND2x4_ASAP7_75t_L g584 ( .A(n_509), .B(n_435), .Y(n_584) );
NOR3xp33_ASAP7_75t_SL g585 ( .A(n_501), .B(n_350), .C(n_347), .Y(n_585) );
BUFx10_ASAP7_75t_L g586 ( .A(n_509), .Y(n_586) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_492), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_509), .Y(n_588) );
OAI22xp5_ASAP7_75t_SL g589 ( .A1(n_523), .A2(n_466), .B1(n_460), .B2(n_313), .Y(n_589) );
INVx4_ASAP7_75t_L g590 ( .A(n_509), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_517), .Y(n_591) );
BUFx3_ASAP7_75t_L g592 ( .A(n_517), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_517), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_517), .B(n_363), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_499), .Y(n_595) );
CKINVDCx5p33_ASAP7_75t_R g596 ( .A(n_517), .Y(n_596) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_492), .Y(n_597) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_492), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_524), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_523), .B(n_374), .Y(n_600) );
CKINVDCx16_ASAP7_75t_R g601 ( .A(n_524), .Y(n_601) );
BUFx10_ASAP7_75t_L g602 ( .A(n_524), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_499), .Y(n_603) );
OR2x6_ASAP7_75t_L g604 ( .A(n_506), .B(n_407), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_504), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_504), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_505), .Y(n_607) );
AND2x4_ASAP7_75t_L g608 ( .A(n_485), .B(n_316), .Y(n_608) );
NOR2xp33_ASAP7_75t_R g609 ( .A(n_505), .B(n_466), .Y(n_609) );
BUFx4f_ASAP7_75t_L g610 ( .A(n_514), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_506), .B(n_374), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_485), .B(n_301), .Y(n_612) );
BUFx4f_ASAP7_75t_SL g613 ( .A(n_514), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_515), .B(n_377), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_515), .B(n_377), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_520), .B(n_388), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_520), .B(n_347), .Y(n_617) );
BUFx2_ASAP7_75t_L g618 ( .A(n_501), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_526), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_592), .Y(n_620) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_532), .Y(n_621) );
OAI21xp5_ASAP7_75t_L g622 ( .A1(n_567), .A2(n_497), .B(n_493), .Y(n_622) );
INVxp67_ASAP7_75t_SL g623 ( .A(n_550), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_568), .Y(n_624) );
BUFx5_ASAP7_75t_L g625 ( .A(n_586), .Y(n_625) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_532), .Y(n_626) );
INVx1_ASAP7_75t_SL g627 ( .A(n_548), .Y(n_627) );
A2O1A1Ixp33_ASAP7_75t_L g628 ( .A1(n_565), .A2(n_318), .B(n_327), .C(n_319), .Y(n_628) );
CKINVDCx16_ASAP7_75t_R g629 ( .A(n_609), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_554), .B(n_350), .Y(n_630) );
AOI22xp33_ASAP7_75t_SL g631 ( .A1(n_574), .A2(n_375), .B1(n_399), .B2(n_355), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_568), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g633 ( .A(n_609), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_556), .Y(n_634) );
BUFx3_ASAP7_75t_L g635 ( .A(n_613), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_571), .B(n_375), .Y(n_636) );
BUFx6f_ASAP7_75t_L g637 ( .A(n_568), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_534), .B(n_399), .Y(n_638) );
BUFx6f_ASAP7_75t_L g639 ( .A(n_568), .Y(n_639) );
INVx8_ASAP7_75t_L g640 ( .A(n_572), .Y(n_640) );
INVx3_ASAP7_75t_L g641 ( .A(n_572), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_556), .Y(n_642) );
INVx3_ASAP7_75t_L g643 ( .A(n_572), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_573), .Y(n_644) );
BUFx2_ASAP7_75t_L g645 ( .A(n_550), .Y(n_645) );
BUFx12f_ASAP7_75t_L g646 ( .A(n_545), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_556), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_567), .A2(n_508), .B(n_490), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_554), .A2(n_355), .B1(n_360), .B2(n_301), .Y(n_649) );
INVx2_ASAP7_75t_SL g650 ( .A(n_613), .Y(n_650) );
OAI321xp33_ASAP7_75t_L g651 ( .A1(n_555), .A2(n_424), .A3(n_395), .B1(n_425), .B2(n_426), .C(n_361), .Y(n_651) );
OR2x2_ASAP7_75t_SL g652 ( .A(n_601), .B(n_328), .Y(n_652) );
INVxp67_ASAP7_75t_L g653 ( .A(n_542), .Y(n_653) );
BUFx3_ASAP7_75t_L g654 ( .A(n_572), .Y(n_654) );
O2A1O1Ixp5_ASAP7_75t_L g655 ( .A1(n_543), .A2(n_493), .B(n_507), .C(n_497), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_583), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_586), .Y(n_657) );
INVx3_ASAP7_75t_L g658 ( .A(n_569), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_588), .A2(n_360), .B1(n_328), .B2(n_334), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_595), .Y(n_660) );
INVx1_ASAP7_75t_SL g661 ( .A(n_574), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_602), .Y(n_662) );
BUFx3_ASAP7_75t_L g663 ( .A(n_538), .Y(n_663) );
BUFx4_ASAP7_75t_SL g664 ( .A(n_545), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_602), .Y(n_665) );
INVx5_ASAP7_75t_L g666 ( .A(n_569), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_578), .B(n_493), .Y(n_667) );
BUFx6f_ASAP7_75t_L g668 ( .A(n_538), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_549), .B(n_323), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_542), .B(n_493), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_562), .B(n_497), .Y(n_671) );
AOI21xp5_ASAP7_75t_L g672 ( .A1(n_533), .A2(n_508), .B(n_490), .Y(n_672) );
O2A1O1Ixp33_ASAP7_75t_L g673 ( .A1(n_565), .A2(n_398), .B(n_390), .C(n_353), .Y(n_673) );
BUFx3_ASAP7_75t_L g674 ( .A(n_538), .Y(n_674) );
INVx3_ASAP7_75t_L g675 ( .A(n_569), .Y(n_675) );
O2A1O1Ixp5_ASAP7_75t_L g676 ( .A1(n_543), .A2(n_497), .B(n_513), .C(n_507), .Y(n_676) );
BUFx4f_ASAP7_75t_L g677 ( .A(n_559), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_604), .A2(n_397), .B1(n_411), .B2(n_388), .Y(n_678) );
AND2x4_ASAP7_75t_L g679 ( .A(n_560), .B(n_331), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g680 ( .A1(n_533), .A2(n_508), .B(n_490), .Y(n_680) );
INVx2_ASAP7_75t_L g681 ( .A(n_607), .Y(n_681) );
BUFx6f_ASAP7_75t_L g682 ( .A(n_538), .Y(n_682) );
OAI21x1_ASAP7_75t_L g683 ( .A1(n_539), .A2(n_525), .B(n_513), .Y(n_683) );
BUFx12f_ASAP7_75t_L g684 ( .A(n_545), .Y(n_684) );
INVx3_ASAP7_75t_L g685 ( .A(n_590), .Y(n_685) );
BUFx3_ASAP7_75t_L g686 ( .A(n_610), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_590), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_603), .Y(n_688) );
INVx2_ASAP7_75t_SL g689 ( .A(n_610), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_605), .Y(n_690) );
NAND2xp5_ASAP7_75t_SL g691 ( .A(n_618), .B(n_507), .Y(n_691) );
BUFx6f_ASAP7_75t_L g692 ( .A(n_576), .Y(n_692) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_576), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_559), .A2(n_596), .B1(n_570), .B2(n_604), .Y(n_694) );
BUFx6f_ASAP7_75t_L g695 ( .A(n_576), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_559), .A2(n_329), .B1(n_411), .B2(n_397), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g697 ( .A1(n_539), .A2(n_544), .B(n_540), .Y(n_697) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_604), .A2(n_433), .B1(n_418), .B2(n_507), .Y(n_698) );
INVx2_ASAP7_75t_SL g699 ( .A(n_576), .Y(n_699) );
BUFx2_ASAP7_75t_L g700 ( .A(n_577), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_557), .B(n_305), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_591), .Y(n_702) );
INVx3_ASAP7_75t_L g703 ( .A(n_531), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_593), .Y(n_704) );
OAI21xp33_ASAP7_75t_L g705 ( .A1(n_611), .A2(n_513), .B(n_382), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_599), .A2(n_331), .B1(n_336), .B2(n_334), .Y(n_706) );
AND2x4_ASAP7_75t_L g707 ( .A(n_560), .B(n_336), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_617), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_563), .A2(n_433), .B1(n_418), .B2(n_513), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_575), .B(n_378), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_575), .B(n_383), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_606), .Y(n_712) );
BUFx6f_ASAP7_75t_L g713 ( .A(n_582), .Y(n_713) );
BUFx2_ASAP7_75t_L g714 ( .A(n_577), .Y(n_714) );
AND2x4_ASAP7_75t_L g715 ( .A(n_563), .B(n_339), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_584), .B(n_339), .Y(n_716) );
BUFx2_ASAP7_75t_L g717 ( .A(n_584), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_580), .A2(n_343), .B1(n_349), .B2(n_340), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_581), .B(n_386), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_608), .B(n_391), .Y(n_720) );
INVx2_ASAP7_75t_L g721 ( .A(n_553), .Y(n_721) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_579), .Y(n_722) );
BUFx3_ASAP7_75t_L g723 ( .A(n_541), .Y(n_723) );
INVx3_ASAP7_75t_L g724 ( .A(n_546), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_608), .B(n_392), .Y(n_725) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_594), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_600), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_558), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_566), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_614), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_615), .Y(n_731) );
BUFx3_ASAP7_75t_L g732 ( .A(n_535), .Y(n_732) );
AND2x4_ASAP7_75t_L g733 ( .A(n_564), .B(n_340), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_616), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_619), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_612), .B(n_404), .Y(n_736) );
OAI222xp33_ASAP7_75t_L g737 ( .A1(n_547), .A2(n_447), .B1(n_446), .B2(n_445), .C1(n_400), .C2(n_429), .Y(n_737) );
OR2x2_ASAP7_75t_L g738 ( .A(n_589), .B(n_343), .Y(n_738) );
AND2x4_ASAP7_75t_L g739 ( .A(n_564), .B(n_349), .Y(n_739) );
AOI21x1_ASAP7_75t_SL g740 ( .A1(n_561), .A2(n_526), .B(n_321), .Y(n_740) );
NAND2x1p5_ASAP7_75t_L g741 ( .A(n_536), .B(n_400), .Y(n_741) );
INVx3_ASAP7_75t_L g742 ( .A(n_537), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_612), .B(n_406), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_551), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_582), .A2(n_432), .B1(n_441), .B2(n_429), .Y(n_745) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_561), .A2(n_441), .B1(n_445), .B2(n_432), .Y(n_746) );
AOI222xp33_ASAP7_75t_L g747 ( .A1(n_547), .A2(n_446), .B1(n_447), .B2(n_419), .C1(n_415), .C2(n_414), .Y(n_747) );
CKINVDCx5p33_ASAP7_75t_R g748 ( .A(n_552), .Y(n_748) );
INVx1_ASAP7_75t_SL g749 ( .A(n_582), .Y(n_749) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_627), .A2(n_585), .B1(n_357), .B2(n_362), .Y(n_750) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_645), .Y(n_751) );
OR2x2_ASAP7_75t_L g752 ( .A(n_661), .B(n_384), .Y(n_752) );
AOI221xp5_ASAP7_75t_L g753 ( .A1(n_708), .A2(n_585), .B1(n_370), .B2(n_437), .C(n_434), .Y(n_753) );
AO21x2_ASAP7_75t_L g754 ( .A1(n_697), .A2(n_521), .B(n_516), .Y(n_754) );
INVx3_ASAP7_75t_L g755 ( .A(n_640), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_638), .B(n_324), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_667), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_712), .Y(n_758) );
CKINVDCx16_ASAP7_75t_R g759 ( .A(n_629), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_688), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_679), .A2(n_370), .B1(n_434), .B2(n_324), .Y(n_761) );
NAND2xp33_ASAP7_75t_L g762 ( .A(n_625), .B(n_379), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g763 ( .A1(n_623), .A2(n_369), .B1(n_376), .B2(n_306), .Y(n_763) );
O2A1O1Ixp33_ASAP7_75t_SL g764 ( .A1(n_628), .A2(n_338), .B(n_342), .C(n_337), .Y(n_764) );
INVx4_ASAP7_75t_L g765 ( .A(n_640), .Y(n_765) );
AND2x4_ASAP7_75t_L g766 ( .A(n_621), .B(n_338), .Y(n_766) );
OR2x2_ASAP7_75t_L g767 ( .A(n_722), .B(n_2), .Y(n_767) );
INVx2_ASAP7_75t_L g768 ( .A(n_637), .Y(n_768) );
AND2x4_ASAP7_75t_L g769 ( .A(n_621), .B(n_342), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_630), .B(n_324), .Y(n_770) );
HB1xp67_ASAP7_75t_L g771 ( .A(n_640), .Y(n_771) );
AOI21xp5_ASAP7_75t_L g772 ( .A1(n_672), .A2(n_587), .B(n_582), .Y(n_772) );
NAND2xp33_ASAP7_75t_R g773 ( .A(n_700), .B(n_714), .Y(n_773) );
OAI21x1_ASAP7_75t_L g774 ( .A1(n_683), .A2(n_521), .B(n_516), .Y(n_774) );
NOR2x1_ASAP7_75t_SL g775 ( .A(n_621), .B(n_428), .Y(n_775) );
INVx3_ASAP7_75t_L g776 ( .A(n_640), .Y(n_776) );
OR2x2_ASAP7_75t_L g777 ( .A(n_652), .B(n_3), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_688), .Y(n_778) );
CKINVDCx5p33_ASAP7_75t_R g779 ( .A(n_664), .Y(n_779) );
AND2x2_ASAP7_75t_L g780 ( .A(n_717), .B(n_324), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_679), .A2(n_370), .B1(n_434), .B2(n_324), .Y(n_781) );
CKINVDCx5p33_ASAP7_75t_R g782 ( .A(n_633), .Y(n_782) );
INVx2_ASAP7_75t_L g783 ( .A(n_690), .Y(n_783) );
AOI21x1_ASAP7_75t_L g784 ( .A1(n_683), .A2(n_521), .B(n_516), .Y(n_784) );
CKINVDCx11_ASAP7_75t_R g785 ( .A(n_633), .Y(n_785) );
AOI22xp33_ASAP7_75t_SL g786 ( .A1(n_694), .A2(n_370), .B1(n_437), .B2(n_434), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g787 ( .A(n_646), .Y(n_787) );
AO21x2_ASAP7_75t_L g788 ( .A1(n_691), .A2(n_521), .B(n_516), .Y(n_788) );
INVx2_ASAP7_75t_SL g789 ( .A(n_635), .Y(n_789) );
OAI221xp5_ASAP7_75t_L g790 ( .A1(n_631), .A2(n_428), .B1(n_430), .B2(n_431), .C(n_439), .Y(n_790) );
AND2x4_ASAP7_75t_L g791 ( .A(n_621), .B(n_430), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_677), .A2(n_431), .B1(n_442), .B2(n_439), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_677), .A2(n_442), .B1(n_444), .B2(n_443), .Y(n_793) );
OR2x6_ASAP7_75t_L g794 ( .A(n_626), .B(n_370), .Y(n_794) );
INVx2_ASAP7_75t_SL g795 ( .A(n_677), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_670), .Y(n_796) );
O2A1O1Ixp33_ASAP7_75t_L g797 ( .A1(n_628), .A2(n_444), .B(n_443), .C(n_303), .Y(n_797) );
INVx1_ASAP7_75t_SL g798 ( .A(n_679), .Y(n_798) );
OR2x2_ASAP7_75t_L g799 ( .A(n_669), .B(n_5), .Y(n_799) );
AOI22xp5_ASAP7_75t_L g800 ( .A1(n_636), .A2(n_311), .B1(n_314), .B2(n_302), .Y(n_800) );
AND2x2_ASAP7_75t_L g801 ( .A(n_716), .B(n_434), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_690), .Y(n_802) );
NOR3xp33_ASAP7_75t_SL g803 ( .A(n_748), .B(n_354), .C(n_352), .Y(n_803) );
INVx1_ASAP7_75t_SL g804 ( .A(n_707), .Y(n_804) );
AO31x2_ASAP7_75t_L g805 ( .A1(n_746), .A2(n_529), .A3(n_527), .B(n_325), .Y(n_805) );
BUFx6f_ASAP7_75t_L g806 ( .A(n_713), .Y(n_806) );
BUFx6f_ASAP7_75t_L g807 ( .A(n_713), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_707), .A2(n_437), .B1(n_482), .B2(n_356), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_636), .B(n_437), .Y(n_809) );
INVx2_ASAP7_75t_L g810 ( .A(n_637), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_701), .B(n_437), .Y(n_811) );
AOI221xp5_ASAP7_75t_L g812 ( .A1(n_701), .A2(n_410), .B1(n_366), .B2(n_408), .C(n_368), .Y(n_812) );
AND2x2_ASAP7_75t_L g813 ( .A(n_653), .B(n_6), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_707), .Y(n_814) );
OAI21xp5_ASAP7_75t_L g815 ( .A1(n_655), .A2(n_529), .B(n_527), .Y(n_815) );
A2O1A1Ixp33_ASAP7_75t_L g816 ( .A1(n_730), .A2(n_325), .B(n_351), .C(n_322), .Y(n_816) );
OAI21xp5_ASAP7_75t_L g817 ( .A1(n_676), .A2(n_529), .B(n_527), .Y(n_817) );
AOI21xp5_ASAP7_75t_R g818 ( .A1(n_733), .A2(n_6), .B(n_7), .Y(n_818) );
CKINVDCx6p67_ASAP7_75t_R g819 ( .A(n_684), .Y(n_819) );
AND2x4_ASAP7_75t_L g820 ( .A(n_626), .B(n_371), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_715), .Y(n_821) );
BUFx3_ASAP7_75t_L g822 ( .A(n_654), .Y(n_822) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_671), .A2(n_367), .B1(n_393), .B2(n_385), .Y(n_823) );
HB1xp67_ASAP7_75t_L g824 ( .A(n_626), .Y(n_824) );
INVx2_ASAP7_75t_L g825 ( .A(n_637), .Y(n_825) );
NAND2xp33_ASAP7_75t_SL g826 ( .A(n_626), .B(n_587), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_715), .A2(n_482), .B1(n_402), .B2(n_405), .Y(n_827) );
OAI21x1_ASAP7_75t_L g828 ( .A1(n_680), .A2(n_525), .B(n_380), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_715), .A2(n_482), .B1(n_413), .B2(n_420), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_727), .B(n_726), .Y(n_830) );
OAI221xp5_ASAP7_75t_L g831 ( .A1(n_738), .A2(n_427), .B1(n_448), .B2(n_422), .C(n_421), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_733), .A2(n_482), .B1(n_394), .B2(n_373), .Y(n_832) );
AOI21xp5_ASAP7_75t_SL g833 ( .A1(n_713), .A2(n_373), .B(n_348), .Y(n_833) );
CKINVDCx6p67_ASAP7_75t_R g834 ( .A(n_684), .Y(n_834) );
AO21x2_ASAP7_75t_L g835 ( .A1(n_691), .A2(n_380), .B(n_351), .Y(n_835) );
AOI22xp5_ASAP7_75t_L g836 ( .A1(n_649), .A2(n_412), .B1(n_387), .B2(n_379), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_649), .A2(n_387), .B1(n_412), .B2(n_348), .Y(n_837) );
CKINVDCx11_ASAP7_75t_R g838 ( .A(n_625), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_731), .B(n_7), .Y(n_839) );
NAND2xp33_ASAP7_75t_L g840 ( .A(n_625), .B(n_379), .Y(n_840) );
CKINVDCx5p33_ASAP7_75t_R g841 ( .A(n_748), .Y(n_841) );
OAI21x1_ASAP7_75t_L g842 ( .A1(n_740), .A2(n_525), .B(n_587), .Y(n_842) );
OAI21x1_ASAP7_75t_L g843 ( .A1(n_648), .A2(n_525), .B(n_587), .Y(n_843) );
INVx2_ASAP7_75t_L g844 ( .A(n_624), .Y(n_844) );
OAI22xp5_ASAP7_75t_L g845 ( .A1(n_741), .A2(n_482), .B1(n_598), .B2(n_597), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_702), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_704), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_733), .A2(n_379), .B1(n_526), .B2(n_525), .Y(n_848) );
INVx2_ASAP7_75t_L g849 ( .A(n_624), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_720), .Y(n_850) );
CKINVDCx5p33_ASAP7_75t_R g851 ( .A(n_678), .Y(n_851) );
CKINVDCx6p67_ASAP7_75t_R g852 ( .A(n_686), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_734), .B(n_8), .Y(n_853) );
OR2x6_ASAP7_75t_L g854 ( .A(n_650), .B(n_597), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_725), .Y(n_855) );
AOI211xp5_ASAP7_75t_L g856 ( .A1(n_737), .A2(n_718), .B(n_673), .C(n_696), .Y(n_856) );
A2O1A1Ixp33_ASAP7_75t_L g857 ( .A1(n_705), .A2(n_526), .B(n_389), .C(n_500), .Y(n_857) );
CKINVDCx5p33_ASAP7_75t_R g858 ( .A(n_698), .Y(n_858) );
HB1xp67_ASAP7_75t_L g859 ( .A(n_625), .Y(n_859) );
AND2x4_ASAP7_75t_L g860 ( .A(n_650), .B(n_9), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_739), .A2(n_379), .B1(n_500), .B2(n_492), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_739), .A2(n_379), .B1(n_500), .B2(n_492), .Y(n_862) );
AND2x4_ASAP7_75t_L g863 ( .A(n_689), .B(n_10), .Y(n_863) );
OR2x2_ASAP7_75t_L g864 ( .A(n_710), .B(n_10), .Y(n_864) );
AOI222xp33_ASAP7_75t_L g865 ( .A1(n_711), .A2(n_492), .B1(n_500), .B2(n_511), .C1(n_15), .C2(n_16), .Y(n_865) );
CKINVDCx20_ASAP7_75t_R g866 ( .A(n_686), .Y(n_866) );
O2A1O1Ixp5_ASAP7_75t_L g867 ( .A1(n_739), .A2(n_500), .B(n_511), .C(n_492), .Y(n_867) );
OA21x2_ASAP7_75t_L g868 ( .A1(n_622), .A2(n_511), .B(n_500), .Y(n_868) );
AND2x4_ASAP7_75t_L g869 ( .A(n_689), .B(n_11), .Y(n_869) );
AND2x2_ASAP7_75t_L g870 ( .A(n_659), .B(n_11), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_741), .Y(n_871) );
OAI222xp33_ASAP7_75t_L g872 ( .A1(n_709), .A2(n_13), .B1(n_14), .B2(n_15), .C1(n_16), .C2(n_17), .Y(n_872) );
AND2x2_ASAP7_75t_L g873 ( .A(n_659), .B(n_14), .Y(n_873) );
OR2x2_ASAP7_75t_L g874 ( .A(n_719), .B(n_21), .Y(n_874) );
INVx2_ASAP7_75t_L g875 ( .A(n_632), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_736), .A2(n_511), .B1(n_500), .B2(n_598), .Y(n_876) );
OAI22xp33_ASAP7_75t_SL g877 ( .A1(n_743), .A2(n_21), .B1(n_22), .B2(n_24), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_687), .Y(n_878) );
OAI22xp33_ASAP7_75t_L g879 ( .A1(n_651), .A2(n_500), .B1(n_511), .B2(n_25), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_620), .Y(n_880) );
BUFx2_ASAP7_75t_L g881 ( .A(n_625), .Y(n_881) );
AOI21xp5_ASAP7_75t_L g882 ( .A1(n_713), .A2(n_598), .B(n_597), .Y(n_882) );
AND2x4_ASAP7_75t_L g883 ( .A(n_654), .B(n_22), .Y(n_883) );
NOR2xp33_ASAP7_75t_R g884 ( .A(n_625), .B(n_24), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_744), .Y(n_885) );
AOI22xp5_ASAP7_75t_L g886 ( .A1(n_625), .A2(n_598), .B1(n_597), .B2(n_511), .Y(n_886) );
CKINVDCx5p33_ASAP7_75t_R g887 ( .A(n_706), .Y(n_887) );
OAI221xp5_ASAP7_75t_L g888 ( .A1(n_856), .A2(n_747), .B1(n_706), .B2(n_745), .C(n_657), .Y(n_888) );
OAI22xp5_ASAP7_75t_L g889 ( .A1(n_887), .A2(n_681), .B1(n_660), .B2(n_745), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_830), .Y(n_890) );
AOI21xp5_ASAP7_75t_L g891 ( .A1(n_772), .A2(n_749), .B(n_681), .Y(n_891) );
AOI22xp5_ASAP7_75t_L g892 ( .A1(n_858), .A2(n_665), .B1(n_662), .B2(n_685), .Y(n_892) );
AOI22xp5_ASAP7_75t_L g893 ( .A1(n_851), .A2(n_685), .B1(n_641), .B2(n_643), .Y(n_893) );
AOI221xp5_ASAP7_75t_L g894 ( .A1(n_831), .A2(n_685), .B1(n_728), .B2(n_660), .C(n_642), .Y(n_894) );
OAI22xp33_ASAP7_75t_L g895 ( .A1(n_777), .A2(n_729), .B1(n_721), .B2(n_643), .Y(n_895) );
AND2x2_ASAP7_75t_L g896 ( .A(n_751), .B(n_699), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_758), .Y(n_897) );
OAI21x1_ASAP7_75t_L g898 ( .A1(n_784), .A2(n_742), .B(n_729), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_870), .A2(n_721), .B1(n_732), .B2(n_647), .Y(n_899) );
OA21x2_ASAP7_75t_L g900 ( .A1(n_828), .A2(n_735), .B(n_656), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_873), .A2(n_732), .B1(n_634), .B2(n_742), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_865), .A2(n_742), .B1(n_723), .B2(n_724), .Y(n_902) );
INVx2_ASAP7_75t_L g903 ( .A(n_760), .Y(n_903) );
NOR2x1_ASAP7_75t_SL g904 ( .A(n_765), .B(n_692), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_801), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_860), .A2(n_723), .B1(n_724), .B2(n_703), .Y(n_906) );
OAI22xp33_ASAP7_75t_L g907 ( .A1(n_751), .A2(n_643), .B1(n_641), .B2(n_637), .Y(n_907) );
AOI22xp5_ASAP7_75t_L g908 ( .A1(n_871), .A2(n_641), .B1(n_699), .B2(n_675), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_850), .B(n_644), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_860), .A2(n_874), .B1(n_809), .B2(n_869), .Y(n_910) );
INVx2_ASAP7_75t_L g911 ( .A(n_778), .Y(n_911) );
OAI31xp33_ASAP7_75t_SL g912 ( .A1(n_879), .A2(n_632), .A3(n_656), .B(n_644), .Y(n_912) );
OAI221xp5_ASAP7_75t_L g913 ( .A1(n_800), .A2(n_675), .B1(n_658), .B2(n_703), .C(n_724), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_863), .A2(n_703), .B1(n_735), .B2(n_639), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_863), .A2(n_639), .B1(n_675), .B2(n_658), .Y(n_915) );
AOI22xp33_ASAP7_75t_SL g916 ( .A1(n_884), .A2(n_639), .B1(n_693), .B2(n_692), .Y(n_916) );
INVxp67_ASAP7_75t_L g917 ( .A(n_859), .Y(n_917) );
OR2x2_ASAP7_75t_SL g918 ( .A(n_759), .B(n_692), .Y(n_918) );
BUFx3_ASAP7_75t_L g919 ( .A(n_838), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_869), .A2(n_639), .B1(n_658), .B2(n_692), .Y(n_920) );
INVx2_ASAP7_75t_L g921 ( .A(n_783), .Y(n_921) );
OAI21x1_ASAP7_75t_L g922 ( .A1(n_843), .A2(n_682), .B(n_668), .Y(n_922) );
INVx3_ASAP7_75t_L g923 ( .A(n_838), .Y(n_923) );
OAI221xp5_ASAP7_75t_L g924 ( .A1(n_790), .A2(n_786), .B1(n_812), .B2(n_855), .C(n_767), .Y(n_924) );
INVx2_ASAP7_75t_L g925 ( .A(n_802), .Y(n_925) );
AND2x4_ASAP7_75t_SL g926 ( .A(n_765), .B(n_695), .Y(n_926) );
OAI22xp5_ASAP7_75t_L g927 ( .A1(n_798), .A2(n_666), .B1(n_663), .B2(n_674), .Y(n_927) );
CKINVDCx20_ASAP7_75t_R g928 ( .A(n_779), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_884), .A2(n_695), .B1(n_693), .B2(n_663), .Y(n_929) );
OAI22xp5_ASAP7_75t_L g930 ( .A1(n_804), .A2(n_666), .B1(n_674), .B2(n_682), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_799), .A2(n_695), .B1(n_693), .B2(n_682), .Y(n_931) );
AND2x2_ASAP7_75t_L g932 ( .A(n_757), .B(n_693), .Y(n_932) );
NOR2xp33_ASAP7_75t_L g933 ( .A(n_814), .B(n_666), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_885), .Y(n_934) );
BUFx2_ASAP7_75t_L g935 ( .A(n_866), .Y(n_935) );
AOI221xp5_ASAP7_75t_L g936 ( .A1(n_797), .A2(n_682), .B1(n_668), .B2(n_666), .C(n_511), .Y(n_936) );
OAI21xp5_ASAP7_75t_L g937 ( .A1(n_816), .A2(n_666), .B(n_668), .Y(n_937) );
INVx2_ASAP7_75t_SL g938 ( .A(n_771), .Y(n_938) );
AOI22xp5_ASAP7_75t_L g939 ( .A1(n_883), .A2(n_27), .B1(n_30), .B2(n_31), .Y(n_939) );
AOI222xp33_ASAP7_75t_L g940 ( .A1(n_785), .A2(n_27), .B1(n_30), .B2(n_32), .C1(n_33), .C2(n_34), .Y(n_940) );
OAI211xp5_ASAP7_75t_SL g941 ( .A1(n_803), .A2(n_33), .B(n_34), .C(n_35), .Y(n_941) );
BUFx6f_ASAP7_75t_L g942 ( .A(n_806), .Y(n_942) );
OAI22xp5_ASAP7_75t_L g943 ( .A1(n_786), .A2(n_37), .B1(n_38), .B2(n_39), .Y(n_943) );
OR2x2_ASAP7_75t_L g944 ( .A(n_752), .B(n_37), .Y(n_944) );
BUFx12f_ASAP7_75t_L g945 ( .A(n_785), .Y(n_945) );
OA21x2_ASAP7_75t_L g946 ( .A1(n_857), .A2(n_106), .B(n_104), .Y(n_946) );
AOI21x1_ASAP7_75t_L g947 ( .A1(n_868), .A2(n_111), .B(n_108), .Y(n_947) );
AOI22xp5_ASAP7_75t_L g948 ( .A1(n_883), .A2(n_38), .B1(n_40), .B2(n_42), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_864), .A2(n_821), .B1(n_853), .B2(n_839), .Y(n_949) );
OAI221xp5_ASAP7_75t_L g950 ( .A1(n_750), .A2(n_43), .B1(n_44), .B2(n_45), .C(n_47), .Y(n_950) );
AND2x4_ASAP7_75t_L g951 ( .A(n_771), .B(n_43), .Y(n_951) );
AOI22xp33_ASAP7_75t_SL g952 ( .A1(n_818), .A2(n_44), .B1(n_45), .B2(n_48), .Y(n_952) );
AND2x2_ASAP7_75t_L g953 ( .A(n_795), .B(n_48), .Y(n_953) );
OAI22xp33_ASAP7_75t_L g954 ( .A1(n_879), .A2(n_49), .B1(n_50), .B2(n_51), .Y(n_954) );
OAI22xp33_ASAP7_75t_L g955 ( .A1(n_773), .A2(n_50), .B1(n_52), .B2(n_53), .Y(n_955) );
AND2x2_ASAP7_75t_L g956 ( .A(n_846), .B(n_54), .Y(n_956) );
INVx4_ASAP7_75t_L g957 ( .A(n_852), .Y(n_957) );
INVx2_ASAP7_75t_L g958 ( .A(n_847), .Y(n_958) );
INVx8_ASAP7_75t_L g959 ( .A(n_794), .Y(n_959) );
AOI211xp5_ASAP7_75t_L g960 ( .A1(n_877), .A2(n_55), .B(n_56), .C(n_58), .Y(n_960) );
AOI22xp5_ASAP7_75t_L g961 ( .A1(n_773), .A2(n_55), .B1(n_56), .B2(n_58), .Y(n_961) );
OAI22xp33_ASAP7_75t_L g962 ( .A1(n_794), .A2(n_59), .B1(n_60), .B2(n_61), .Y(n_962) );
NOR2x1_ASAP7_75t_SL g963 ( .A(n_794), .B(n_59), .Y(n_963) );
OAI21x1_ASAP7_75t_L g964 ( .A1(n_774), .A2(n_114), .B(n_113), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_796), .A2(n_60), .B1(n_61), .B2(n_62), .Y(n_965) );
AND2x2_ASAP7_75t_L g966 ( .A(n_803), .B(n_62), .Y(n_966) );
BUFx3_ASAP7_75t_L g967 ( .A(n_755), .Y(n_967) );
AO21x2_ASAP7_75t_L g968 ( .A1(n_857), .A2(n_117), .B(n_115), .Y(n_968) );
BUFx2_ASAP7_75t_L g969 ( .A(n_859), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_756), .Y(n_970) );
OAI211xp5_ASAP7_75t_L g971 ( .A1(n_836), .A2(n_63), .B(n_64), .C(n_66), .Y(n_971) );
OAI22xp33_ASAP7_75t_L g972 ( .A1(n_792), .A2(n_63), .B1(n_64), .B2(n_66), .Y(n_972) );
AND2x2_ASAP7_75t_L g973 ( .A(n_819), .B(n_834), .Y(n_973) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_827), .A2(n_67), .B1(n_68), .B2(n_69), .Y(n_974) );
OAI221xp5_ASAP7_75t_L g975 ( .A1(n_816), .A2(n_68), .B1(n_69), .B2(n_70), .C(n_71), .Y(n_975) );
OAI332xp33_ASAP7_75t_L g976 ( .A1(n_837), .A2(n_72), .A3(n_73), .B1(n_74), .B2(n_75), .B3(n_76), .C1(n_77), .C2(n_78), .Y(n_976) );
AND2x2_ASAP7_75t_L g977 ( .A(n_813), .B(n_72), .Y(n_977) );
BUFx2_ASAP7_75t_L g978 ( .A(n_822), .Y(n_978) );
CKINVDCx5p33_ASAP7_75t_R g979 ( .A(n_787), .Y(n_979) );
AOI21x1_ASAP7_75t_L g980 ( .A1(n_868), .A2(n_121), .B(n_120), .Y(n_980) );
INVx1_ASAP7_75t_L g981 ( .A(n_878), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_753), .A2(n_76), .B1(n_77), .B2(n_78), .Y(n_982) );
AND2x2_ASAP7_75t_L g983 ( .A(n_780), .B(n_79), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_766), .A2(n_79), .B1(n_81), .B2(n_84), .Y(n_984) );
OAI22xp5_ASAP7_75t_L g985 ( .A1(n_827), .A2(n_81), .B1(n_85), .B2(n_86), .Y(n_985) );
OR2x6_ASAP7_75t_L g986 ( .A(n_881), .B(n_85), .Y(n_986) );
AOI21xp33_ASAP7_75t_SL g987 ( .A1(n_841), .A2(n_86), .B(n_87), .Y(n_987) );
OAI22xp5_ASAP7_75t_L g988 ( .A1(n_829), .A2(n_87), .B1(n_88), .B2(n_89), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_766), .A2(n_88), .B1(n_89), .B2(n_91), .Y(n_989) );
OAI22xp5_ASAP7_75t_L g990 ( .A1(n_829), .A2(n_91), .B1(n_92), .B2(n_93), .Y(n_990) );
OAI21x1_ASAP7_75t_L g991 ( .A1(n_882), .A2(n_207), .B(n_297), .Y(n_991) );
AOI22xp5_ASAP7_75t_L g992 ( .A1(n_793), .A2(n_93), .B1(n_94), .B2(n_95), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_769), .A2(n_94), .B1(n_95), .B2(n_96), .Y(n_993) );
AND2x4_ASAP7_75t_L g994 ( .A(n_755), .B(n_97), .Y(n_994) );
INVx1_ASAP7_75t_L g995 ( .A(n_880), .Y(n_995) );
AOI211xp5_ASAP7_75t_L g996 ( .A1(n_872), .A2(n_97), .B(n_98), .C(n_99), .Y(n_996) );
AOI222xp33_ASAP7_75t_L g997 ( .A1(n_872), .A2(n_98), .B1(n_100), .B2(n_122), .C1(n_125), .C2(n_126), .Y(n_997) );
OAI21xp5_ASAP7_75t_SL g998 ( .A1(n_823), .A2(n_127), .B(n_129), .Y(n_998) );
AOI211xp5_ASAP7_75t_L g999 ( .A1(n_763), .A2(n_130), .B(n_131), .C(n_134), .Y(n_999) );
INVx1_ASAP7_75t_SL g1000 ( .A(n_822), .Y(n_1000) );
INVx2_ASAP7_75t_L g1001 ( .A(n_844), .Y(n_1001) );
INVx2_ASAP7_75t_L g1002 ( .A(n_849), .Y(n_1002) );
AOI22xp33_ASAP7_75t_SL g1003 ( .A1(n_775), .A2(n_136), .B1(n_138), .B2(n_139), .Y(n_1003) );
INVx2_ASAP7_75t_L g1004 ( .A(n_875), .Y(n_1004) );
OR2x2_ASAP7_75t_L g1005 ( .A(n_782), .B(n_140), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_811), .Y(n_1006) );
OAI221xp5_ASAP7_75t_L g1007 ( .A1(n_832), .A2(n_141), .B1(n_143), .B2(n_145), .C(n_149), .Y(n_1007) );
OA21x2_ASAP7_75t_L g1008 ( .A1(n_842), .A2(n_150), .B(n_151), .Y(n_1008) );
INVx2_ASAP7_75t_L g1009 ( .A(n_754), .Y(n_1009) );
INVx4_ASAP7_75t_L g1010 ( .A(n_776), .Y(n_1010) );
OAI22xp5_ASAP7_75t_L g1011 ( .A1(n_832), .A2(n_153), .B1(n_158), .B2(n_159), .Y(n_1011) );
AOI21xp33_ASAP7_75t_L g1012 ( .A1(n_770), .A2(n_299), .B(n_161), .Y(n_1012) );
AND2x4_ASAP7_75t_L g1013 ( .A(n_776), .B(n_160), .Y(n_1013) );
INVx2_ASAP7_75t_L g1014 ( .A(n_903), .Y(n_1014) );
OR2x2_ASAP7_75t_L g1015 ( .A(n_890), .B(n_769), .Y(n_1015) );
OAI221xp5_ASAP7_75t_L g1016 ( .A1(n_952), .A2(n_761), .B1(n_781), .B2(n_848), .C(n_862), .Y(n_1016) );
AOI221xp5_ASAP7_75t_L g1017 ( .A1(n_924), .A2(n_764), .B1(n_761), .B2(n_781), .C(n_808), .Y(n_1017) );
NAND2xp5_ASAP7_75t_L g1018 ( .A(n_897), .B(n_791), .Y(n_1018) );
INVx2_ASAP7_75t_L g1019 ( .A(n_903), .Y(n_1019) );
NOR2x2_ASAP7_75t_L g1020 ( .A(n_986), .B(n_854), .Y(n_1020) );
NAND2xp5_ASAP7_75t_L g1021 ( .A(n_934), .B(n_820), .Y(n_1021) );
AND2x2_ASAP7_75t_L g1022 ( .A(n_951), .B(n_789), .Y(n_1022) );
NOR3xp33_ASAP7_75t_L g1023 ( .A(n_976), .B(n_764), .C(n_867), .Y(n_1023) );
OA21x2_ASAP7_75t_L g1024 ( .A1(n_922), .A2(n_867), .B(n_817), .Y(n_1024) );
AOI221xp5_ASAP7_75t_L g1025 ( .A1(n_955), .A2(n_972), .B1(n_888), .B2(n_954), .C(n_895), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_958), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_981), .Y(n_1027) );
INVx2_ASAP7_75t_L g1028 ( .A(n_921), .Y(n_1028) );
CKINVDCx5p33_ASAP7_75t_R g1029 ( .A(n_928), .Y(n_1029) );
INVx8_ASAP7_75t_L g1030 ( .A(n_959), .Y(n_1030) );
OAI221xp5_ASAP7_75t_L g1031 ( .A1(n_952), .A2(n_848), .B1(n_861), .B2(n_862), .C(n_876), .Y(n_1031) );
AOI21xp5_ASAP7_75t_L g1032 ( .A1(n_916), .A2(n_826), .B(n_845), .Y(n_1032) );
OR2x2_ASAP7_75t_L g1033 ( .A(n_944), .B(n_824), .Y(n_1033) );
OR2x2_ASAP7_75t_L g1034 ( .A(n_938), .B(n_824), .Y(n_1034) );
INVx1_ASAP7_75t_L g1035 ( .A(n_995), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_951), .B(n_805), .Y(n_1036) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_956), .B(n_805), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_896), .B(n_805), .Y(n_1038) );
INVx2_ASAP7_75t_L g1039 ( .A(n_921), .Y(n_1039) );
OR2x2_ASAP7_75t_L g1040 ( .A(n_1000), .B(n_805), .Y(n_1040) );
OAI211xp5_ASAP7_75t_SL g1041 ( .A1(n_940), .A2(n_861), .B(n_833), .C(n_762), .Y(n_1041) );
INVxp67_ASAP7_75t_L g1042 ( .A(n_935), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g1043 ( .A1(n_941), .A2(n_835), .B1(n_840), .B2(n_854), .Y(n_1043) );
AOI211xp5_ASAP7_75t_SL g1044 ( .A1(n_962), .A2(n_886), .B(n_825), .C(n_768), .Y(n_1044) );
AO21x2_ASAP7_75t_L g1045 ( .A1(n_937), .A2(n_835), .B(n_815), .Y(n_1045) );
NAND3xp33_ASAP7_75t_L g1046 ( .A(n_960), .B(n_876), .C(n_826), .Y(n_1046) );
OAI21xp5_ASAP7_75t_L g1047 ( .A1(n_902), .A2(n_768), .B(n_825), .Y(n_1047) );
AND2x2_ASAP7_75t_L g1048 ( .A(n_977), .B(n_854), .Y(n_1048) );
CKINVDCx5p33_ASAP7_75t_R g1049 ( .A(n_945), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_909), .Y(n_1050) );
INVx3_ASAP7_75t_L g1051 ( .A(n_926), .Y(n_1051) );
OAI22xp33_ASAP7_75t_L g1052 ( .A1(n_986), .A2(n_810), .B1(n_807), .B2(n_806), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1053 ( .A(n_966), .B(n_810), .Y(n_1053) );
OAI22xp5_ASAP7_75t_SL g1054 ( .A1(n_918), .A2(n_868), .B1(n_807), .B2(n_806), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_986), .B(n_788), .Y(n_1055) );
OA21x2_ASAP7_75t_L g1056 ( .A1(n_1009), .A2(n_788), .B(n_807), .Y(n_1056) );
OA21x2_ASAP7_75t_L g1057 ( .A1(n_898), .A2(n_807), .B(n_806), .Y(n_1057) );
INVx2_ASAP7_75t_L g1058 ( .A(n_900), .Y(n_1058) );
OAI211xp5_ASAP7_75t_SL g1059 ( .A1(n_892), .A2(n_163), .B(n_164), .C(n_165), .Y(n_1059) );
INVx1_ASAP7_75t_L g1060 ( .A(n_911), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_925), .Y(n_1061) );
NOR5xp2_ASAP7_75t_SL g1062 ( .A(n_943), .B(n_166), .C(n_167), .D(n_168), .E(n_169), .Y(n_1062) );
OAI22xp5_ASAP7_75t_L g1063 ( .A1(n_910), .A2(n_171), .B1(n_175), .B2(n_177), .Y(n_1063) );
OAI22xp33_ASAP7_75t_L g1064 ( .A1(n_961), .A2(n_178), .B1(n_179), .B2(n_183), .Y(n_1064) );
OR2x2_ASAP7_75t_L g1065 ( .A(n_978), .B(n_294), .Y(n_1065) );
AOI22xp5_ASAP7_75t_L g1066 ( .A1(n_895), .A2(n_186), .B1(n_187), .B2(n_188), .Y(n_1066) );
AOI33xp33_ASAP7_75t_L g1067 ( .A1(n_972), .A2(n_288), .A3(n_190), .B1(n_197), .B2(n_200), .B3(n_201), .Y(n_1067) );
OR2x6_ASAP7_75t_L g1068 ( .A(n_959), .B(n_189), .Y(n_1068) );
BUFx6f_ASAP7_75t_L g1069 ( .A(n_942), .Y(n_1069) );
HB1xp67_ASAP7_75t_L g1070 ( .A(n_969), .Y(n_1070) );
NAND2xp33_ASAP7_75t_SL g1071 ( .A(n_929), .B(n_910), .Y(n_1071) );
OAI221xp5_ASAP7_75t_SL g1072 ( .A1(n_996), .A2(n_202), .B1(n_203), .B2(n_204), .C(n_205), .Y(n_1072) );
OAI211xp5_ASAP7_75t_L g1073 ( .A1(n_987), .A2(n_206), .B(n_208), .C(n_209), .Y(n_1073) );
NAND3xp33_ASAP7_75t_L g1074 ( .A(n_997), .B(n_214), .C(n_215), .Y(n_1074) );
INVxp67_ASAP7_75t_SL g1075 ( .A(n_916), .Y(n_1075) );
INVxp33_ASAP7_75t_L g1076 ( .A(n_904), .Y(n_1076) );
BUFx6f_ASAP7_75t_L g1077 ( .A(n_942), .Y(n_1077) );
BUFx2_ASAP7_75t_L g1078 ( .A(n_919), .Y(n_1078) );
OAI22xp5_ASAP7_75t_SL g1079 ( .A1(n_957), .A2(n_216), .B1(n_217), .B2(n_219), .Y(n_1079) );
OAI21xp5_ASAP7_75t_L g1080 ( .A1(n_902), .A2(n_220), .B(n_223), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_975), .A2(n_224), .B1(n_229), .B2(n_230), .Y(n_1081) );
NAND2xp5_ASAP7_75t_L g1082 ( .A(n_949), .B(n_232), .Y(n_1082) );
OAI31xp33_ASAP7_75t_L g1083 ( .A1(n_962), .A2(n_234), .A3(n_235), .B(n_240), .Y(n_1083) );
OAI21x1_ASAP7_75t_L g1084 ( .A1(n_947), .A2(n_241), .B(n_242), .Y(n_1084) );
OAI211xp5_ASAP7_75t_L g1085 ( .A1(n_939), .A2(n_244), .B(n_245), .C(n_248), .Y(n_1085) );
BUFx2_ASAP7_75t_L g1086 ( .A(n_919), .Y(n_1086) );
AND2x2_ASAP7_75t_L g1087 ( .A(n_932), .B(n_250), .Y(n_1087) );
INVxp67_ASAP7_75t_L g1088 ( .A(n_994), .Y(n_1088) );
HB1xp67_ASAP7_75t_L g1089 ( .A(n_917), .Y(n_1089) );
OAI211xp5_ASAP7_75t_L g1090 ( .A1(n_948), .A2(n_251), .B(n_252), .C(n_253), .Y(n_1090) );
OAI22xp5_ASAP7_75t_L g1091 ( .A1(n_906), .A2(n_254), .B1(n_255), .B2(n_256), .Y(n_1091) );
NAND2xp5_ASAP7_75t_L g1092 ( .A(n_949), .B(n_257), .Y(n_1092) );
OAI31xp33_ASAP7_75t_L g1093 ( .A1(n_954), .A2(n_258), .A3(n_259), .B(n_262), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_950), .A2(n_263), .B1(n_264), .B2(n_265), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_994), .Y(n_1095) );
AND2x4_ASAP7_75t_L g1096 ( .A(n_923), .B(n_266), .Y(n_1096) );
AOI21xp5_ASAP7_75t_L g1097 ( .A1(n_907), .A2(n_267), .B(n_268), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_974), .A2(n_269), .B1(n_273), .B2(n_274), .Y(n_1098) );
AOI221xp5_ASAP7_75t_L g1099 ( .A1(n_985), .A2(n_275), .B1(n_277), .B2(n_278), .C(n_279), .Y(n_1099) );
INVx2_ASAP7_75t_L g1100 ( .A(n_900), .Y(n_1100) );
INVxp67_ASAP7_75t_SL g1101 ( .A(n_917), .Y(n_1101) );
HB1xp67_ASAP7_75t_L g1102 ( .A(n_907), .Y(n_1102) );
AOI221xp5_ASAP7_75t_L g1103 ( .A1(n_988), .A2(n_280), .B1(n_281), .B2(n_284), .C(n_286), .Y(n_1103) );
OAI31xp33_ASAP7_75t_L g1104 ( .A1(n_971), .A2(n_287), .A3(n_990), .B(n_998), .Y(n_1104) );
NAND4xp25_ASAP7_75t_L g1105 ( .A(n_984), .B(n_989), .C(n_993), .D(n_965), .Y(n_1105) );
BUFx10_ASAP7_75t_L g1106 ( .A(n_926), .Y(n_1106) );
INVx3_ASAP7_75t_L g1107 ( .A(n_959), .Y(n_1107) );
OAI221xp5_ASAP7_75t_SL g1108 ( .A1(n_984), .A2(n_989), .B1(n_993), .B2(n_992), .C(n_965), .Y(n_1108) );
BUFx3_ASAP7_75t_L g1109 ( .A(n_923), .Y(n_1109) );
OAI21xp5_ASAP7_75t_L g1110 ( .A1(n_982), .A2(n_889), .B(n_899), .Y(n_1110) );
BUFx2_ASAP7_75t_L g1111 ( .A(n_957), .Y(n_1111) );
AND2x4_ASAP7_75t_L g1112 ( .A(n_1010), .B(n_1013), .Y(n_1112) );
INVx2_ASAP7_75t_L g1113 ( .A(n_900), .Y(n_1113) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_1038), .B(n_1002), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_1037), .B(n_1001), .Y(n_1115) );
AOI211xp5_ASAP7_75t_L g1116 ( .A1(n_1108), .A2(n_1005), .B(n_953), .C(n_973), .Y(n_1116) );
OAI21xp5_ASAP7_75t_L g1117 ( .A1(n_1046), .A2(n_999), .B(n_914), .Y(n_1117) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1058), .Y(n_1118) );
AND2x4_ASAP7_75t_SL g1119 ( .A(n_1106), .B(n_1010), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_1014), .B(n_1004), .Y(n_1120) );
INVx1_ASAP7_75t_SL g1121 ( .A(n_1111), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1058), .Y(n_1122) );
INVx2_ASAP7_75t_L g1123 ( .A(n_1100), .Y(n_1123) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1100), .Y(n_1124) );
BUFx2_ASAP7_75t_L g1125 ( .A(n_1020), .Y(n_1125) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1113), .Y(n_1126) );
OAI22xp5_ASAP7_75t_L g1127 ( .A1(n_1068), .A2(n_929), .B1(n_914), .B2(n_920), .Y(n_1127) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1113), .Y(n_1128) );
OR2x2_ASAP7_75t_L g1129 ( .A(n_1070), .B(n_931), .Y(n_1129) );
OAI31xp33_ASAP7_75t_L g1130 ( .A1(n_1071), .A2(n_1013), .A3(n_1007), .B(n_933), .Y(n_1130) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1019), .Y(n_1131) );
INVx2_ASAP7_75t_SL g1132 ( .A(n_1106), .Y(n_1132) );
OR2x2_ASAP7_75t_L g1133 ( .A(n_1089), .B(n_920), .Y(n_1133) );
BUFx2_ASAP7_75t_L g1134 ( .A(n_1020), .Y(n_1134) );
INVx2_ASAP7_75t_L g1135 ( .A(n_1019), .Y(n_1135) );
AOI33xp33_ASAP7_75t_L g1136 ( .A1(n_1027), .A2(n_901), .A3(n_905), .B1(n_1003), .B2(n_915), .B3(n_893), .Y(n_1136) );
INVx2_ASAP7_75t_L g1137 ( .A(n_1028), .Y(n_1137) );
HB1xp67_ASAP7_75t_L g1138 ( .A(n_1089), .Y(n_1138) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1039), .Y(n_1139) );
NAND2xp5_ASAP7_75t_L g1140 ( .A(n_1050), .B(n_983), .Y(n_1140) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1035), .Y(n_1141) );
NAND2xp5_ASAP7_75t_SL g1142 ( .A(n_1112), .B(n_912), .Y(n_1142) );
INVxp67_ASAP7_75t_L g1143 ( .A(n_1078), .Y(n_1143) );
AND2x4_ASAP7_75t_L g1144 ( .A(n_1036), .B(n_963), .Y(n_1144) );
AOI22xp5_ASAP7_75t_L g1145 ( .A1(n_1105), .A2(n_894), .B1(n_933), .B2(n_915), .Y(n_1145) );
BUFx2_ASAP7_75t_L g1146 ( .A(n_1054), .Y(n_1146) );
HB1xp67_ASAP7_75t_L g1147 ( .A(n_1101), .Y(n_1147) );
NAND2xp5_ASAP7_75t_L g1148 ( .A(n_1026), .B(n_908), .Y(n_1148) );
INVx2_ASAP7_75t_L g1149 ( .A(n_1056), .Y(n_1149) );
OAI33xp33_ASAP7_75t_L g1150 ( .A1(n_1042), .A2(n_1011), .A3(n_970), .B1(n_1006), .B2(n_927), .B3(n_979), .Y(n_1150) );
OAI221xp5_ASAP7_75t_L g1151 ( .A1(n_1025), .A2(n_913), .B1(n_967), .B2(n_936), .C(n_946), .Y(n_1151) );
OAI33xp33_ASAP7_75t_L g1152 ( .A1(n_1064), .A2(n_930), .A3(n_968), .B1(n_946), .B2(n_967), .B3(n_980), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_1060), .B(n_946), .Y(n_1153) );
NAND2xp5_ASAP7_75t_L g1154 ( .A(n_1061), .B(n_891), .Y(n_1154) );
INVx1_ASAP7_75t_SL g1155 ( .A(n_1106), .Y(n_1155) );
OAI221xp5_ASAP7_75t_L g1156 ( .A1(n_1088), .A2(n_1012), .B1(n_1008), .B2(n_942), .C(n_991), .Y(n_1156) );
BUFx2_ASAP7_75t_L g1157 ( .A(n_1112), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1040), .Y(n_1158) );
OAI33xp33_ASAP7_75t_L g1159 ( .A1(n_1064), .A2(n_942), .A3(n_964), .B1(n_1008), .B2(n_1021), .B3(n_1095), .Y(n_1159) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1056), .Y(n_1160) );
CKINVDCx16_ASAP7_75t_R g1161 ( .A(n_1068), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1055), .B(n_1008), .Y(n_1162) );
INVx2_ASAP7_75t_L g1163 ( .A(n_1056), .Y(n_1163) );
OR2x2_ASAP7_75t_L g1164 ( .A(n_1033), .B(n_1015), .Y(n_1164) );
AND3x2_ASAP7_75t_L g1165 ( .A(n_1086), .B(n_1112), .C(n_1096), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1053), .B(n_1110), .Y(n_1166) );
INVx6_ASAP7_75t_L g1167 ( .A(n_1030), .Y(n_1167) );
NAND2xp5_ASAP7_75t_L g1168 ( .A(n_1018), .B(n_1022), .Y(n_1168) );
INVx1_ASAP7_75t_SL g1169 ( .A(n_1029), .Y(n_1169) );
OAI33xp33_ASAP7_75t_L g1170 ( .A1(n_1049), .A2(n_1079), .A3(n_1052), .B1(n_1092), .B2(n_1082), .B3(n_1034), .Y(n_1170) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1057), .Y(n_1171) );
AOI221xp5_ASAP7_75t_L g1172 ( .A1(n_1071), .A2(n_1023), .B1(n_1017), .B2(n_1075), .C(n_1072), .Y(n_1172) );
OAI31xp33_ASAP7_75t_L g1173 ( .A1(n_1052), .A2(n_1041), .A3(n_1044), .B(n_1074), .Y(n_1173) );
NOR2xp33_ASAP7_75t_L g1174 ( .A(n_1029), .B(n_1107), .Y(n_1174) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1109), .Y(n_1175) );
INVx2_ASAP7_75t_L g1176 ( .A(n_1057), .Y(n_1176) );
AND2x4_ASAP7_75t_L g1177 ( .A(n_1096), .B(n_1069), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1102), .B(n_1047), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1102), .B(n_1045), .Y(n_1179) );
OR2x2_ASAP7_75t_L g1180 ( .A(n_1068), .B(n_1076), .Y(n_1180) );
NAND2xp5_ASAP7_75t_L g1181 ( .A(n_1048), .B(n_1107), .Y(n_1181) );
OAI211xp5_ASAP7_75t_L g1182 ( .A1(n_1104), .A2(n_1083), .B(n_1030), .C(n_1080), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1045), .B(n_1087), .Y(n_1183) );
HB1xp67_ASAP7_75t_L g1184 ( .A(n_1076), .Y(n_1184) );
AOI21xp33_ASAP7_75t_L g1185 ( .A1(n_1016), .A2(n_1043), .B(n_1073), .Y(n_1185) );
INVx2_ASAP7_75t_L g1186 ( .A(n_1057), .Y(n_1186) );
INVx1_ASAP7_75t_SL g1187 ( .A(n_1030), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1024), .Y(n_1188) );
INVx2_ASAP7_75t_L g1189 ( .A(n_1123), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1115), .B(n_1024), .Y(n_1190) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1166), .B(n_1051), .Y(n_1191) );
HB1xp67_ASAP7_75t_L g1192 ( .A(n_1147), .Y(n_1192) );
OR2x2_ASAP7_75t_L g1193 ( .A(n_1158), .B(n_1065), .Y(n_1193) );
AOI21xp5_ASAP7_75t_L g1194 ( .A1(n_1159), .A2(n_1032), .B(n_1097), .Y(n_1194) );
INVx2_ASAP7_75t_L g1195 ( .A(n_1123), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1115), .B(n_1024), .Y(n_1196) );
INVx1_ASAP7_75t_SL g1197 ( .A(n_1121), .Y(n_1197) );
OR2x2_ASAP7_75t_L g1198 ( .A(n_1158), .B(n_1051), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1199 ( .A(n_1114), .B(n_1069), .Y(n_1199) );
NAND2xp5_ASAP7_75t_L g1200 ( .A(n_1166), .B(n_1096), .Y(n_1200) );
INVx2_ASAP7_75t_L g1201 ( .A(n_1118), .Y(n_1201) );
NAND2xp33_ASAP7_75t_R g1202 ( .A(n_1125), .B(n_1049), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1114), .B(n_1069), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1204 ( .A(n_1178), .B(n_1069), .Y(n_1204) );
AND2x4_ASAP7_75t_L g1205 ( .A(n_1125), .B(n_1077), .Y(n_1205) );
NAND2xp33_ASAP7_75t_SL g1206 ( .A(n_1134), .B(n_1067), .Y(n_1206) );
INVx2_ASAP7_75t_L g1207 ( .A(n_1118), .Y(n_1207) );
INVx2_ASAP7_75t_L g1208 ( .A(n_1122), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1131), .Y(n_1209) );
NAND2xp5_ASAP7_75t_L g1210 ( .A(n_1141), .B(n_1043), .Y(n_1210) );
OR2x2_ASAP7_75t_L g1211 ( .A(n_1138), .B(n_1077), .Y(n_1211) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1164), .Y(n_1212) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1131), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1139), .Y(n_1214) );
NAND2x1p5_ASAP7_75t_L g1215 ( .A(n_1180), .B(n_1077), .Y(n_1215) );
NOR2xp33_ASAP7_75t_R g1216 ( .A(n_1161), .B(n_1077), .Y(n_1216) );
OR2x2_ASAP7_75t_L g1217 ( .A(n_1164), .B(n_1093), .Y(n_1217) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1139), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1219 ( .A(n_1168), .B(n_1094), .Y(n_1219) );
INVx2_ASAP7_75t_L g1220 ( .A(n_1122), .Y(n_1220) );
NAND2xp5_ASAP7_75t_L g1221 ( .A(n_1140), .B(n_1081), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1178), .B(n_1066), .Y(n_1222) );
BUFx12f_ASAP7_75t_L g1223 ( .A(n_1167), .Y(n_1223) );
OR2x2_ASAP7_75t_L g1224 ( .A(n_1129), .B(n_1031), .Y(n_1224) );
AOI21xp33_ASAP7_75t_L g1225 ( .A1(n_1116), .A2(n_1090), .B(n_1085), .Y(n_1225) );
OR2x2_ASAP7_75t_L g1226 ( .A(n_1129), .B(n_1063), .Y(n_1226) );
INVx2_ASAP7_75t_L g1227 ( .A(n_1124), .Y(n_1227) );
NAND2xp5_ASAP7_75t_L g1228 ( .A(n_1120), .B(n_1098), .Y(n_1228) );
NAND4xp25_ASAP7_75t_L g1229 ( .A(n_1172), .B(n_1098), .C(n_1099), .D(n_1103), .Y(n_1229) );
AND2x4_ASAP7_75t_SL g1230 ( .A(n_1132), .B(n_1062), .Y(n_1230) );
NAND2xp5_ASAP7_75t_L g1231 ( .A(n_1120), .B(n_1091), .Y(n_1231) );
NAND2xp33_ASAP7_75t_L g1232 ( .A(n_1180), .B(n_1062), .Y(n_1232) );
INVx1_ASAP7_75t_SL g1233 ( .A(n_1187), .Y(n_1233) );
NAND2xp33_ASAP7_75t_SL g1234 ( .A(n_1134), .B(n_1059), .Y(n_1234) );
INVx2_ASAP7_75t_L g1235 ( .A(n_1124), .Y(n_1235) );
NAND2xp5_ASAP7_75t_L g1236 ( .A(n_1143), .B(n_1084), .Y(n_1236) );
CKINVDCx5p33_ASAP7_75t_R g1237 ( .A(n_1167), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1238 ( .A(n_1175), .B(n_1084), .Y(n_1238) );
NAND2xp5_ASAP7_75t_L g1239 ( .A(n_1181), .B(n_1184), .Y(n_1239) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1133), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1126), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1179), .B(n_1128), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1133), .Y(n_1243) );
NOR4xp25_ASAP7_75t_SL g1244 ( .A(n_1146), .B(n_1185), .C(n_1142), .D(n_1151), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_1179), .B(n_1126), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1128), .B(n_1162), .Y(n_1246) );
XNOR2xp5_ASAP7_75t_L g1247 ( .A(n_1169), .B(n_1165), .Y(n_1247) );
INVx2_ASAP7_75t_L g1248 ( .A(n_1201), .Y(n_1248) );
AOI21xp5_ASAP7_75t_L g1249 ( .A1(n_1206), .A2(n_1170), .B(n_1152), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1250 ( .A(n_1246), .B(n_1162), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g1251 ( .A(n_1192), .B(n_1157), .Y(n_1251) );
AOI22xp33_ASAP7_75t_L g1252 ( .A1(n_1206), .A2(n_1150), .B1(n_1173), .B2(n_1145), .Y(n_1252) );
NAND2xp5_ASAP7_75t_L g1253 ( .A(n_1212), .B(n_1157), .Y(n_1253) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1199), .B(n_1144), .Y(n_1254) );
AND2x4_ASAP7_75t_L g1255 ( .A(n_1242), .B(n_1245), .Y(n_1255) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1224), .B(n_1144), .Y(n_1256) );
AOI22xp5_ASAP7_75t_L g1257 ( .A1(n_1221), .A2(n_1182), .B1(n_1144), .B2(n_1127), .Y(n_1257) );
NOR2x1_ASAP7_75t_SL g1258 ( .A(n_1223), .B(n_1132), .Y(n_1258) );
A2O1A1Ixp33_ASAP7_75t_L g1259 ( .A1(n_1225), .A2(n_1119), .B(n_1130), .C(n_1136), .Y(n_1259) );
OAI22xp5_ASAP7_75t_L g1260 ( .A1(n_1247), .A2(n_1167), .B1(n_1155), .B2(n_1119), .Y(n_1260) );
INVx1_ASAP7_75t_SL g1261 ( .A(n_1233), .Y(n_1261) );
AOI21xp33_ASAP7_75t_L g1262 ( .A1(n_1224), .A2(n_1232), .B(n_1210), .Y(n_1262) );
NAND2xp5_ASAP7_75t_L g1263 ( .A(n_1240), .B(n_1243), .Y(n_1263) );
OAI22xp5_ASAP7_75t_L g1264 ( .A1(n_1247), .A2(n_1167), .B1(n_1117), .B2(n_1177), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1199), .B(n_1183), .Y(n_1265) );
NOR2xp33_ASAP7_75t_L g1266 ( .A(n_1197), .B(n_1148), .Y(n_1266) );
NAND2x1_ASAP7_75t_L g1267 ( .A(n_1205), .B(n_1177), .Y(n_1267) );
AOI21xp33_ASAP7_75t_SL g1268 ( .A1(n_1202), .A2(n_1174), .B(n_1177), .Y(n_1268) );
INVx2_ASAP7_75t_SL g1269 ( .A(n_1216), .Y(n_1269) );
OAI22xp33_ASAP7_75t_L g1270 ( .A1(n_1200), .A2(n_1156), .B1(n_1135), .B2(n_1137), .Y(n_1270) );
NOR4xp25_ASAP7_75t_SL g1271 ( .A(n_1237), .B(n_1160), .C(n_1171), .D(n_1188), .Y(n_1271) );
CKINVDCx16_ASAP7_75t_R g1272 ( .A(n_1223), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_1203), .B(n_1183), .Y(n_1273) );
OAI32xp33_ASAP7_75t_L g1274 ( .A1(n_1237), .A2(n_1160), .A3(n_1171), .B1(n_1163), .B2(n_1149), .Y(n_1274) );
AOI21xp5_ASAP7_75t_L g1275 ( .A1(n_1232), .A2(n_1163), .B(n_1149), .Y(n_1275) );
NOR2xp33_ASAP7_75t_L g1276 ( .A(n_1239), .B(n_1154), .Y(n_1276) );
INVx2_ASAP7_75t_SL g1277 ( .A(n_1211), .Y(n_1277) );
OAI21x1_ASAP7_75t_SL g1278 ( .A1(n_1191), .A2(n_1135), .B(n_1137), .Y(n_1278) );
AOI21xp5_ASAP7_75t_L g1279 ( .A1(n_1234), .A2(n_1176), .B(n_1186), .Y(n_1279) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1209), .Y(n_1280) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1209), .Y(n_1281) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1213), .Y(n_1282) );
NOR2xp33_ASAP7_75t_L g1283 ( .A(n_1217), .B(n_1153), .Y(n_1283) );
INVx2_ASAP7_75t_L g1284 ( .A(n_1201), .Y(n_1284) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1213), .Y(n_1285) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1214), .Y(n_1286) );
INVx3_ASAP7_75t_SL g1287 ( .A(n_1272), .Y(n_1287) );
AOI21xp5_ASAP7_75t_L g1288 ( .A1(n_1249), .A2(n_1234), .B(n_1230), .Y(n_1288) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1248), .Y(n_1289) );
OR2x2_ASAP7_75t_L g1290 ( .A(n_1255), .B(n_1245), .Y(n_1290) );
NAND2xp5_ASAP7_75t_L g1291 ( .A(n_1276), .B(n_1242), .Y(n_1291) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1248), .Y(n_1292) );
NOR2xp33_ASAP7_75t_L g1293 ( .A(n_1261), .B(n_1193), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1255), .B(n_1246), .Y(n_1294) );
NOR2x1_ASAP7_75t_L g1295 ( .A(n_1260), .B(n_1211), .Y(n_1295) );
AOI31xp33_ASAP7_75t_L g1296 ( .A1(n_1268), .A2(n_1217), .A3(n_1193), .B(n_1226), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g1297 ( .A(n_1276), .B(n_1196), .Y(n_1297) );
NOR3xp33_ASAP7_75t_SL g1298 ( .A(n_1264), .B(n_1229), .C(n_1219), .Y(n_1298) );
OR2x2_ASAP7_75t_L g1299 ( .A(n_1255), .B(n_1196), .Y(n_1299) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1284), .Y(n_1300) );
NOR3xp33_ASAP7_75t_SL g1301 ( .A(n_1259), .B(n_1194), .C(n_1244), .Y(n_1301) );
OAI211xp5_ASAP7_75t_L g1302 ( .A1(n_1252), .A2(n_1226), .B(n_1222), .C(n_1198), .Y(n_1302) );
AOI322xp5_ASAP7_75t_L g1303 ( .A1(n_1252), .A2(n_1222), .A3(n_1190), .B1(n_1204), .B2(n_1228), .C1(n_1241), .C2(n_1203), .Y(n_1303) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1284), .Y(n_1304) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1250), .B(n_1190), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1250), .B(n_1204), .Y(n_1306) );
INVx2_ASAP7_75t_L g1307 ( .A(n_1280), .Y(n_1307) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1281), .Y(n_1308) );
AOI211xp5_ASAP7_75t_L g1309 ( .A1(n_1262), .A2(n_1259), .B(n_1274), .C(n_1270), .Y(n_1309) );
NOR2xp33_ASAP7_75t_L g1310 ( .A(n_1266), .B(n_1198), .Y(n_1310) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1282), .Y(n_1311) );
AOI22xp5_ASAP7_75t_L g1312 ( .A1(n_1302), .A2(n_1257), .B1(n_1283), .B2(n_1256), .Y(n_1312) );
A2O1A1Ixp33_ASAP7_75t_L g1313 ( .A1(n_1288), .A2(n_1269), .B(n_1279), .C(n_1230), .Y(n_1313) );
XOR2x2_ASAP7_75t_L g1314 ( .A(n_1287), .B(n_1258), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1305), .B(n_1265), .Y(n_1315) );
A2O1A1Ixp33_ASAP7_75t_L g1316 ( .A1(n_1309), .A2(n_1283), .B(n_1267), .C(n_1251), .Y(n_1316) );
BUFx2_ASAP7_75t_L g1317 ( .A(n_1287), .Y(n_1317) );
OAI211xp5_ASAP7_75t_L g1318 ( .A1(n_1298), .A2(n_1271), .B(n_1253), .C(n_1263), .Y(n_1318) );
OAI22xp5_ASAP7_75t_L g1319 ( .A1(n_1296), .A2(n_1270), .B1(n_1277), .B2(n_1275), .Y(n_1319) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1308), .Y(n_1320) );
AOI21xp33_ASAP7_75t_L g1321 ( .A1(n_1295), .A2(n_1236), .B(n_1278), .Y(n_1321) );
NOR3xp33_ASAP7_75t_L g1322 ( .A(n_1293), .B(n_1238), .C(n_1285), .Y(n_1322) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1308), .Y(n_1323) );
AO22x2_ASAP7_75t_L g1324 ( .A1(n_1311), .A2(n_1286), .B1(n_1214), .B2(n_1218), .Y(n_1324) );
XOR2xp5_ASAP7_75t_L g1325 ( .A(n_1297), .B(n_1254), .Y(n_1325) );
AOI221xp5_ASAP7_75t_L g1326 ( .A1(n_1310), .A2(n_1273), .B1(n_1231), .B2(n_1235), .C(n_1227), .Y(n_1326) );
NOR2x1p5_ASAP7_75t_L g1327 ( .A(n_1314), .B(n_1290), .Y(n_1327) );
OAI21xp33_ASAP7_75t_L g1328 ( .A1(n_1316), .A2(n_1301), .B(n_1303), .Y(n_1328) );
A2O1A1Ixp33_ASAP7_75t_L g1329 ( .A1(n_1317), .A2(n_1290), .B(n_1294), .C(n_1291), .Y(n_1329) );
AOI22xp5_ASAP7_75t_L g1330 ( .A1(n_1312), .A2(n_1294), .B1(n_1305), .B2(n_1306), .Y(n_1330) );
NOR2xp33_ASAP7_75t_R g1331 ( .A(n_1313), .B(n_1205), .Y(n_1331) );
NAND2xp5_ASAP7_75t_L g1332 ( .A(n_1322), .B(n_1306), .Y(n_1332) );
INVx2_ASAP7_75t_L g1333 ( .A(n_1324), .Y(n_1333) );
XOR2xp5_ASAP7_75t_L g1334 ( .A(n_1319), .B(n_1299), .Y(n_1334) );
NAND2xp5_ASAP7_75t_L g1335 ( .A(n_1326), .B(n_1311), .Y(n_1335) );
OAI21xp33_ASAP7_75t_SL g1336 ( .A1(n_1321), .A2(n_1307), .B(n_1304), .Y(n_1336) );
CKINVDCx20_ASAP7_75t_R g1337 ( .A(n_1325), .Y(n_1337) );
AOI22x1_ASAP7_75t_L g1338 ( .A1(n_1324), .A2(n_1215), .B1(n_1300), .B2(n_1292), .Y(n_1338) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1324), .Y(n_1339) );
HB1xp67_ASAP7_75t_L g1340 ( .A(n_1320), .Y(n_1340) );
NOR3xp33_ASAP7_75t_SL g1341 ( .A(n_1319), .B(n_1304), .C(n_1292), .Y(n_1341) );
NOR3x1_ASAP7_75t_L g1342 ( .A(n_1318), .B(n_1289), .C(n_1188), .Y(n_1342) );
A2O1A1Ixp33_ASAP7_75t_L g1343 ( .A1(n_1321), .A2(n_1289), .B(n_1207), .C(n_1208), .Y(n_1343) );
OAI31xp33_ASAP7_75t_L g1344 ( .A1(n_1315), .A2(n_1215), .A3(n_1227), .B(n_1220), .Y(n_1344) );
NAND3xp33_ASAP7_75t_SL g1345 ( .A(n_1328), .B(n_1341), .C(n_1331), .Y(n_1345) );
NAND2xp5_ASAP7_75t_L g1346 ( .A(n_1335), .B(n_1330), .Y(n_1346) );
INVx2_ASAP7_75t_L g1347 ( .A(n_1333), .Y(n_1347) );
BUFx3_ASAP7_75t_L g1348 ( .A(n_1337), .Y(n_1348) );
AND2x4_ASAP7_75t_L g1349 ( .A(n_1327), .B(n_1339), .Y(n_1349) );
NOR3x2_ASAP7_75t_L g1350 ( .A(n_1348), .B(n_1342), .C(n_1336), .Y(n_1350) );
AOI22xp33_ASAP7_75t_L g1351 ( .A1(n_1345), .A2(n_1334), .B1(n_1338), .B2(n_1332), .Y(n_1351) );
NAND2xp5_ASAP7_75t_L g1352 ( .A(n_1346), .B(n_1343), .Y(n_1352) );
OAI322xp33_ASAP7_75t_L g1353 ( .A1(n_1347), .A2(n_1340), .A3(n_1323), .B1(n_1329), .B2(n_1215), .C1(n_1343), .C2(n_1344), .Y(n_1353) );
INVx1_ASAP7_75t_SL g1354 ( .A(n_1350), .Y(n_1354) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1352), .Y(n_1355) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1353), .Y(n_1356) );
OAI22xp33_ASAP7_75t_L g1357 ( .A1(n_1356), .A2(n_1349), .B1(n_1347), .B2(n_1351), .Y(n_1357) );
AOI22xp33_ASAP7_75t_L g1358 ( .A1(n_1357), .A2(n_1354), .B1(n_1355), .B2(n_1349), .Y(n_1358) );
AOI21xp5_ASAP7_75t_L g1359 ( .A1(n_1358), .A2(n_1189), .B(n_1195), .Y(n_1359) );
endmodule