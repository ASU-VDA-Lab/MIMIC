module fake_jpeg_24162_n_338 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx2_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx4f_ASAP7_75t_SL g65 ( 
.A(n_35),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_19),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_42),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_16),
.B(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_17),
.B1(n_29),
.B2(n_22),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_45),
.A2(n_36),
.B1(n_22),
.B2(n_29),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_36),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_29),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_42),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_57),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_33),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_61),
.Y(n_71)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_75),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_48),
.A2(n_38),
.B1(n_40),
.B2(n_56),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_70),
.A2(n_72),
.B1(n_34),
.B2(n_67),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_40),
.B1(n_38),
.B2(n_22),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_73),
.A2(n_17),
.B1(n_30),
.B2(n_32),
.Y(n_101)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

CKINVDCx6p67_ASAP7_75t_R g112 ( 
.A(n_82),
.Y(n_112)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_83),
.B(n_88),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_33),
.B1(n_29),
.B2(n_40),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_84),
.A2(n_33),
.B1(n_32),
.B2(n_30),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_20),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_87),
.Y(n_103)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_62),
.B(n_24),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_20),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_89),
.B(n_90),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_60),
.B(n_24),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_21),
.Y(n_107)
);

BUFx16f_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_94),
.B(n_106),
.Y(n_146)
);

OA21x2_ASAP7_75t_L g139 ( 
.A1(n_95),
.A2(n_104),
.B(n_112),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_27),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_97),
.B(n_103),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_101),
.B1(n_105),
.B2(n_116),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx3_ASAP7_75t_SL g130 ( 
.A(n_99),
.Y(n_130)
);

AND2x4_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_84),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_104),
.A2(n_39),
.B(n_16),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_70),
.A2(n_34),
.B1(n_50),
.B2(n_67),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_84),
.Y(n_124)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

NOR3xp33_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_30),
.C(n_32),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_113),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_68),
.A2(n_53),
.B1(n_17),
.B2(n_58),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_117),
.B(n_16),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_75),
.A2(n_58),
.B1(n_44),
.B2(n_31),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_69),
.A2(n_17),
.B1(n_28),
.B2(n_25),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

INVxp33_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

BUFx10_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_112),
.Y(n_121)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_123),
.A2(n_132),
.B(n_141),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_124),
.B(n_126),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_76),
.C(n_74),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_96),
.C(n_114),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_102),
.B(n_27),
.Y(n_126)
);

FAx1_ASAP7_75t_SL g127 ( 
.A(n_104),
.B(n_84),
.CI(n_39),
.CON(n_127),
.SN(n_127)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_137),
.C(n_139),
.Y(n_164)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_95),
.B(n_105),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_109),
.B(n_27),
.Y(n_136)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_137),
.A2(n_28),
.B(n_26),
.Y(n_172)
);

OA21x2_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_112),
.B(n_54),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_98),
.B(n_54),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_95),
.A2(n_34),
.B1(n_77),
.B2(n_93),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_142),
.A2(n_118),
.B1(n_69),
.B2(n_93),
.Y(n_156)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_143),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_119),
.B(n_24),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_141),
.A2(n_95),
.B1(n_101),
.B2(n_120),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_142),
.B1(n_127),
.B2(n_140),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_151),
.A2(n_164),
.B(n_167),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_165),
.C(n_170),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_97),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_154),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_86),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_134),
.A2(n_111),
.B1(n_106),
.B2(n_77),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_155),
.A2(n_156),
.B1(n_159),
.B2(n_163),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_134),
.A2(n_54),
.B1(n_63),
.B2(n_46),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_131),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_124),
.B(n_119),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_L g167 ( 
.A1(n_123),
.A2(n_0),
.B(n_110),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_146),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_169),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_124),
.B(n_64),
.C(n_66),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_172),
.A2(n_122),
.B(n_147),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_131),
.A2(n_20),
.B1(n_25),
.B2(n_26),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_138),
.Y(n_187)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

INVx11_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_139),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_189),
.C(n_121),
.Y(n_213)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_182),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_179),
.A2(n_184),
.B1(n_130),
.B2(n_110),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_135),
.Y(n_180)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_150),
.A2(n_127),
.B1(n_129),
.B2(n_128),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_186),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_155),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_187),
.Y(n_202)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_133),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_149),
.B(n_153),
.Y(n_190)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_122),
.Y(n_192)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_193),
.A2(n_196),
.B1(n_158),
.B2(n_152),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_145),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_194),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_195),
.A2(n_197),
.B(n_200),
.Y(n_209)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_164),
.A2(n_147),
.B(n_143),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_145),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_198),
.Y(n_201)
);

AO22x2_ASAP7_75t_L g199 ( 
.A1(n_151),
.A2(n_63),
.B1(n_46),
.B2(n_140),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_SL g205 ( 
.A1(n_199),
.A2(n_151),
.B(n_167),
.C(n_63),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_170),
.A2(n_121),
.B(n_130),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_205),
.A2(n_178),
.B1(n_191),
.B2(n_174),
.Y(n_236)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_206),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_183),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_210),
.B(n_216),
.Y(n_228)
);

AO21x1_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_166),
.B(n_171),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_212),
.A2(n_222),
.B(n_217),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_214),
.C(n_224),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_119),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_180),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_199),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_219),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

INVxp33_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_197),
.A2(n_130),
.B(n_94),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_174),
.A2(n_94),
.B(n_51),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_223),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_177),
.B(n_52),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_176),
.B(n_49),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_181),
.C(n_189),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_195),
.Y(n_227)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_204),
.B(n_175),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_235),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_208),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_230),
.A2(n_1),
.B(n_2),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_200),
.Y(n_232)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_232),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_234),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_225),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_236),
.A2(n_243),
.B1(n_246),
.B2(n_247),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_224),
.C(n_223),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_239),
.A2(n_21),
.B(n_2),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_201),
.B(n_212),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_240),
.Y(n_257)
);

NOR4xp25_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_190),
.C(n_181),
.D(n_191),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_1),
.Y(n_259)
);

NAND5xp2_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_21),
.C(n_18),
.D(n_37),
.E(n_43),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_220),
.A2(n_213),
.B1(n_209),
.B2(n_205),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_205),
.A2(n_17),
.B1(n_55),
.B2(n_64),
.Y(n_247)
);

INVx13_ASAP7_75t_L g248 ( 
.A(n_211),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_1),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_242),
.A2(n_202),
.B1(n_207),
.B2(n_205),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_250),
.A2(n_251),
.B1(n_265),
.B2(n_266),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_219),
.B1(n_222),
.B2(n_215),
.Y(n_251)
);

XOR2x2_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_232),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_252),
.B(n_259),
.Y(n_272)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_254),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_256),
.C(n_264),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_214),
.C(n_37),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_245),
.Y(n_261)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_261),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_18),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_242),
.A2(n_43),
.B1(n_41),
.B2(n_37),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_SL g267 ( 
.A1(n_239),
.A2(n_43),
.B(n_41),
.C(n_21),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_267),
.A2(n_21),
.B1(n_41),
.B2(n_18),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_268),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_231),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_282),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_230),
.Y(n_274)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_274),
.Y(n_300)
);

XOR2x2_ASAP7_75t_SL g275 ( 
.A(n_252),
.B(n_237),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_275),
.B(n_21),
.Y(n_299)
);

INVx4_ASAP7_75t_SL g276 ( 
.A(n_261),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_265),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_260),
.A2(n_233),
.B1(n_244),
.B2(n_227),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_277),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_240),
.C(n_228),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_283),
.C(n_257),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_248),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_279),
.B(n_267),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_236),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_249),
.B(n_243),
.C(n_247),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_284),
.Y(n_292)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_258),
.C(n_251),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_290),
.Y(n_301)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_288),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_259),
.C(n_267),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_270),
.B(n_267),
.C(n_3),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_293),
.B(n_295),
.Y(n_312)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_294),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_2),
.C(n_4),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_18),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_5),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_283),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_297),
.A2(n_4),
.B(n_5),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_4),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_298),
.A2(n_292),
.B1(n_7),
.B2(n_8),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_5),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_297),
.A2(n_281),
.B1(n_276),
.B2(n_275),
.Y(n_303)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_303),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_292),
.A2(n_280),
.B1(n_269),
.B2(n_273),
.Y(n_304)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_304),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_15),
.C(n_8),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_310),
.Y(n_314)
);

FAx1_ASAP7_75t_SL g309 ( 
.A(n_299),
.B(n_291),
.CI(n_300),
.CON(n_309),
.SN(n_309)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_311),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_301),
.A2(n_289),
.B1(n_8),
.B2(n_9),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_317),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_306),
.A2(n_307),
.B1(n_302),
.B2(n_305),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_6),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_319),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_6),
.Y(n_321)
);

AND2x2_ASAP7_75t_SL g327 ( 
.A(n_321),
.B(n_6),
.Y(n_327)
);

INVx11_ASAP7_75t_L g323 ( 
.A(n_321),
.Y(n_323)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_323),
.Y(n_331)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_312),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_324),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_310),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_326),
.C(n_327),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_320),
.C(n_316),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_330),
.B(n_328),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_331),
.B(n_329),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_333),
.A2(n_322),
.B(n_328),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_334),
.A2(n_11),
.B(n_12),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_335),
.A2(n_11),
.B(n_13),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_336),
.B(n_14),
.Y(n_337)
);

OA21x2_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_14),
.B(n_210),
.Y(n_338)
);


endmodule