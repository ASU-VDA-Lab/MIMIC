module fake_jpeg_21166_n_214 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_214);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_214;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_20),
.B(n_2),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_37),
.Y(n_59)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_11),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_2),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_40),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_9),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_17),
.B(n_28),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_60),
.B(n_40),
.Y(n_66)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_53),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_55),
.B(n_3),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_25),
.B1(n_28),
.B2(n_13),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_61),
.B1(n_15),
.B2(n_42),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_25),
.B1(n_21),
.B2(n_24),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_35),
.B1(n_36),
.B2(n_5),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_32),
.A2(n_33),
.B(n_37),
.C(n_43),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_21),
.B1(n_18),
.B2(n_24),
.Y(n_61)
);

NOR2x1_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_18),
.Y(n_63)
);

OR2x2_ASAP7_75t_SL g93 ( 
.A(n_63),
.B(n_26),
.Y(n_93)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_66),
.A2(n_82),
.B1(n_85),
.B2(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_44),
.B(n_15),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_67),
.B(n_73),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_69),
.A2(n_47),
.B1(n_56),
.B2(n_6),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_36),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_70),
.B(n_97),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_45),
.A2(n_35),
.B1(n_31),
.B2(n_19),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_36),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_98),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_27),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_27),
.Y(n_74)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_77),
.Y(n_106)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_14),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_80),
.Y(n_120)
);

BUFx8_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_41),
.B1(n_29),
.B2(n_23),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

HB1xp67_ASAP7_75t_SL g107 ( 
.A(n_87),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_14),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_89),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_57),
.B(n_63),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_53),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_93),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_64),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_95),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_65),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_29),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_78),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_97),
.A2(n_52),
.B(n_26),
.C(n_19),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_113),
.B(n_99),
.C(n_84),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_110),
.A2(n_114),
.B1(n_119),
.B2(n_82),
.Y(n_141)
);

OR2x6_ASAP7_75t_SL g113 ( 
.A(n_93),
.B(n_39),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_66),
.A2(n_29),
.B1(n_23),
.B2(n_6),
.Y(n_114)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_70),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_4),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_92),
.Y(n_132)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_140),
.Y(n_156)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_107),
.A2(n_90),
.B(n_92),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_134),
.A2(n_124),
.B(n_119),
.Y(n_162)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_135),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_125),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_136),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_118),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_137),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_90),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_139),
.C(n_144),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_86),
.C(n_68),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_141),
.A2(n_123),
.B1(n_101),
.B2(n_112),
.Y(n_149)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_143),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_94),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_94),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_146),
.A2(n_147),
.B(n_113),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_113),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_141),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_149),
.A2(n_131),
.B1(n_134),
.B2(n_143),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_153),
.A2(n_157),
.B(n_145),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_147),
.A2(n_101),
.B(n_115),
.Y(n_157)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_117),
.A3(n_106),
.B1(n_120),
.B2(n_108),
.C1(n_110),
.C2(n_122),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_L g176 ( 
.A1(n_160),
.A2(n_133),
.B(n_124),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_145),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_150),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_164),
.B(n_167),
.Y(n_183)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_163),
.Y(n_165)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_144),
.C(n_139),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_154),
.C(n_148),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_128),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_132),
.Y(n_168)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_152),
.B(n_156),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_169),
.A2(n_171),
.B1(n_174),
.B2(n_176),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_150),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_170),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_L g179 ( 
.A1(n_172),
.A2(n_163),
.B(n_153),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_175),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_127),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_177),
.A2(n_172),
.B1(n_151),
.B2(n_164),
.Y(n_182)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_186),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_182),
.A2(n_161),
.B1(n_158),
.B2(n_155),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_148),
.C(n_149),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_102),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_165),
.A2(n_162),
.B1(n_151),
.B2(n_157),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_187),
.A2(n_155),
.B1(n_105),
.B2(n_79),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_179),
.A2(n_175),
.B(n_173),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_192),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_190),
.A2(n_194),
.B1(n_195),
.B2(n_142),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_183),
.A2(n_161),
.B(n_158),
.Y(n_191)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_191),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_185),
.A2(n_105),
.B1(n_103),
.B2(n_75),
.Y(n_194)
);

MAJx2_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_189),
.C(n_192),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_193),
.A2(n_188),
.B1(n_178),
.B2(n_184),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_199),
.Y(n_203)
);

NAND4xp25_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_188),
.C(n_181),
.D(n_180),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_202),
.Y(n_206)
);

OAI321xp33_ASAP7_75t_L g204 ( 
.A1(n_198),
.A2(n_184),
.A3(n_180),
.B1(n_196),
.B2(n_8),
.C(n_9),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_204),
.B(n_205),
.Y(n_207)
);

FAx1_ASAP7_75t_SL g205 ( 
.A(n_197),
.B(n_9),
.CI(n_83),
.CON(n_205),
.SN(n_205)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_201),
.C(n_200),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_208),
.B(n_81),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_206),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_209),
.A2(n_205),
.B1(n_201),
.B2(n_96),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_210),
.B(n_211),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_211),
.C(n_207),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_96),
.Y(n_214)
);


endmodule