module fake_jpeg_14872_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_12),
.B(n_6),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

CKINVDCx6p67_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_12),
.Y(n_48)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_31),
.A2(n_25),
.B(n_22),
.Y(n_44)
);

NAND2xp33_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_18),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_32),
.B1(n_28),
.B2(n_26),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_45),
.A2(n_54),
.B1(n_63),
.B2(n_15),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_43),
.A2(n_23),
.B1(n_13),
.B2(n_18),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_47),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_48),
.B(n_49),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_30),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_52),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_21),
.Y(n_52)
);

AND2x6_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_7),
.Y(n_53)
);

AND2x6_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_7),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_13),
.B1(n_14),
.B2(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_57),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_62),
.A2(n_47),
.B1(n_59),
.B2(n_61),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_13),
.B1(n_18),
.B2(n_12),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_21),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_14),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_61),
.B(n_47),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_49),
.A2(n_13),
.B1(n_21),
.B2(n_14),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_68),
.A2(n_70),
.B1(n_74),
.B2(n_77),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_14),
.B1(n_36),
.B2(n_24),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_50),
.B(n_22),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_76),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_48),
.B(n_22),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_52),
.B(n_17),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_79),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_29),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_54),
.C(n_51),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_51),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_83),
.B(n_84),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_75),
.B(n_64),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_69),
.A2(n_77),
.B1(n_79),
.B2(n_75),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_88),
.B1(n_19),
.B2(n_20),
.Y(n_109)
);

AOI22x1_ASAP7_75t_L g88 ( 
.A1(n_69),
.A2(n_46),
.B1(n_53),
.B2(n_63),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_90),
.C(n_92),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_82),
.B(n_19),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_91),
.A2(n_72),
.B1(n_62),
.B2(n_56),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_29),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_55),
.C(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_65),
.Y(n_100)
);

INVxp67_ASAP7_75t_SL g94 ( 
.A(n_66),
.Y(n_94)
);

INVxp33_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_62),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_96),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_97),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_87),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_102),
.A2(n_108),
.B1(n_89),
.B2(n_41),
.Y(n_110)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_19),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_74),
.B(n_16),
.C(n_17),
.Y(n_105)
);

A2O1A1O1Ixp25_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_19),
.B(n_20),
.C(n_16),
.D(n_3),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_71),
.B(n_66),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_106),
.A2(n_109),
.B(n_41),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_71),
.B1(n_60),
.B2(n_56),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_110),
.A2(n_111),
.B1(n_114),
.B2(n_115),
.Y(n_123)
);

AO22x1_ASAP7_75t_L g111 ( 
.A1(n_109),
.A2(n_85),
.B1(n_90),
.B2(n_92),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_116),
.C(n_107),
.Y(n_119)
);

NAND3xp33_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_86),
.C(n_105),
.Y(n_113)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_117),
.B(n_6),
.C(n_1),
.D(n_2),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_104),
.A2(n_15),
.B1(n_25),
.B2(n_24),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_24),
.B1(n_17),
.B2(n_16),
.Y(n_115)
);

OAI321xp33_ASAP7_75t_L g122 ( 
.A1(n_118),
.A2(n_106),
.A3(n_98),
.B1(n_99),
.B2(n_19),
.C(n_20),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_120),
.C(n_121),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_107),
.C(n_101),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_103),
.C(n_102),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_124),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_115),
.Y(n_125)
);

AOI321xp33_ASAP7_75t_L g128 ( 
.A1(n_120),
.A2(n_111),
.A3(n_117),
.B1(n_2),
.B2(n_5),
.C(n_8),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_128),
.A2(n_127),
.B(n_125),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_8),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_129),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_126),
.A2(n_2),
.B(n_5),
.C(n_9),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_132),
.A2(n_10),
.B(n_11),
.Y(n_134)
);

OAI21x1_ASAP7_75t_SL g135 ( 
.A1(n_134),
.A2(n_132),
.B(n_131),
.Y(n_135)
);

BUFx24_ASAP7_75t_SL g136 ( 
.A(n_135),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_133),
.Y(n_137)
);


endmodule