module real_jpeg_24093_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_206;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_1),
.A2(n_37),
.B1(n_39),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_1),
.A2(n_43),
.B1(n_55),
.B2(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_1),
.A2(n_49),
.B1(n_50),
.B2(n_55),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_1),
.A2(n_55),
.B1(n_63),
.B2(n_64),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_2),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_4),
.A2(n_63),
.B1(n_64),
.B2(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_4),
.Y(n_90)
);

INVx8_ASAP7_75t_SL g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_6),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_6),
.B(n_36),
.Y(n_168)
);

O2A1O1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_6),
.A2(n_39),
.B(n_51),
.C(n_198),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_6),
.A2(n_37),
.B1(n_39),
.B2(n_114),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_6),
.B(n_64),
.C(n_81),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_6),
.A2(n_49),
.B1(n_50),
.B2(n_114),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_6),
.A2(n_61),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_6),
.B(n_109),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_7),
.A2(n_37),
.B1(n_39),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_7),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_7),
.A2(n_47),
.B1(n_63),
.B2(n_64),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_8),
.A2(n_27),
.B1(n_37),
.B2(n_39),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_8),
.A2(n_27),
.B1(n_49),
.B2(n_50),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_8),
.A2(n_27),
.B1(n_63),
.B2(n_64),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_10),
.A2(n_28),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_10),
.A2(n_37),
.B1(n_39),
.B2(n_41),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_10),
.A2(n_41),
.B1(n_49),
.B2(n_50),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_10),
.A2(n_41),
.B1(n_63),
.B2(n_64),
.Y(n_226)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_12),
.A2(n_63),
.B1(n_64),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_12),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_12),
.A2(n_49),
.B1(n_50),
.B2(n_75),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_13),
.A2(n_49),
.B1(n_50),
.B2(n_86),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_13),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_13),
.A2(n_63),
.B1(n_64),
.B2(n_86),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_13),
.A2(n_37),
.B1(n_39),
.B2(n_86),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_14),
.A2(n_63),
.B1(n_64),
.B2(n_70),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_14),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_14),
.A2(n_49),
.B1(n_50),
.B2(n_70),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_16),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_16),
.A2(n_62),
.B1(n_69),
.B2(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_16),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_16),
.A2(n_62),
.B1(n_223),
.B2(n_225),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_145),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_143),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_120),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_20),
.B(n_120),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_87),
.C(n_98),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_21),
.A2(n_22),
.B1(n_87),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_59),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_44),
.B2(n_45),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_25),
.B(n_44),
.C(n_59),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_36),
.B2(n_40),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_26),
.Y(n_100)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_29),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_30),
.B(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_30),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_30),
.A2(n_140),
.B(n_159),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_35),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_32),
.A2(n_33),
.B1(n_37),
.B2(n_39),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_32),
.A2(n_37),
.B(n_113),
.C(n_115),
.Y(n_112)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND3xp33_ASAP7_75t_SL g115 ( 
.A(n_33),
.B(n_39),
.C(n_116),
.Y(n_115)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_34),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_35),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_35),
.B(n_103),
.Y(n_140)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_SL g39 ( 
.A(n_37),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_39),
.B1(n_51),
.B2(n_52),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_40),
.Y(n_137)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_43),
.B(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_48),
.B(n_53),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_46),
.A2(n_48),
.B1(n_57),
.B2(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_48),
.A2(n_53),
.B(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_49),
.A2(n_50),
.B1(n_81),
.B2(n_83),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_49),
.A2(n_52),
.B(n_114),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_50),
.B(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_56),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_54),
.B(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_56),
.A2(n_107),
.B1(n_109),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_57),
.A2(n_106),
.B(n_108),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g209 ( 
.A1(n_57),
.A2(n_108),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_76),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_60),
.B(n_76),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_68),
.B1(n_71),
.B2(n_74),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_61),
.A2(n_74),
.B1(n_89),
.B2(n_91),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_61),
.A2(n_89),
.B(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_61),
.A2(n_119),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_61),
.A2(n_226),
.B(n_232),
.Y(n_246)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_62),
.B(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_64),
.B1(n_81),
.B2(n_83),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_63),
.B(n_230),
.Y(n_229)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_84),
.B2(n_85),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_77),
.A2(n_84),
.B(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_78),
.A2(n_192),
.B(n_194),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_78),
.A2(n_194),
.B(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_79),
.A2(n_94),
.B1(n_95),
.B2(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_79),
.B(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_79),
.A2(n_95),
.B1(n_193),
.B2(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_84),
.Y(n_79)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_81),
.Y(n_83)
);

BUFx24_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_84),
.B(n_114),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_84),
.A2(n_156),
.B(n_207),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_87),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_92),
.B1(n_96),
.B2(n_97),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_88),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_97),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_91),
.B(n_114),
.Y(n_230)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_91),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_91),
.A2(n_200),
.B(n_224),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_92),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_95),
.B(n_157),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_98),
.B(n_265),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_105),
.C(n_110),
.Y(n_98)
);

FAx1_ASAP7_75t_SL g173 ( 
.A(n_99),
.B(n_105),
.CI(n_110),
.CON(n_173),
.SN(n_173)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_117),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_111),
.A2(n_112),
.B1(n_117),
.B2(n_163),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_113),
.A2(n_114),
.B(n_160),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_117),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_142),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_130),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_126),
.B2(n_127),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_141),
.Y(n_130)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B(n_139),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_179),
.B(n_263),
.C(n_268),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_172),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_147),
.B(n_172),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_161),
.C(n_164),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_148),
.A2(n_149),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_158),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_154),
.B2(n_155),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_154),
.C(n_158),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_153),
.Y(n_166)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_161),
.A2(n_162),
.B1(n_164),
.B2(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_164),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.C(n_169),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_170),
.A2(n_171),
.B(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_178),
.Y(n_172)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_173),
.Y(n_178)
);

BUFx24_ASAP7_75t_SL g270 ( 
.A(n_173),
.Y(n_270)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_176),
.B(n_177),
.C(n_178),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_256),
.B(n_262),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_211),
.B(n_255),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_203),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_184),
.B(n_203),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_189),
.B2(n_202),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_185),
.B(n_191),
.C(n_195),
.Y(n_261)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_195),
.B2(n_196),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_197),
.B(n_199),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.C(n_208),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_204),
.B(n_251),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_205),
.A2(n_208),
.B1(n_209),
.B2(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_205),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_249),
.B(n_254),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_239),
.B(n_248),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_227),
.B(n_238),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_222),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_222),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_219),
.Y(n_247)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_234),
.B(n_237),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_236),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_247),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_247),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_246),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_245),
.C(n_246),
.Y(n_253)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_253),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_253),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_261),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_261),
.Y(n_262)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_267),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_267),
.Y(n_268)
);


endmodule