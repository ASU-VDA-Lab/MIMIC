module fake_jpeg_21094_n_292 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_292);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_292;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_266;
wire n_218;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_44),
.Y(n_55)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_20),
.B(n_7),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_47),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_20),
.B(n_7),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_49),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_28),
.B(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_30),
.Y(n_88)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_16),
.B1(n_33),
.B2(n_37),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_53),
.A2(n_76),
.B1(n_91),
.B2(n_99),
.Y(n_107)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_57),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_28),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_22),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_58),
.B(n_60),
.Y(n_104)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

CKINVDCx12_ASAP7_75t_R g63 ( 
.A(n_41),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_64),
.B(n_67),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_49),
.B(n_21),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_66),
.B(n_68),
.Y(n_125)
);

CKINVDCx12_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_43),
.Y(n_68)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_72),
.B(n_74),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_73),
.Y(n_115)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_29),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_75),
.B(n_80),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_40),
.A2(n_16),
.B1(n_33),
.B2(n_22),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_77),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_38),
.A2(n_16),
.B1(n_33),
.B2(n_30),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_78),
.A2(n_94),
.B1(n_97),
.B2(n_34),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_17),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_18),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_83),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_82),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_48),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_84),
.B(n_86),
.Y(n_127)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_88),
.Y(n_124)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_50),
.A2(n_18),
.B1(n_21),
.B2(n_17),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

CKINVDCx12_ASAP7_75t_R g94 ( 
.A(n_51),
.Y(n_94)
);

BUFx10_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_25),
.Y(n_130)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_45),
.B(n_29),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_27),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_38),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_69),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_24),
.C(n_25),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_79),
.C(n_71),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_78),
.A2(n_19),
.B1(n_35),
.B2(n_27),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_118),
.B1(n_131),
.B2(n_90),
.Y(n_138)
);

AO22x1_ASAP7_75t_SL g116 ( 
.A1(n_99),
.A2(n_34),
.B1(n_25),
.B2(n_24),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_116),
.A2(n_89),
.B1(n_52),
.B2(n_100),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_83),
.A2(n_19),
.B1(n_31),
.B2(n_26),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_34),
.B1(n_19),
.B2(n_31),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_119),
.A2(n_117),
.B(n_115),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_122),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_130),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_55),
.A2(n_26),
.B1(n_24),
.B2(n_34),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_132),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_127),
.B(n_75),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_144),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_134),
.A2(n_164),
.B(n_109),
.Y(n_172)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_136),
.A2(n_103),
.B1(n_117),
.B2(n_115),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_138),
.A2(n_140),
.B1(n_151),
.B2(n_153),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_139),
.A2(n_142),
.B1(n_148),
.B2(n_150),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_53),
.B1(n_89),
.B2(n_100),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_141),
.B(n_146),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_107),
.A2(n_52),
.B1(n_70),
.B2(n_96),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_143),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_124),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_105),
.A2(n_112),
.B1(n_114),
.B2(n_124),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_145),
.A2(n_1),
.B(n_2),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_62),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_73),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_149),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_70),
.B1(n_65),
.B2(n_82),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_116),
.A2(n_71),
.B1(n_65),
.B2(n_92),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_116),
.A2(n_114),
.B1(n_113),
.B2(n_102),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_102),
.B(n_36),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_158),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_116),
.A2(n_93),
.B1(n_79),
.B2(n_61),
.Y(n_153)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_154),
.Y(n_183)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_114),
.A2(n_104),
.B1(n_125),
.B2(n_131),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_156),
.A2(n_159),
.B1(n_111),
.B2(n_110),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_95),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_157),
.B(n_161),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_104),
.B(n_95),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_105),
.A2(n_7),
.B1(n_15),
.B2(n_14),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_119),
.B(n_129),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_162),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_6),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_119),
.A2(n_36),
.B(n_6),
.C(n_9),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_163),
.B(n_121),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_119),
.A2(n_106),
.B(n_109),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_120),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_165),
.B(n_168),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_106),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_SL g197 ( 
.A(n_169),
.B(n_173),
.C(n_186),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_163),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_177),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_101),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_174),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_172),
.A2(n_182),
.B(n_161),
.Y(n_206)
);

NOR2x1_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_121),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_101),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_158),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_178),
.B(n_193),
.Y(n_201)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_135),
.A2(n_103),
.B(n_111),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_110),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_191),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_L g186 ( 
.A1(n_160),
.A2(n_0),
.B(n_1),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_133),
.B(n_5),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_188),
.B(n_189),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_141),
.B(n_5),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_137),
.B(n_0),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_137),
.B(n_1),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_195),
.A2(n_186),
.B1(n_173),
.B2(n_177),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_151),
.B(n_2),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_138),
.Y(n_210)
);

OAI32xp33_ASAP7_75t_L g199 ( 
.A1(n_196),
.A2(n_145),
.A3(n_164),
.B1(n_152),
.B2(n_134),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_212),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_149),
.C(n_135),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_176),
.C(n_179),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_202),
.A2(n_206),
.B(n_215),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_188),
.B(n_146),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_204),
.B(n_207),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_187),
.B(n_159),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_167),
.A2(n_150),
.B1(n_139),
.B2(n_153),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_209),
.A2(n_217),
.B1(n_178),
.B2(n_184),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_210),
.B(n_214),
.Y(n_237)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_181),
.Y(n_211)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_136),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_140),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_195),
.A2(n_155),
.B1(n_154),
.B2(n_148),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_185),
.A2(n_2),
.B(n_3),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_195),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_167),
.A2(n_5),
.B1(n_9),
.B2(n_10),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_171),
.Y(n_219)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_219),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_228),
.C(n_234),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_200),
.B(n_179),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_227),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_205),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_224),
.B(n_225),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_198),
.B(n_189),
.Y(n_225)
);

OR2x2_ASAP7_75t_SL g226 ( 
.A(n_197),
.B(n_173),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_226),
.A2(n_216),
.B1(n_197),
.B2(n_199),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_213),
.C(n_206),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_205),
.Y(n_230)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_230),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_233),
.A2(n_238),
.B1(n_209),
.B2(n_214),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_174),
.C(n_172),
.Y(n_234)
);

AOI221xp5_ASAP7_75t_L g235 ( 
.A1(n_207),
.A2(n_185),
.B1(n_180),
.B2(n_175),
.C(n_187),
.Y(n_235)
);

BUFx24_ASAP7_75t_SL g244 ( 
.A(n_235),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_175),
.C(n_180),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_203),
.C(n_202),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_210),
.A2(n_190),
.B1(n_168),
.B2(n_191),
.Y(n_238)
);

BUFx12_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_245),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_203),
.Y(n_241)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_241),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_246),
.Y(n_264)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_249),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_208),
.C(n_211),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_250),
.Y(n_261)
);

AO221x1_ASAP7_75t_L g251 ( 
.A1(n_222),
.A2(n_166),
.B1(n_212),
.B2(n_183),
.C(n_192),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_251),
.A2(n_252),
.B1(n_198),
.B2(n_234),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_204),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_223),
.Y(n_253)
);

NOR3xp33_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_170),
.C(n_229),
.Y(n_260)
);

OA21x2_ASAP7_75t_SL g254 ( 
.A1(n_240),
.A2(n_231),
.B(n_227),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_242),
.C(n_250),
.Y(n_269)
);

OAI21xp33_ASAP7_75t_L g255 ( 
.A1(n_240),
.A2(n_232),
.B(n_247),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_242),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_241),
.A2(n_233),
.B1(n_232),
.B2(n_238),
.Y(n_257)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_257),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_248),
.A2(n_231),
.B(n_249),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_258),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_260),
.A2(n_208),
.B1(n_165),
.B2(n_183),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_246),
.A2(n_237),
.B(n_182),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_266),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_263),
.B(n_239),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_243),
.A2(n_201),
.B(n_215),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_SL g267 ( 
.A1(n_257),
.A2(n_217),
.B(n_190),
.C(n_228),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_267),
.A2(n_271),
.B(n_218),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_270),
.C(n_274),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_269),
.A2(n_275),
.B(n_273),
.Y(n_281)
);

A2O1A1Ixp33_ASAP7_75t_SL g271 ( 
.A1(n_258),
.A2(n_220),
.B(n_201),
.C(n_169),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_239),
.Y(n_274)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_267),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_280),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_261),
.C(n_264),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_271),
.C(n_218),
.Y(n_285)
);

AOI322xp5_ASAP7_75t_L g280 ( 
.A1(n_276),
.A2(n_265),
.A3(n_266),
.B1(n_244),
.B2(n_262),
.C1(n_259),
.C2(n_254),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_281),
.A2(n_282),
.B(n_271),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_283),
.B(n_285),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_277),
.A2(n_259),
.B1(n_267),
.B2(n_256),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_279),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_286),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_288),
.B(n_289),
.Y(n_290)
);

BUFx24_ASAP7_75t_SL g291 ( 
.A(n_290),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_287),
.Y(n_292)
);


endmodule