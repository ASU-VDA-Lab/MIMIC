module fake_jpeg_13481_n_177 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_177);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_10),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_5),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_2),
.B(n_43),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx4f_ASAP7_75t_SL g71 ( 
.A(n_49),
.Y(n_71)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_1),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_51),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_55),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_84),
.Y(n_99)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_61),
.B(n_0),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_0),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_3),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_67),
.B1(n_53),
.B2(n_65),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_90),
.A2(n_100),
.B1(n_82),
.B2(n_72),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_81),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_93),
.B(n_95),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_53),
.B1(n_58),
.B2(n_59),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_52),
.B1(n_6),
.B2(n_7),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_57),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_1),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_75),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_66),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_65),
.B1(n_54),
.B2(n_72),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_113),
.B1(n_115),
.B2(n_116),
.Y(n_121)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_100),
.A2(n_54),
.B1(n_69),
.B2(n_64),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_103),
.A2(n_118),
.B1(n_8),
.B2(n_9),
.Y(n_128)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_99),
.A2(n_74),
.B1(n_68),
.B2(n_63),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_105),
.A2(n_11),
.B(n_12),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_106),
.B(n_112),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_119),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_66),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_111),
.Y(n_137)
);

AND2x6_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_25),
.Y(n_110)
);

FAx1_ASAP7_75t_SL g131 ( 
.A(n_110),
.B(n_115),
.CI(n_101),
.CON(n_131),
.SN(n_131)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_88),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_60),
.B1(n_70),
.B2(n_62),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_73),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_120),
.Y(n_126)
);

AO21x2_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_52),
.B(n_20),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_116)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_117),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_88),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_50),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_128),
.Y(n_147)
);

NAND2x1p5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_7),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_16),
.B(n_18),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_8),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_138),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_136),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_115),
.B(n_26),
.Y(n_132)
);

A2O1A1O1Ixp25_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_24),
.B(n_27),
.C(n_29),
.D(n_30),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_9),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_133),
.B(n_134),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_11),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_12),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

OAI22x1_ASAP7_75t_L g142 ( 
.A1(n_131),
.A2(n_121),
.B1(n_128),
.B2(n_132),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_124),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_143),
.A2(n_123),
.B1(n_136),
.B2(n_127),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_13),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_144),
.B(n_153),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_155),
.Y(n_164)
);

AOI21xp33_ASAP7_75t_L g146 ( 
.A1(n_137),
.A2(n_19),
.B(n_22),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_146),
.A2(n_150),
.B(n_31),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_122),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_130),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_142),
.B(n_137),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_159),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_148),
.A2(n_125),
.B(n_139),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_149),
.B(n_36),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_161),
.A2(n_165),
.B1(n_145),
.B2(n_144),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_147),
.A2(n_38),
.B1(n_45),
.B2(n_46),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_164),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_162),
.B1(n_157),
.B2(n_143),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_171),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_170),
.B1(n_162),
.B2(n_156),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_173),
.A2(n_167),
.B(n_163),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_168),
.B1(n_154),
.B2(n_151),
.Y(n_175)
);

NOR4xp25_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_146),
.C(n_168),
.D(n_150),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_152),
.Y(n_177)
);


endmodule