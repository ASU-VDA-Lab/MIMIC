module fake_aes_7440_n_24 (n_1, n_2, n_4, n_3, n_5, n_0, n_24);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_24;
wire n_20;
wire n_23;
wire n_8;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
wire n_6;
wire n_7;
CKINVDCx5p33_ASAP7_75t_R g6 ( .A(n_5), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_3), .Y(n_7) );
HB1xp67_ASAP7_75t_L g8 ( .A(n_0), .Y(n_8) );
CKINVDCx5p33_ASAP7_75t_R g9 ( .A(n_2), .Y(n_9) );
INVx1_ASAP7_75t_SL g10 ( .A(n_4), .Y(n_10) );
BUFx2_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
BUFx6f_ASAP7_75t_L g12 ( .A(n_7), .Y(n_12) );
INVx4_ASAP7_75t_L g13 ( .A(n_6), .Y(n_13) );
BUFx6f_ASAP7_75t_L g14 ( .A(n_9), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_13), .B(n_10), .Y(n_15) );
NAND2xp33_ASAP7_75t_R g16 ( .A(n_11), .B(n_0), .Y(n_16) );
OR2x2_ASAP7_75t_L g17 ( .A(n_15), .B(n_13), .Y(n_17) );
OR2x2_ASAP7_75t_L g18 ( .A(n_16), .B(n_14), .Y(n_18) );
NAND3xp33_ASAP7_75t_L g19 ( .A(n_17), .B(n_18), .C(n_14), .Y(n_19) );
NOR3xp33_ASAP7_75t_L g20 ( .A(n_19), .B(n_1), .C(n_12), .Y(n_20) );
INVx1_ASAP7_75t_SL g21 ( .A(n_20), .Y(n_21) );
BUFx6f_ASAP7_75t_L g22 ( .A(n_20), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
AOI22xp33_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_22), .B1(n_21), .B2(n_20), .Y(n_24) );
endmodule