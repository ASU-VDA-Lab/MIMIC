module fake_jpeg_9697_n_205 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_205);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_0),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_32),
.B1(n_18),
.B2(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_22),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_41),
.B(n_2),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_21),
.B(n_31),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_50),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_35),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_28),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_49),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_41),
.B(n_25),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_28),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_26),
.Y(n_82)
);

HB1xp67_ASAP7_75t_SL g69 ( 
.A(n_53),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_32),
.B1(n_18),
.B2(n_16),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_55),
.A2(n_24),
.B1(n_21),
.B2(n_25),
.Y(n_65)
);

OR2x4_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_23),
.Y(n_57)
);

NOR2x1_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_30),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_58),
.B(n_66),
.Y(n_94)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_59),
.B(n_60),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_61),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_35),
.C(n_37),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_62),
.A2(n_78),
.B(n_80),
.Y(n_99)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_63),
.B(n_67),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_73),
.B1(n_84),
.B2(n_29),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_31),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_70),
.B(n_75),
.Y(n_86)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_71),
.A2(n_27),
.B1(n_30),
.B2(n_8),
.Y(n_107)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

AO22x1_ASAP7_75t_SL g73 ( 
.A1(n_49),
.A2(n_51),
.B1(n_36),
.B2(n_39),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_2),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_76),
.B(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_3),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_40),
.C(n_37),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_15),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_79),
.B(n_81),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_4),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_4),
.Y(n_83)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

AO22x2_ASAP7_75t_L g84 ( 
.A1(n_54),
.A2(n_38),
.B1(n_23),
.B2(n_34),
.Y(n_84)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_104),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_73),
.B1(n_68),
.B2(n_82),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_92),
.B1(n_96),
.B2(n_97),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_27),
.B(n_64),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_73),
.A2(n_38),
.B1(n_40),
.B2(n_34),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_57),
.A2(n_26),
.B1(n_22),
.B2(n_19),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_6),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_61),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_105),
.B(n_6),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_107),
.Y(n_124)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_111),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_94),
.B(n_56),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_94),
.B(n_68),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_115),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_62),
.C(n_67),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_125),
.C(n_86),
.Y(n_138)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_95),
.B(n_67),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_116),
.A2(n_118),
.B(n_119),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_64),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_117),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_88),
.A2(n_65),
.B(n_80),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_93),
.B(n_90),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_7),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_74),
.Y(n_122)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_85),
.B(n_12),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_128),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_6),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_72),
.Y(n_126)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_92),
.B(n_7),
.Y(n_127)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_98),
.Y(n_129)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_129),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_130),
.B(n_149),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_128),
.A2(n_87),
.B1(n_103),
.B2(n_100),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_133),
.A2(n_136),
.B1(n_149),
.B2(n_137),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_100),
.B1(n_97),
.B2(n_89),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_140),
.C(n_143),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_89),
.C(n_91),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_141),
.B(n_147),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_91),
.C(n_93),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_90),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_146),
.A2(n_119),
.B(n_116),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_117),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_136),
.A2(n_124),
.B1(n_110),
.B2(n_120),
.Y(n_150)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_139),
.B1(n_142),
.B2(n_143),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_125),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_153),
.A2(n_155),
.B(n_160),
.Y(n_166)
);

OAI322xp33_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_118),
.A3(n_122),
.B1(n_113),
.B2(n_116),
.C1(n_115),
.C2(n_111),
.Y(n_154)
);

NOR3xp33_ASAP7_75t_SL g171 ( 
.A(n_154),
.B(n_123),
.C(n_109),
.Y(n_171)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_146),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_138),
.C(n_132),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_159),
.C(n_161),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_131),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_148),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_116),
.C(n_108),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_134),
.A2(n_127),
.B(n_124),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_141),
.B(n_133),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_9),
.C(n_10),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_163),
.Y(n_169)
);

OAI321xp33_ASAP7_75t_L g165 ( 
.A1(n_152),
.A2(n_135),
.A3(n_139),
.B1(n_145),
.B2(n_121),
.C(n_148),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_168),
.Y(n_179)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_162),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_71),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_173),
.C(n_175),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_11),
.C(n_12),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_170),
.A2(n_159),
.B(n_155),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_176),
.B(n_178),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_169),
.Y(n_177)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_170),
.A2(n_156),
.B(n_151),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_181),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_174),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_158),
.C(n_160),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_173),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_179),
.B(n_182),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_187),
.B(n_188),
.Y(n_194)
);

OAI211xp5_ASAP7_75t_L g189 ( 
.A1(n_181),
.A2(n_171),
.B(n_153),
.C(n_161),
.Y(n_189)
);

NOR2x1_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_166),
.Y(n_192)
);

INVxp33_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_10),
.C(n_13),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_192),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_183),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_195),
.C(n_14),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_186),
.A2(n_153),
.B1(n_11),
.B2(n_13),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_196),
.B(n_191),
.C(n_190),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_194),
.B(n_193),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_198),
.C(n_199),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_200),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_15),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_192),
.C(n_196),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_204),
.Y(n_205)
);


endmodule