module real_jpeg_16969_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_286;
wire n_166;
wire n_176;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AND2x2_ASAP7_75t_L g55 ( 
.A(n_0),
.B(n_56),
.Y(n_55)
);

AND2x4_ASAP7_75t_SL g80 ( 
.A(n_0),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_0),
.B(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g149 ( 
.A(n_0),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_0),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_1),
.B(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_1),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_1),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_1),
.B(n_121),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_1),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_1),
.B(n_224),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_1),
.B(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_2),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_3),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g158 ( 
.A(n_3),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_3),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_4),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_4),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_4),
.B(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_4),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_4),
.B(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_4),
.B(n_228),
.Y(n_227)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_5),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_5),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_6),
.B(n_33),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_6),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_7),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_7),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_7),
.Y(n_118)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_7),
.Y(n_163)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_7),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_8),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_8),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_8),
.B(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_8),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_8),
.B(n_210),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_8),
.B(n_150),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_8),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_8),
.B(n_323),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_9),
.B(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_9),
.A2(n_15),
.B1(n_36),
.B2(n_39),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_9),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_9),
.B(n_187),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_9),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_10),
.Y(n_102)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_10),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_11),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_11),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_11),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_11),
.B(n_50),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_11),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_11),
.B(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_11),
.B(n_359),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_12),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_13),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_13),
.B(n_68),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_14),
.Y(n_226)
);

BUFx4f_ASAP7_75t_L g363 ( 
.A(n_14),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_15),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_15),
.B(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_15),
.B(n_153),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_15),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_15),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_15),
.B(n_298),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_15),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_15),
.B(n_340),
.Y(n_339)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_16),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_215),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_213),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_170),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_20),
.B(n_170),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_92),
.C(n_135),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_21),
.A2(n_22),
.B1(n_92),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_57),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_23),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_34),
.C(n_43),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_24),
.B(n_277),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_27),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_25),
.B(n_28),
.C(n_32),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_30),
.B(n_194),
.Y(n_193)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_31),
.Y(n_132)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_31),
.Y(n_147)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_31),
.Y(n_310)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_33),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_34),
.A2(n_35),
.B1(n_43),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_35),
.A2(n_237),
.B(n_243),
.Y(n_236)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_42),
.Y(n_207)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_42),
.Y(n_268)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_43),
.Y(n_278)
);

MAJx2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_49),
.C(n_55),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_44),
.A2(n_45),
.B1(n_55),
.B2(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_44),
.A2(n_45),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_49),
.B(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_55),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_70),
.B1(n_90),
.B2(n_91),
.Y(n_57)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

MAJx2_ASAP7_75t_L g199 ( 
.A(n_59),
.B(n_67),
.C(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_66),
.B2(n_67),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_62),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_62),
.B(n_222),
.C(n_232),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_62),
.A2(n_232),
.B1(n_233),
.B2(n_380),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_62),
.Y(n_380)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVxp67_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_69),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g91 ( 
.A(n_70),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_70),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_79),
.C(n_84),
.Y(n_70)
);

XOR2x2_ASAP7_75t_SL g164 ( 
.A(n_71),
.B(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_74),
.C(n_77),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_72),
.A2(n_77),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_72),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_72),
.B(n_295),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_74),
.B(n_250),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_76),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_77),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_79),
.A2(n_80),
.B1(n_84),
.B2(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_81),
.Y(n_354)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_84),
.Y(n_166)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_88),
.Y(n_242)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_90),
.Y(n_174)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_92),
.Y(n_286)
);

XNOR2x2_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_107),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_93),
.B(n_108),
.C(n_123),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_97),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_94),
.B(n_98),
.C(n_103),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_103),
.Y(n_97)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_106),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_123),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_114),
.C(n_119),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_109),
.A2(n_119),
.B1(n_120),
.B2(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_109),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_112),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_114),
.B(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_119),
.B(n_261),
.C(n_265),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_119),
.A2(n_120),
.B1(n_265),
.B2(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_124),
.B(n_130),
.C(n_133),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_133),
.B2(n_134),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_133),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_133),
.A2(n_134),
.B1(n_193),
.B2(n_195),
.Y(n_192)
);

INVxp33_ASAP7_75t_SL g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_136),
.B(n_285),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_164),
.C(n_167),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_137),
.B(n_280),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.C(n_151),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2x2_ASAP7_75t_L g271 ( 
.A(n_139),
.B(n_272),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_143),
.B(n_151),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_149),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_144),
.B(n_149),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_157),
.C(n_159),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_152),
.A2(n_157),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_152),
.Y(n_257)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_157),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_157),
.A2(n_258),
.B1(n_345),
.B2(n_346),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_157),
.B(n_345),
.C(n_348),
.Y(n_370)
);

XOR2x1_ASAP7_75t_L g255 ( 
.A(n_159),
.B(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_164),
.B(n_167),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.C(n_174),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_196),
.B1(n_211),
.B2(n_212),
.Y(n_175)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_176),
.Y(n_212)
);

XOR2x2_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_190),
.Y(n_176)
);

XNOR2x1_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

XNOR2x2_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_186),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_188),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_189),
.Y(n_264)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_193),
.Y(n_195)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

XNOR2x1_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_208),
.B2(n_209),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_287),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_281),
.C(n_283),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_273),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_219),
.B(n_273),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_253),
.C(n_271),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_220),
.B(n_390),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_235),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_221),
.B(n_236),
.C(n_249),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_222),
.B(n_379),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_227),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_223),
.B(n_227),
.Y(n_321)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_223),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_223),
.A2(n_338),
.B1(n_339),
.B2(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_226),
.Y(n_305)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_230),
.Y(n_248)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_230),
.Y(n_341)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_249),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_251),
.B(n_296),
.C(n_297),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_254),
.B(n_271),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_259),
.C(n_269),
.Y(n_254)
);

XOR2x1_ASAP7_75t_L g384 ( 
.A(n_255),
.B(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_260),
.B(n_270),
.Y(n_385)
);

XOR2x1_ASAP7_75t_L g331 ( 
.A(n_261),
.B(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_265),
.Y(n_333)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_279),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_276),
.C(n_279),
.Y(n_282)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_282),
.B(n_284),
.Y(n_393)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NAND3xp33_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_289),
.C(n_393),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_388),
.B(n_392),
.Y(n_289)
);

AOI21x1_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_373),
.B(n_387),
.Y(n_290)
);

OAI21x1_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_334),
.B(n_372),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_317),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_293),
.B(n_317),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_299),
.C(n_307),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_294),
.B(n_368),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_299),
.A2(n_300),
.B1(n_307),
.B2(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_306),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_301),
.B(n_306),
.Y(n_349)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_307),
.Y(n_369)
);

AO22x1_ASAP7_75t_SL g307 ( 
.A1(n_308),
.A2(n_311),
.B1(n_315),
.B2(n_316),
.Y(n_307)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_308),
.Y(n_315)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_311),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_315),
.Y(n_319)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_316),
.B(n_358),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_329),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_318),
.B(n_330),
.C(n_331),
.Y(n_386)
);

XOR2x1_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

MAJx2_ASAP7_75t_L g382 ( 
.A(n_319),
.B(n_321),
.C(n_322),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx6_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

AOI21x1_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_366),
.B(n_371),
.Y(n_334)
);

OAI21x1_ASAP7_75t_SL g335 ( 
.A1(n_336),
.A2(n_350),
.B(n_365),
.Y(n_335)
);

NOR2x1_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_342),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_337),
.B(n_342),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_339),
.Y(n_356)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_343),
.A2(n_344),
.B1(n_348),
.B2(n_349),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

AOI21x1_ASAP7_75t_SL g350 ( 
.A1(n_351),
.A2(n_357),
.B(n_364),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_355),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_352),
.B(n_355),
.Y(n_364)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_367),
.B(n_370),
.Y(n_366)
);

NOR2x1_ASAP7_75t_SL g371 ( 
.A(n_367),
.B(n_370),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_374),
.B(n_386),
.Y(n_373)
);

NOR2x1_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_386),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_375),
.A2(n_376),
.B1(n_383),
.B2(n_384),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_376),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_377),
.A2(n_378),
.B1(n_381),
.B2(n_382),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_377),
.B(n_382),
.C(n_383),
.Y(n_391)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

NOR2xp67_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_391),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_389),
.B(n_391),
.Y(n_392)
);


endmodule