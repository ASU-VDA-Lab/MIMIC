module fake_jpeg_11596_n_143 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_143);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_20),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_26),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx4f_ASAP7_75t_SL g53 ( 
.A(n_37),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_5),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_46),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_60),
.A2(n_52),
.B1(n_41),
.B2(n_47),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_57),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_56),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_70),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_48),
.Y(n_70)
);

CKINVDCx6p67_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_71),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_60),
.B1(n_55),
.B2(n_49),
.Y(n_83)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_73),
.A2(n_41),
.B1(n_55),
.B2(n_47),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_82),
.A2(n_83),
.B(n_95),
.Y(n_110)
);

NOR2x1_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_53),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_89),
.Y(n_100)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_69),
.B(n_42),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_93),
.C(n_97),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_71),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_98),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_79),
.A2(n_49),
.B1(n_51),
.B2(n_54),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_92),
.A2(n_94),
.B1(n_8),
.B2(n_9),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_40),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_44),
.B1(n_40),
.B2(n_4),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_76),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_95)
);

AND2x6_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_23),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_72),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_101),
.B(n_106),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_6),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_104),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_7),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_8),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_88),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_107),
.B(n_113),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_112),
.Y(n_126)
);

AND2x4_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_25),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_109),
.A2(n_28),
.B(n_29),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_82),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_109),
.B1(n_114),
.B2(n_110),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_12),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_85),
.B(n_14),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_82),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_114),
.A2(n_18),
.B1(n_21),
.B2(n_24),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_123),
.Y(n_131)
);

NAND2x1_ASAP7_75t_SL g127 ( 
.A(n_117),
.B(n_125),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_30),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_119),
.B(n_121),
.Y(n_128)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_31),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_103),
.Y(n_123)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_32),
.C(n_33),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_122),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_130),
.A2(n_115),
.B1(n_118),
.B2(n_126),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_133),
.B(n_134),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_124),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_129),
.A2(n_117),
.B1(n_109),
.B2(n_125),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_135),
.A2(n_128),
.B(n_131),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_134),
.Y(n_138)
);

A2O1A1O1Ixp25_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_137),
.B(n_129),
.C(n_127),
.D(n_39),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_140),
.B(n_36),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_127),
.Y(n_143)
);


endmodule