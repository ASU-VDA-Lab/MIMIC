module fake_ariane_3179_n_4335 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_332, n_294, n_197, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_57, n_424, n_387, n_406, n_117, n_139, n_85, n_130, n_349, n_391, n_346, n_214, n_348, n_2, n_32, n_410, n_379, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_267, n_335, n_350, n_291, n_344, n_381, n_426, n_398, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_390, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_413, n_392, n_376, n_221, n_321, n_86, n_361, n_89, n_149, n_383, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_409, n_171, n_384, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_418, n_223, n_403, n_25, n_83, n_389, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_378, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_428, n_159, n_358, n_105, n_30, n_131, n_263, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_425, n_118, n_121, n_411, n_353, n_22, n_241, n_29, n_357, n_412, n_191, n_382, n_80, n_211, n_97, n_408, n_322, n_251, n_116, n_397, n_351, n_39, n_393, n_359, n_155, n_127, n_4335);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_57;
input n_424;
input n_387;
input n_406;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_391;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_410;
input n_379;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_398;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_413;
input n_392;
input n_376;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_409;
input n_171;
input n_384;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_418;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_378;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_425;
input n_118;
input n_121;
input n_411;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_191;
input n_382;
input n_80;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_116;
input n_397;
input n_351;
input n_39;
input n_393;
input n_359;
input n_155;
input n_127;

output n_4335;

wire n_2752;
wire n_3527;
wire n_913;
wire n_1681;
wire n_2163;
wire n_3432;
wire n_4030;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_3619;
wire n_589;
wire n_2484;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_4013;
wire n_3152;
wire n_2346;
wire n_3434;
wire n_1469;
wire n_691;
wire n_1353;
wire n_3056;
wire n_3500;
wire n_3480;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_3268;
wire n_3853;
wire n_2559;
wire n_4213;
wire n_4127;
wire n_2500;
wire n_2509;
wire n_4085;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_4259;
wire n_3264;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_3181;
wire n_850;
wire n_2993;
wire n_4299;
wire n_4283;
wire n_1916;
wire n_2879;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2818;
wire n_2407;
wire n_690;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_1430;
wire n_525;
wire n_3745;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_3487;
wire n_1238;
wire n_2694;
wire n_3668;
wire n_2011;
wire n_3742;
wire n_2729;
wire n_4302;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_4178;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_717;
wire n_3765;
wire n_2006;
wire n_4090;
wire n_952;
wire n_864;
wire n_4058;
wire n_2446;
wire n_1096;
wire n_4116;
wire n_1379;
wire n_2436;
wire n_3352;
wire n_3517;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2702;
wire n_2461;
wire n_3719;
wire n_524;
wire n_2731;
wire n_3703;
wire n_634;
wire n_1214;
wire n_3561;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_3526;
wire n_3888;
wire n_3954;
wire n_2042;
wire n_2123;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_4103;
wire n_1196;
wire n_462;
wire n_1181;
wire n_1999;
wire n_3435;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_3154;
wire n_2646;
wire n_1298;
wire n_737;
wire n_2653;
wire n_2873;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_3115;
wire n_3938;
wire n_568;
wire n_2278;
wire n_4028;
wire n_3330;
wire n_3514;
wire n_1088;
wire n_1424;
wire n_766;
wire n_2976;
wire n_1835;
wire n_3383;
wire n_3965;
wire n_1457;
wire n_2482;
wire n_3905;
wire n_1682;
wire n_2750;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_520;
wire n_870;
wire n_2547;
wire n_3382;
wire n_1453;
wire n_945;
wire n_958;
wire n_3943;
wire n_3930;
wire n_2554;
wire n_3145;
wire n_3808;
wire n_2248;
wire n_3665;
wire n_3063;
wire n_4321;
wire n_813;
wire n_3281;
wire n_3535;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_3081;
wire n_3858;
wire n_4106;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_3220;
wire n_2960;
wire n_500;
wire n_754;
wire n_665;
wire n_4260;
wire n_903;
wire n_3270;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_3348;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_3261;
wire n_829;
wire n_1761;
wire n_4148;
wire n_1062;
wire n_738;
wire n_3679;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_3283;
wire n_4038;
wire n_4132;
wire n_3856;
wire n_2442;
wire n_2735;
wire n_4159;
wire n_953;
wire n_1364;
wire n_4214;
wire n_2390;
wire n_4331;
wire n_1888;
wire n_1224;
wire n_3657;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_3451;
wire n_625;
wire n_557;
wire n_2322;
wire n_2746;
wire n_3419;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_2370;
wire n_559;
wire n_2663;
wire n_2233;
wire n_495;
wire n_2914;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_3545;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_2878;
wire n_1284;
wire n_1428;
wire n_1241;
wire n_3890;
wire n_3830;
wire n_821;
wire n_561;
wire n_770;
wire n_3252;
wire n_1514;
wire n_4143;
wire n_4273;
wire n_2539;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_2782;
wire n_3879;
wire n_569;
wire n_4136;
wire n_2078;
wire n_3315;
wire n_3929;
wire n_1145;
wire n_3523;
wire n_971;
wire n_3144;
wire n_2359;
wire n_3999;
wire n_2201;
wire n_787;
wire n_4012;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_4176;
wire n_1207;
wire n_4124;
wire n_3606;
wire n_786;
wire n_1404;
wire n_3347;
wire n_3420;
wire n_3859;
wire n_868;
wire n_3474;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_4320;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_3150;
wire n_2950;
wire n_1542;
wire n_3552;
wire n_1314;
wire n_3756;
wire n_3639;
wire n_3254;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_3121;
wire n_2847;
wire n_884;
wire n_3412;
wire n_4077;
wire n_1851;
wire n_2162;
wire n_3209;
wire n_3324;
wire n_3015;
wire n_1415;
wire n_3870;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_3749;
wire n_1085;
wire n_2988;
wire n_1636;
wire n_3482;
wire n_432;
wire n_823;
wire n_1900;
wire n_620;
wire n_3948;
wire n_1074;
wire n_3230;
wire n_859;
wire n_3793;
wire n_4268;
wire n_1765;
wire n_4031;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_1254;
wire n_3960;
wire n_4147;
wire n_929;
wire n_3207;
wire n_3641;
wire n_2433;
wire n_899;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_3828;
wire n_3975;
wire n_3073;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_3183;
wire n_3571;
wire n_1013;
wire n_3883;
wire n_4032;
wire n_4018;
wire n_1495;
wire n_3607;
wire n_1637;
wire n_3297;
wire n_2571;
wire n_2427;
wire n_3325;
wire n_3613;
wire n_2885;
wire n_661;
wire n_2098;
wire n_4227;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_3003;
wire n_4117;
wire n_533;
wire n_3049;
wire n_3136;
wire n_2867;
wire n_3634;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_3066;
wire n_1811;
wire n_2045;
wire n_3274;
wire n_3877;
wire n_4284;
wire n_440;
wire n_3913;
wire n_3817;
wire n_3013;
wire n_3612;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_3739;
wire n_1230;
wire n_612;
wire n_1840;
wire n_2739;
wire n_3728;
wire n_3962;
wire n_512;
wire n_1597;
wire n_4082;
wire n_2942;
wire n_1771;
wire n_2902;
wire n_1544;
wire n_579;
wire n_3271;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_3164;
wire n_2094;
wire n_3854;
wire n_3861;
wire n_2956;
wire n_1354;
wire n_1790;
wire n_2512;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_4171;
wire n_3652;
wire n_3449;
wire n_2788;
wire n_4119;
wire n_1021;
wire n_1443;
wire n_4000;
wire n_3089;
wire n_491;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_3084;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_3458;
wire n_570;
wire n_2727;
wire n_942;
wire n_3580;
wire n_1437;
wire n_3860;
wire n_3511;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_461;
wire n_1416;
wire n_2909;
wire n_490;
wire n_3554;
wire n_1461;
wire n_2717;
wire n_3012;
wire n_1391;
wire n_2981;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_3850;
wire n_575;
wire n_546;
wire n_3472;
wire n_503;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_700;
wire n_772;
wire n_1216;
wire n_4174;
wire n_3126;
wire n_3754;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_676;
wire n_3758;
wire n_2038;
wire n_2263;
wire n_3518;
wire n_3958;
wire n_2800;
wire n_2568;
wire n_2271;
wire n_2116;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_3485;
wire n_1594;
wire n_680;
wire n_1935;
wire n_2806;
wire n_3191;
wire n_1716;
wire n_4109;
wire n_3777;
wire n_4108;
wire n_1872;
wire n_3562;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_3359;
wire n_3767;
wire n_3841;
wire n_3119;
wire n_1108;
wire n_3588;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_3234;
wire n_3280;
wire n_3413;
wire n_3692;
wire n_3900;
wire n_2216;
wire n_4115;
wire n_1274;
wire n_3539;
wire n_2426;
wire n_652;
wire n_1819;
wire n_475;
wire n_3095;
wire n_947;
wire n_2134;
wire n_3862;
wire n_1260;
wire n_930;
wire n_3698;
wire n_3716;
wire n_4226;
wire n_1179;
wire n_468;
wire n_3284;
wire n_3909;
wire n_4311;
wire n_4220;
wire n_2703;
wire n_2926;
wire n_1442;
wire n_696;
wire n_482;
wire n_2620;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_3391;
wire n_3506;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_2549;
wire n_2499;
wire n_3678;
wire n_762;
wire n_1253;
wire n_1661;
wire n_1468;
wire n_2791;
wire n_555;
wire n_2683;
wire n_3212;
wire n_804;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_3529;
wire n_4180;
wire n_2970;
wire n_4235;
wire n_3159;
wire n_966;
wire n_992;
wire n_955;
wire n_3549;
wire n_3885;
wire n_3914;
wire n_3624;
wire n_4264;
wire n_1182;
wire n_794;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_3192;
wire n_2611;
wire n_1562;
wire n_514;
wire n_2748;
wire n_2185;
wire n_3306;
wire n_3250;
wire n_4223;
wire n_3029;
wire n_2398;
wire n_4233;
wire n_3538;
wire n_3915;
wire n_1376;
wire n_3839;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2925;
wire n_2015;
wire n_1435;
wire n_3407;
wire n_3717;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_3460;
wire n_3544;
wire n_1610;
wire n_3875;
wire n_4029;
wire n_2202;
wire n_2072;
wire n_3852;
wire n_2952;
wire n_3530;
wire n_4206;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_4099;
wire n_3120;
wire n_2922;
wire n_436;
wire n_3000;
wire n_2871;
wire n_2930;
wire n_3193;
wire n_3240;
wire n_2745;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_2628;
wire n_3219;
wire n_3362;
wire n_619;
wire n_967;
wire n_437;
wire n_1083;
wire n_4130;
wire n_3937;
wire n_2161;
wire n_1418;
wire n_4175;
wire n_746;
wire n_1357;
wire n_1079;
wire n_4170;
wire n_1787;
wire n_2462;
wire n_3510;
wire n_1389;
wire n_3393;
wire n_3172;
wire n_2155;
wire n_2659;
wire n_4033;
wire n_615;
wire n_3747;
wire n_1139;
wire n_2836;
wire n_3688;
wire n_2439;
wire n_2864;
wire n_517;
wire n_1312;
wire n_1717;
wire n_3604;
wire n_4045;
wire n_1812;
wire n_3651;
wire n_824;
wire n_2172;
wire n_2601;
wire n_3614;
wire n_3871;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_3757;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_4272;
wire n_2219;
wire n_3116;
wire n_4141;
wire n_1855;
wire n_3784;
wire n_2100;
wire n_2333;
wire n_3176;
wire n_3629;
wire n_3666;
wire n_3372;
wire n_3891;
wire n_990;
wire n_1623;
wire n_3559;
wire n_1903;
wire n_3792;
wire n_867;
wire n_2147;
wire n_4267;
wire n_3479;
wire n_4020;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_3998;
wire n_3724;
wire n_4150;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_3287;
wire n_2167;
wire n_4285;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_470;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_3046;
wire n_1087;
wire n_4055;
wire n_3980;
wire n_2701;
wire n_3021;
wire n_2400;
wire n_632;
wire n_3257;
wire n_477;
wire n_650;
wire n_3741;
wire n_2388;
wire n_3730;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_1911;
wire n_3979;
wire n_3912;
wire n_2567;
wire n_3950;
wire n_3496;
wire n_3493;
wire n_2557;
wire n_2695;
wire n_2898;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_3727;
wire n_3700;
wire n_976;
wire n_712;
wire n_3567;
wire n_909;
wire n_4003;
wire n_1392;
wire n_767;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_4307;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_3014;
wire n_489;
wire n_2294;
wire n_2274;
wire n_3342;
wire n_2895;
wire n_2903;
wire n_974;
wire n_506;
wire n_3814;
wire n_3812;
wire n_3127;
wire n_3796;
wire n_1731;
wire n_799;
wire n_3884;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_3625;
wire n_2467;
wire n_3375;
wire n_2768;
wire n_471;
wire n_965;
wire n_1914;
wire n_4195;
wire n_3760;
wire n_2253;
wire n_934;
wire n_2213;
wire n_3515;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_4056;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_3010;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_3744;
wire n_4015;
wire n_2924;
wire n_1209;
wire n_4022;
wire n_1020;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_646;
wire n_4254;
wire n_2507;
wire n_4219;
wire n_3438;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_2896;
wire n_1913;
wire n_2495;
wire n_2069;
wire n_3187;
wire n_1058;
wire n_2328;
wire n_4043;
wire n_2434;
wire n_1042;
wire n_3170;
wire n_1234;
wire n_2311;
wire n_479;
wire n_3936;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_3147;
wire n_2287;
wire n_836;
wire n_2223;
wire n_3082;
wire n_1279;
wire n_3415;
wire n_3661;
wire n_2473;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_2511;
wire n_3464;
wire n_564;
wire n_3414;
wire n_1029;
wire n_2649;
wire n_3981;
wire n_1247;
wire n_4234;
wire n_760;
wire n_522;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_3210;
wire n_1483;
wire n_3108;
wire n_1363;
wire n_2681;
wire n_3867;
wire n_3397;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_3467;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_598;
wire n_3031;
wire n_2262;
wire n_3179;
wire n_2565;
wire n_3889;
wire n_1237;
wire n_3262;
wire n_4314;
wire n_927;
wire n_1095;
wire n_2980;
wire n_1728;
wire n_2335;
wire n_3078;
wire n_3699;
wire n_3971;
wire n_4315;
wire n_706;
wire n_2120;
wire n_3239;
wire n_2631;
wire n_3215;
wire n_3311;
wire n_3869;
wire n_3516;
wire n_1401;
wire n_1419;
wire n_3138;
wire n_1531;
wire n_776;
wire n_2860;
wire n_3816;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_3528;
wire n_1651;
wire n_3087;
wire n_2697;
wire n_1387;
wire n_466;
wire n_1263;
wire n_1817;
wire n_3711;
wire n_4207;
wire n_4201;
wire n_2404;
wire n_2757;
wire n_2168;
wire n_3704;
wire n_552;
wire n_2312;
wire n_670;
wire n_2677;
wire n_4296;
wire n_1826;
wire n_3171;
wire n_3577;
wire n_2834;
wire n_4051;
wire n_2483;
wire n_4242;
wire n_4074;
wire n_3994;
wire n_441;
wire n_1951;
wire n_3185;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_2996;
wire n_637;
wire n_1592;
wire n_2812;
wire n_3660;
wire n_2662;
wire n_1259;
wire n_3300;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_3104;
wire n_3074;
wire n_2655;
wire n_1231;
wire n_3917;
wire n_4122;
wire n_3246;
wire n_2132;
wire n_3299;
wire n_980;
wire n_1618;
wire n_4275;
wire n_3774;
wire n_1869;
wire n_3589;
wire n_3623;
wire n_1743;
wire n_905;
wire n_2718;
wire n_4263;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_3876;
wire n_3615;
wire n_3267;
wire n_1802;
wire n_2178;
wire n_3946;
wire n_4243;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_3054;
wire n_2811;
wire n_3019;
wire n_1795;
wire n_3200;
wire n_1384;
wire n_4225;
wire n_3642;
wire n_2237;
wire n_4153;
wire n_2146;
wire n_4274;
wire n_2983;
wire n_1868;
wire n_3276;
wire n_3601;
wire n_4089;
wire n_1501;
wire n_4186;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_3513;
wire n_3498;
wire n_3682;
wire n_2350;
wire n_3881;
wire n_1068;
wire n_1198;
wire n_4096;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_3759;
wire n_3377;
wire n_487;
wire n_1518;
wire n_3323;
wire n_1456;
wire n_4007;
wire n_1879;
wire n_1886;
wire n_4138;
wire n_1648;
wire n_2187;
wire n_3961;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_3863;
wire n_2129;
wire n_855;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_808;
wire n_1365;
wire n_2476;
wire n_553;
wire n_2814;
wire n_2059;
wire n_3675;
wire n_3968;
wire n_4133;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_578;
wire n_3466;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_3572;
wire n_2975;
wire n_3332;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_3374;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2998;
wire n_3465;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_3118;
wire n_4072;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_4323;
wire n_529;
wire n_1899;
wire n_3039;
wire n_2195;
wire n_3922;
wire n_502;
wire n_2194;
wire n_2937;
wire n_4293;
wire n_3508;
wire n_1467;
wire n_4039;
wire n_1828;
wire n_4129;
wire n_2159;
wire n_1798;
wire n_3057;
wire n_1304;
wire n_1608;
wire n_3831;
wire n_1744;
wire n_3335;
wire n_3007;
wire n_2267;
wire n_1105;
wire n_547;
wire n_3599;
wire n_3618;
wire n_604;
wire n_439;
wire n_677;
wire n_3705;
wire n_3022;
wire n_478;
wire n_703;
wire n_3983;
wire n_1349;
wire n_1709;
wire n_3318;
wire n_1061;
wire n_3385;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_681;
wire n_3286;
wire n_3734;
wire n_3370;
wire n_874;
wire n_3773;
wire n_3949;
wire n_2286;
wire n_3494;
wire n_2023;
wire n_1278;
wire n_4247;
wire n_707;
wire n_3974;
wire n_3443;
wire n_3401;
wire n_983;
wire n_3036;
wire n_2783;
wire n_2599;
wire n_3988;
wire n_3788;
wire n_3939;
wire n_699;
wire n_727;
wire n_590;
wire n_1726;
wire n_2075;
wire n_3263;
wire n_3542;
wire n_2523;
wire n_1945;
wire n_3569;
wire n_3837;
wire n_3835;
wire n_545;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2496;
wire n_3260;
wire n_3349;
wire n_3819;
wire n_3761;
wire n_3996;
wire n_4292;
wire n_2118;
wire n_3222;
wire n_1740;
wire n_1602;
wire n_688;
wire n_3139;
wire n_636;
wire n_2853;
wire n_3350;
wire n_3801;
wire n_1098;
wire n_3009;
wire n_1490;
wire n_2338;
wire n_442;
wire n_777;
wire n_3764;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_3025;
wire n_3636;
wire n_3051;
wire n_3205;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_3653;
wire n_3951;
wire n_3868;
wire n_3035;
wire n_3823;
wire n_729;
wire n_887;
wire n_3403;
wire n_4261;
wire n_2218;
wire n_2057;
wire n_1122;
wire n_1408;
wire n_1205;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_501;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2944;
wire n_2861;
wire n_4236;
wire n_2780;
wire n_3023;
wire n_1120;
wire n_3439;
wire n_3942;
wire n_1202;
wire n_4084;
wire n_627;
wire n_2254;
wire n_3130;
wire n_3290;
wire n_1498;
wire n_1188;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_2618;
wire n_4121;
wire n_3602;
wire n_4216;
wire n_957;
wire n_1402;
wire n_1242;
wire n_3957;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_3418;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_3611;
wire n_3781;
wire n_2217;
wire n_2226;
wire n_3959;
wire n_3984;
wire n_1586;
wire n_4313;
wire n_861;
wire n_3338;
wire n_2962;
wire n_1543;
wire n_1431;
wire n_877;
wire n_3995;
wire n_1119;
wire n_3713;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_3908;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_2763;
wire n_4297;
wire n_4229;
wire n_3156;
wire n_2256;
wire n_1189;
wire n_3337;
wire n_1089;
wire n_3750;
wire n_3424;
wire n_3326;
wire n_3356;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_1502;
wire n_3044;
wire n_1523;
wire n_2190;
wire n_3501;
wire n_3492;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_3737;
wire n_2516;
wire n_3931;
wire n_4094;
wire n_2776;
wire n_2555;
wire n_3216;
wire n_3224;
wire n_3568;
wire n_1969;
wire n_2708;
wire n_735;
wire n_3070;
wire n_1005;
wire n_3275;
wire n_527;
wire n_2379;
wire n_3579;
wire n_3245;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_845;
wire n_888;
wire n_2949;
wire n_2894;
wire n_2300;
wire n_4049;
wire n_4067;
wire n_3896;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_4182;
wire n_4269;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_3214;
wire n_551;
wire n_3551;
wire n_1708;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_1222;
wire n_2284;
wire n_3005;
wire n_3710;
wire n_1844;
wire n_2283;
wire n_582;
wire n_2526;
wire n_1957;
wire n_3364;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_3803;
wire n_3766;
wire n_3985;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_2994;
wire n_534;
wire n_1791;
wire n_2508;
wire n_3186;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_3826;
wire n_2266;
wire n_3944;
wire n_3417;
wire n_2449;
wire n_560;
wire n_890;
wire n_4324;
wire n_842;
wire n_3626;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_3180;
wire n_3648;
wire n_3423;
wire n_742;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2742;
wire n_2119;
wire n_769;
wire n_3671;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_2821;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_3696;
wire n_2474;
wire n_4104;
wire n_2623;
wire n_3392;
wire n_982;
wire n_1800;
wire n_915;
wire n_3791;
wire n_1075;
wire n_2008;
wire n_454;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_3064;
wire n_3199;
wire n_4034;
wire n_1529;
wire n_4228;
wire n_3353;
wire n_1227;
wire n_3531;
wire n_2127;
wire n_655;
wire n_2946;
wire n_3166;
wire n_4237;
wire n_3151;
wire n_3649;
wire n_3684;
wire n_3333;
wire n_3512;
wire n_1734;
wire n_1860;
wire n_3065;
wire n_3016;
wire n_4114;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_3135;
wire n_657;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_3924;
wire n_4081;
wire n_837;
wire n_812;
wire n_2448;
wire n_3997;
wire n_2211;
wire n_4172;
wire n_4040;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_3024;
wire n_2772;
wire n_3564;
wire n_862;
wire n_1700;
wire n_2637;
wire n_659;
wire n_1332;
wire n_3795;
wire n_2306;
wire n_509;
wire n_4328;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_3990;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_3953;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_2893;
wire n_1532;
wire n_3277;
wire n_1171;
wire n_1030;
wire n_785;
wire n_3208;
wire n_3161;
wire n_2389;
wire n_4069;
wire n_1309;
wire n_3582;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_4280;
wire n_456;
wire n_1867;
wire n_3993;
wire n_852;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_3459;
wire n_3617;
wire n_704;
wire n_2958;
wire n_3365;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_4113;
wire n_2696;
wire n_3340;
wire n_4192;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_3977;
wire n_1400;
wire n_4112;
wire n_3400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_3735;
wire n_3486;
wire n_1513;
wire n_1527;
wire n_2581;
wire n_1783;
wire n_3656;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_3069;
wire n_2992;
wire n_4221;
wire n_1037;
wire n_3650;
wire n_4071;
wire n_1329;
wire n_3197;
wire n_1993;
wire n_1545;
wire n_3586;
wire n_2629;
wire n_3369;
wire n_4035;
wire n_4160;
wire n_3256;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_3670;
wire n_1668;
wire n_1878;
wire n_3964;
wire n_2540;
wire n_3836;
wire n_4190;
wire n_3302;
wire n_1605;
wire n_4137;
wire n_1078;
wire n_3060;
wire n_2486;
wire n_1897;
wire n_2984;
wire n_4009;
wire n_3646;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_3685;
wire n_811;
wire n_4145;
wire n_3097;
wire n_624;
wire n_3507;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_2492;
wire n_3864;
wire n_2939;
wire n_3425;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_3450;
wire n_3748;
wire n_2337;
wire n_2265;
wire n_687;
wire n_2900;
wire n_797;
wire n_2026;
wire n_2912;
wire n_3524;
wire n_1786;
wire n_2627;
wire n_4050;
wire n_3173;
wire n_480;
wire n_1327;
wire n_3732;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_595;
wire n_4306;
wire n_1405;
wire n_2684;
wire n_3174;
wire n_3314;
wire n_2726;
wire n_602;
wire n_3813;
wire n_2622;
wire n_3447;
wire n_4006;
wire n_2272;
wire n_3266;
wire n_1757;
wire n_592;
wire n_3102;
wire n_1499;
wire n_854;
wire n_1318;
wire n_4288;
wire n_3452;
wire n_2091;
wire n_1769;
wire n_1632;
wire n_474;
wire n_1929;
wire n_4098;
wire n_4312;
wire n_1950;
wire n_2691;
wire n_2264;
wire n_3789;
wire n_805;
wire n_4319;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_3124;
wire n_3811;
wire n_3422;
wire n_1658;
wire n_4200;
wire n_2249;
wire n_1072;
wire n_3411;
wire n_695;
wire n_1526;
wire n_2991;
wire n_3463;
wire n_1305;
wire n_2785;
wire n_730;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_516;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_4289;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1856;
wire n_1733;
wire n_2016;
wire n_2667;
wire n_2723;
wire n_1524;
wire n_2725;
wire n_3925;
wire n_2928;
wire n_943;
wire n_1118;
wire n_678;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_651;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_3167;
wire n_3746;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_3780;
wire n_1657;
wire n_878;
wire n_2857;
wire n_3694;
wire n_4118;
wire n_1784;
wire n_3110;
wire n_3857;
wire n_771;
wire n_3787;
wire n_4025;
wire n_4239;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_3157;
wire n_3893;
wire n_3753;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_3702;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_4076;
wire n_806;
wire n_3142;
wire n_1984;
wire n_1350;
wire n_3453;
wire n_3129;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_2720;
wire n_3298;
wire n_3107;
wire n_3495;
wire n_1352;
wire n_3843;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_4065;
wire n_2383;
wire n_2764;
wire n_1822;
wire n_1441;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_3708;
wire n_819;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_2945;
wire n_586;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_3543;
wire n_3640;
wire n_1776;
wire n_3448;
wire n_686;
wire n_4279;
wire n_605;
wire n_2936;
wire n_1154;
wire n_584;
wire n_3609;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_4330;
wire n_1130;
wire n_1450;
wire n_4152;
wire n_3718;
wire n_756;
wire n_2022;
wire n_3390;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_3740;
wire n_2986;
wire n_2320;
wire n_3017;
wire n_979;
wire n_2570;
wire n_2329;
wire n_3140;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_3976;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_2911;
wire n_2890;
wire n_515;
wire n_3381;
wire n_807;
wire n_3455;
wire n_3736;
wire n_891;
wire n_3313;
wire n_885;
wire n_1659;
wire n_3955;
wire n_2354;
wire n_3591;
wire n_1864;
wire n_2760;
wire n_3907;
wire n_3086;
wire n_4332;
wire n_1887;
wire n_3165;
wire n_1208;
wire n_4281;
wire n_3317;
wire n_3945;
wire n_3726;
wire n_3336;
wire n_1987;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_3635;
wire n_2352;
wire n_3541;
wire n_2502;
wire n_1256;
wire n_714;
wire n_3605;
wire n_3345;
wire n_2170;
wire n_3560;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_725;
wire n_2377;
wire n_1577;
wire n_3566;
wire n_3840;
wire n_3421;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_3548;
wire n_2652;
wire n_1133;
wire n_3067;
wire n_883;
wire n_4097;
wire n_4054;
wire n_3809;
wire n_4162;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_3169;
wire n_594;
wire n_3236;
wire n_2222;
wire n_3468;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_4173;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_4301;
wire n_3573;
wire n_2203;
wire n_2133;
wire n_2076;
wire n_833;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_3319;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_3321;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_3291;
wire n_3654;
wire n_4188;
wire n_2001;
wire n_1047;
wire n_3783;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_4008;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_4140;
wire n_1050;
wire n_2626;
wire n_566;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_3643;
wire n_2285;
wire n_3343;
wire n_3184;
wire n_3309;
wire n_2892;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_2796;
wire n_858;
wire n_2804;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_3982;
wire n_2715;
wire n_3206;
wire n_3647;
wire n_1035;
wire n_3475;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_433;
wire n_3973;
wire n_3134;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_3755;
wire n_2947;
wire n_1367;
wire n_3842;
wire n_4202;
wire n_2044;
wire n_928;
wire n_4304;
wire n_3886;
wire n_1153;
wire n_465;
wire n_3769;
wire n_4078;
wire n_825;
wire n_1103;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_3738;
wire n_894;
wire n_3098;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_3055;
wire n_1291;
wire n_562;
wire n_4070;
wire n_2020;
wire n_748;
wire n_3987;
wire n_2310;
wire n_510;
wire n_4249;
wire n_1045;
wire n_3341;
wire n_3600;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_4125;
wire n_1023;
wire n_2711;
wire n_3223;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_3386;
wire n_4139;
wire n_914;
wire n_689;
wire n_1116;
wire n_4327;
wire n_3921;
wire n_3043;
wire n_3190;
wire n_1958;
wire n_2747;
wire n_3667;
wire n_3027;
wire n_4011;
wire n_467;
wire n_1511;
wire n_2177;
wire n_3695;
wire n_2713;
wire n_1422;
wire n_3800;
wire n_2766;
wire n_1965;
wire n_644;
wire n_3462;
wire n_4196;
wire n_1197;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_2613;
wire n_3226;
wire n_497;
wire n_3733;
wire n_1165;
wire n_3378;
wire n_2934;
wire n_1641;
wire n_3967;
wire n_3731;
wire n_4291;
wire n_538;
wire n_2845;
wire n_4151;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_2647;
wire n_455;
wire n_429;
wire n_588;
wire n_3358;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_3920;
wire n_1307;
wire n_3444;
wire n_1128;
wire n_3141;
wire n_2053;
wire n_4091;
wire n_3851;
wire n_1671;
wire n_1417;
wire n_3476;
wire n_1048;
wire n_2343;
wire n_775;
wire n_3096;
wire n_667;
wire n_2419;
wire n_1049;
wire n_3380;
wire n_2330;
wire n_2826;
wire n_869;
wire n_4184;
wire n_846;
wire n_1398;
wire n_1921;
wire n_4166;
wire n_2777;
wire n_3238;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_3189;
wire n_3233;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_3175;
wire n_1440;
wire n_3289;
wire n_2666;
wire n_3322;
wire n_1370;
wire n_1603;
wire n_728;
wire n_4191;
wire n_2935;
wire n_2401;
wire n_4246;
wire n_715;
wire n_889;
wire n_3822;
wire n_3255;
wire n_3818;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2886;
wire n_3827;
wire n_2478;
wire n_685;
wire n_911;
wire n_4061;
wire n_2658;
wire n_623;
wire n_3509;
wire n_3587;
wire n_2608;
wire n_3620;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1948;
wire n_1534;
wire n_3006;
wire n_2767;
wire n_4155;
wire n_810;
wire n_3376;
wire n_4278;
wire n_1290;
wire n_1959;
wire n_3497;
wire n_617;
wire n_3770;
wire n_2396;
wire n_3243;
wire n_543;
wire n_3368;
wire n_1362;
wire n_4326;
wire n_1559;
wire n_2121;
wire n_3456;
wire n_3865;
wire n_3123;
wire n_2692;
wire n_601;
wire n_683;
wire n_565;
wire n_3927;
wire n_628;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_2068;
wire n_3117;
wire n_3595;
wire n_4308;
wire n_743;
wire n_1194;
wire n_2862;
wire n_4060;
wire n_1647;
wire n_1546;
wire n_3384;
wire n_4325;
wire n_1420;
wire n_2645;
wire n_2553;
wire n_3790;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_660;
wire n_464;
wire n_3490;
wire n_2459;
wire n_962;
wire n_941;
wire n_3396;
wire n_1210;
wire n_847;
wire n_747;
wire n_4241;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_3113;
wire n_4183;
wire n_3101;
wire n_918;
wire n_1968;
wire n_3307;
wire n_3662;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_3251;
wire n_3288;
wire n_4093;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_4123;
wire n_1038;
wire n_3603;
wire n_3723;
wire n_4135;
wire n_2371;
wire n_1978;
wire n_4257;
wire n_571;
wire n_4282;
wire n_4294;
wire n_3880;
wire n_3720;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_3683;
wire n_3904;
wire n_3887;
wire n_593;
wire n_3195;
wire n_3008;
wire n_1695;
wire n_3242;
wire n_4027;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_3405;
wire n_4309;
wire n_2313;
wire n_609;
wire n_3077;
wire n_1193;
wire n_3048;
wire n_3339;
wire n_1345;
wire n_613;
wire n_3037;
wire n_1022;
wire n_4126;
wire n_4164;
wire n_1336;
wire n_1033;
wire n_3478;
wire n_4333;
wire n_3062;
wire n_1774;
wire n_2963;
wire n_3532;
wire n_519;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_3363;
wire n_3533;
wire n_3978;
wire n_1767;
wire n_1040;
wire n_674;
wire n_3131;
wire n_1158;
wire n_3168;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_3409;
wire n_4079;
wire n_3522;
wire n_3583;
wire n_4088;
wire n_4316;
wire n_2882;
wire n_2303;
wire n_2669;
wire n_3540;
wire n_3911;
wire n_3241;
wire n_3802;
wire n_3899;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_3481;
wire n_629;
wire n_3563;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_1814;
wire n_4210;
wire n_532;
wire n_3689;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_4041;
wire n_2174;
wire n_2688;
wire n_540;
wire n_2624;
wire n_692;
wire n_3442;
wire n_4208;
wire n_3972;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_3926;
wire n_4209;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_4004;
wire n_1552;
wire n_750;
wire n_2938;
wire n_834;
wire n_3630;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_3992;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_2189;
wire n_621;
wire n_2648;
wire n_3305;
wire n_1587;
wire n_3810;
wire n_4062;
wire n_2093;
wire n_2340;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_3354;
wire n_1014;
wire n_724;
wire n_2204;
wire n_2931;
wire n_3433;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2977;
wire n_3106;
wire n_3597;
wire n_3991;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_3092;
wire n_3437;
wire n_2231;
wire n_3786;
wire n_697;
wire n_2828;
wire n_4212;
wire n_4270;
wire n_622;
wire n_1626;
wire n_3436;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_3806;
wire n_4204;
wire n_3553;
wire n_4044;
wire n_2305;
wire n_3645;
wire n_880;
wire n_793;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3304;
wire n_3833;
wire n_3574;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_3751;
wire n_3402;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_3247;
wire n_1621;
wire n_4110;
wire n_739;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_1221;
wire n_4217;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_4271;
wire n_2180;
wire n_1942;
wire n_3406;
wire n_4317;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_580;
wire n_3664;
wire n_1579;
wire n_494;
wire n_2809;
wire n_4218;
wire n_2181;
wire n_3550;
wire n_434;
wire n_2014;
wire n_975;
wire n_2974;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_2870;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_3686;
wire n_3722;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_3969;
wire n_1805;
wire n_2282;
wire n_3301;
wire n_981;
wire n_4068;
wire n_2910;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_3873;
wire n_2270;
wire n_3470;
wire n_4163;
wire n_3785;
wire n_3294;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_3610;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_3279;
wire n_994;
wire n_2428;
wire n_2972;
wire n_2586;
wire n_2989;
wire n_1360;
wire n_973;
wire n_3178;
wire n_2858;
wire n_972;
wire n_3844;
wire n_3259;
wire n_4262;
wire n_2251;
wire n_2923;
wire n_3076;
wire n_2843;
wire n_3714;
wire n_3410;
wire n_856;
wire n_3100;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_3721;
wire n_3677;
wire n_1564;
wire n_2010;
wire n_3676;
wire n_1054;
wire n_508;
wire n_1679;
wire n_3292;
wire n_3389;
wire n_2872;
wire n_2126;
wire n_3701;
wire n_3109;
wire n_3706;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_3989;
wire n_1858;
wire n_3125;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_3537;
wire n_1057;
wire n_4131;
wire n_2487;
wire n_1834;
wire n_4215;
wire n_1011;
wire n_978;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_2941;
wire n_4158;
wire n_1411;
wire n_1359;
wire n_4286;
wire n_3079;
wire n_3638;
wire n_3269;
wire n_558;
wire n_3536;
wire n_1721;
wire n_2564;
wire n_3558;
wire n_3576;
wire n_3782;
wire n_4231;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_3034;
wire n_2050;
wire n_2197;
wire n_3502;
wire n_3248;
wire n_783;
wire n_4053;
wire n_2550;
wire n_1127;
wire n_556;
wire n_1536;
wire n_3177;
wire n_3594;
wire n_1471;
wire n_2385;
wire n_3440;
wire n_2387;
wire n_1008;
wire n_3963;
wire n_4318;
wire n_3658;
wire n_581;
wire n_3091;
wire n_1024;
wire n_830;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_4177;
wire n_2501;
wire n_2542;
wire n_3227;
wire n_3570;
wire n_3105;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_541;
wire n_499;
wire n_2604;
wire n_1775;
wire n_788;
wire n_908;
wire n_2639;
wire n_3521;
wire n_3855;
wire n_1036;
wire n_2169;
wire n_2985;
wire n_2603;
wire n_4083;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_2630;
wire n_591;
wire n_4105;
wire n_2794;
wire n_969;
wire n_3663;
wire n_2028;
wire n_919;
wire n_1663;
wire n_3114;
wire n_2901;
wire n_2092;
wire n_3940;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_3225;
wire n_3622;
wire n_2817;
wire n_2773;
wire n_1926;
wire n_2402;
wire n_3621;
wire n_1458;
wire n_679;
wire n_1630;
wire n_3473;
wire n_3644;
wire n_3047;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3163;
wire n_3680;
wire n_443;
wire n_3431;
wire n_2176;
wire n_3565;
wire n_1412;
wire n_3355;
wire n_3059;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_826;
wire n_3897;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_3331;
wire n_1735;
wire n_1788;
wire n_940;
wire n_3520;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_4005;
wire n_3272;
wire n_3122;
wire n_3040;
wire n_4230;
wire n_4181;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_607;
wire n_956;
wire n_445;
wire n_3360;
wire n_4187;
wire n_1930;
wire n_3687;
wire n_765;
wire n_1809;
wire n_2787;
wire n_4092;
wire n_3585;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_4037;
wire n_1268;
wire n_3804;
wire n_2676;
wire n_4255;
wire n_2758;
wire n_3211;
wire n_2395;
wire n_917;
wire n_2868;
wire n_1271;
wire n_2096;
wire n_2556;
wire n_2440;
wire n_2186;
wire n_2215;
wire n_1530;
wire n_4057;
wire n_2770;
wire n_631;
wire n_3847;
wire n_1170;
wire n_2724;
wire n_4073;
wire n_3575;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_3633;
wire n_857;
wire n_898;
wire n_3042;
wire n_968;
wire n_1067;
wire n_4144;
wire n_1323;
wire n_1235;
wire n_2584;
wire n_2375;
wire n_3278;
wire n_1462;
wire n_3328;
wire n_4001;
wire n_1937;
wire n_2012;
wire n_3182;
wire n_4167;
wire n_2967;
wire n_3608;
wire n_1064;
wire n_633;
wire n_900;
wire n_4142;
wire n_1446;
wire n_1282;
wire n_3004;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_4021;
wire n_1285;
wire n_3379;
wire n_3111;
wire n_761;
wire n_733;
wire n_2212;
wire n_3838;
wire n_731;
wire n_1813;
wire n_2268;
wire n_2997;
wire n_3469;
wire n_4059;
wire n_2835;
wire n_1452;
wire n_1573;
wire n_3258;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_4019;
wire n_4199;
wire n_3691;
wire n_2252;
wire n_3598;
wire n_2111;
wire n_3743;
wire n_2420;
wire n_2948;
wire n_3099;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_816;
wire n_2897;
wire n_1322;
wire n_3273;
wire n_3829;
wire n_2583;
wire n_2918;
wire n_2987;
wire n_1473;
wire n_835;
wire n_3155;
wire n_4300;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_1003;
wire n_701;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_2358;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_3632;
wire n_2463;
wire n_3546;
wire n_1344;
wire n_2580;
wire n_2355;
wire n_1390;
wire n_2699;
wire n_485;
wire n_1792;
wire n_4064;
wire n_504;
wire n_3351;
wire n_2062;
wire n_483;
wire n_435;
wire n_3068;
wire n_1141;
wire n_3457;
wire n_1629;
wire n_3901;
wire n_1640;
wire n_822;
wire n_1094;
wire n_2973;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_3454;
wire n_3002;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_3146;
wire n_3394;
wire n_3038;
wire n_759;
wire n_567;
wire n_4156;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_3693;
wire n_3878;
wire n_4197;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_3132;
wire n_2615;
wire n_614;
wire n_3776;
wire n_4066;
wire n_2775;
wire n_3903;
wire n_1212;
wire n_3581;
wire n_3778;
wire n_831;
wire n_3681;
wire n_4310;
wire n_3933;
wire n_3970;
wire n_778;
wire n_1619;
wire n_2351;
wire n_4322;
wire n_3303;
wire n_2260;
wire n_550;
wire n_1315;
wire n_1660;
wire n_4080;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2784;
wire n_3898;
wire n_2541;
wire n_694;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_3232;
wire n_3001;
wire n_3188;
wire n_1113;
wire n_3218;
wire n_2347;
wire n_3768;
wire n_1152;
wire n_2657;
wire n_2990;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_4295;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2101;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_4193;
wire n_4100;
wire n_2104;
wire n_1265;
wire n_2552;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1806;
wire n_1533;
wire n_2372;
wire n_1576;
wire n_3445;
wire n_4087;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2933;
wire n_3729;
wire n_3253;
wire n_2856;
wire n_3235;
wire n_3387;
wire n_2088;
wire n_3265;
wire n_3952;
wire n_1275;
wire n_3103;
wire n_488;
wire n_3018;
wire n_4238;
wire n_904;
wire n_505;
wire n_2005;
wire n_3584;
wire n_2048;
wire n_1696;
wire n_3446;
wire n_498;
wire n_3028;
wire n_1875;
wire n_1059;
wire n_3148;
wire n_3775;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_3966;
wire n_3285;
wire n_3824;
wire n_3825;
wire n_4198;
wire n_1039;
wire n_2246;
wire n_3616;
wire n_539;
wire n_1150;
wire n_4266;
wire n_977;
wire n_449;
wire n_2339;
wire n_3846;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_2971;
wire n_3874;
wire n_1497;
wire n_4189;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_4165;
wire n_4154;
wire n_2056;
wire n_2852;
wire n_459;
wire n_1136;
wire n_2515;
wire n_3845;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_3203;
wire n_838;
wire n_1558;
wire n_4107;
wire n_1941;
wire n_3628;
wire n_1316;
wire n_2519;
wire n_3637;
wire n_950;
wire n_1017;
wire n_711;
wire n_3941;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_4168;
wire n_1369;
wire n_4258;
wire n_2846;
wire n_4298;
wire n_3371;
wire n_1781;
wire n_709;
wire n_2917;
wire n_3137;
wire n_4250;
wire n_2544;
wire n_809;
wire n_3143;
wire n_3194;
wire n_3690;
wire n_2085;
wire n_2432;
wire n_3229;
wire n_3032;
wire n_3872;
wire n_1686;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_4232;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_2097;
wire n_1982;
wire n_662;
wire n_641;
wire n_3366;
wire n_3461;
wire n_2430;
wire n_2504;
wire n_910;
wire n_4211;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_3094;
wire n_4276;
wire n_3441;
wire n_4203;
wire n_3020;
wire n_4146;
wire n_4002;
wire n_2964;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_3815;
wire n_2545;
wire n_2513;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_2957;
wire n_865;
wire n_1273;
wire n_1983;
wire n_2982;
wire n_1041;
wire n_2451;
wire n_3312;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_3752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_1810;
wire n_3061;
wire n_448;
wire n_2587;
wire n_3504;
wire n_1347;
wire n_2839;
wire n_3237;
wire n_860;
wire n_3555;
wire n_3820;
wire n_3072;
wire n_4128;
wire n_1043;
wire n_2961;
wire n_2869;
wire n_3534;
wire n_450;
wire n_4036;
wire n_1923;
wire n_3848;
wire n_3655;
wire n_2955;
wire n_2670;
wire n_3631;
wire n_1764;
wire n_2674;
wire n_3556;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_3026;
wire n_2644;
wire n_902;
wire n_1031;
wire n_2979;
wire n_1723;
wire n_3674;
wire n_1638;
wire n_853;
wire n_3071;
wire n_4010;
wire n_716;
wire n_3918;
wire n_4329;
wire n_1571;
wire n_1698;
wire n_3902;
wire n_4101;
wire n_3866;
wire n_1337;
wire n_3763;
wire n_774;
wire n_2148;
wire n_1946;
wire n_933;
wire n_3244;
wire n_3499;
wire n_1779;
wire n_2562;
wire n_596;
wire n_954;
wire n_2051;
wire n_3112;
wire n_1168;
wire n_1821;
wire n_4095;
wire n_1310;
wire n_3296;
wire n_3196;
wire n_3794;
wire n_3910;
wire n_3947;
wire n_3762;
wire n_656;
wire n_492;
wire n_574;
wire n_4205;
wire n_3593;
wire n_2673;
wire n_664;
wire n_1591;
wire n_2585;
wire n_2995;
wire n_3361;
wire n_3293;
wire n_4287;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_3228;
wire n_3327;
wire n_2548;
wire n_3488;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_3707;
wire n_1091;
wire n_2485;
wire n_2052;
wire n_3779;
wire n_3895;
wire n_3149;
wire n_537;
wire n_1063;
wire n_3934;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_3088;
wire n_4224;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_3590;
wire n_2058;
wire n_3231;
wire n_1126;
wire n_3834;
wire n_2761;
wire n_2357;
wire n_4303;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_3923;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_4161;
wire n_2875;
wire n_1639;
wire n_583;
wire n_3519;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_1000;
wire n_626;
wire n_4042;
wire n_1581;
wire n_3849;
wire n_4244;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_3058;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_3398;
wire n_3709;
wire n_1634;
wire n_4265;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_3557;
wire n_3592;
wire n_3725;
wire n_3986;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_4026;
wire n_4245;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_3399;
wire n_3894;
wire n_3202;
wire n_1794;
wire n_4290;
wire n_1375;
wire n_3053;
wire n_1232;
wire n_1211;
wire n_1368;
wire n_996;
wire n_963;
wire n_3772;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_3128;
wire n_4149;
wire n_4120;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2819;
wire n_1115;
wire n_2229;
wire n_2361;
wire n_2880;
wire n_3030;
wire n_3075;
wire n_3505;
wire n_4277;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_3547;
wire n_4014;
wire n_3771;
wire n_2551;
wire n_1102;
wire n_719;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_3045;
wire n_1464;
wire n_1296;
wire n_3158;
wire n_773;
wire n_2798;
wire n_3221;
wire n_2316;
wire n_3217;
wire n_2464;
wire n_3697;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_4222;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_3821;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_3201;
wire n_3334;
wire n_4016;
wire n_2573;
wire n_2940;
wire n_3503;
wire n_548;
wire n_3427;
wire n_2336;
wire n_523;
wire n_1662;
wire n_3162;
wire n_457;
wire n_1299;
wire n_1870;
wire n_3249;
wire n_3483;
wire n_3430;
wire n_4046;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2915;
wire n_3489;
wire n_3083;
wire n_431;
wire n_2654;
wire n_3935;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_3213;
wire n_2517;
wire n_1931;
wire n_4047;
wire n_1244;
wire n_3484;
wire n_1796;
wire n_484;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2965;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_3041;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_2689;
wire n_2423;
wire n_4063;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_3798;
wire n_3080;
wire n_1808;
wire n_1574;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_3033;
wire n_1704;
wire n_3832;
wire n_893;
wire n_3525;
wire n_3308;
wire n_3712;
wire n_1582;
wire n_841;
wire n_2479;
wire n_3204;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_4134;
wire n_2037;
wire n_4305;
wire n_2953;
wire n_3428;
wire n_1308;
wire n_573;
wire n_796;
wire n_2851;
wire n_2823;
wire n_4017;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_146),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_376),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_264),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_338),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_5),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_278),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_395),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_190),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_423),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_308),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g439 ( 
.A(n_384),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_191),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_64),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_337),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_189),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_154),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_107),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_204),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_249),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_394),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_121),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_327),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_303),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_413),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_210),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_17),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_276),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_162),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_26),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g458 ( 
.A(n_267),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_240),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_225),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_291),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_367),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_202),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_304),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_305),
.Y(n_465)
);

BUFx10_ASAP7_75t_L g466 ( 
.A(n_352),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_419),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_343),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_240),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_196),
.Y(n_470)
);

BUFx10_ASAP7_75t_L g471 ( 
.A(n_380),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_3),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_239),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_288),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_195),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_140),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_185),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_125),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_244),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_58),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_351),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_102),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_391),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_165),
.Y(n_484)
);

BUFx10_ASAP7_75t_L g485 ( 
.A(n_271),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_322),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_314),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_397),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_183),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_173),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_16),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_424),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_262),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_289),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_7),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_74),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_398),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_252),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_387),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_283),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_345),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_385),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_130),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_7),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_46),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_127),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_307),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_52),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_18),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_269),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_313),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_116),
.Y(n_512)
);

BUFx10_ASAP7_75t_L g513 ( 
.A(n_184),
.Y(n_513)
);

CKINVDCx14_ASAP7_75t_R g514 ( 
.A(n_127),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_426),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_188),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_120),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_360),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_273),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_173),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_62),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_184),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_411),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_174),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_96),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_321),
.Y(n_526)
);

BUFx10_ASAP7_75t_L g527 ( 
.A(n_97),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_223),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_73),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_146),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_123),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g532 ( 
.A(n_63),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_138),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_57),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_25),
.Y(n_535)
);

BUFx2_ASAP7_75t_SL g536 ( 
.A(n_382),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_231),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_378),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_350),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_275),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_98),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_324),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_417),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_368),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_86),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_56),
.Y(n_546)
);

CKINVDCx14_ASAP7_75t_R g547 ( 
.A(n_138),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_414),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_191),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_249),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_330),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_244),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_185),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_0),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_318),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_356),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_342),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_104),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_422),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_346),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_111),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_386),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_399),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_246),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_235),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_50),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_210),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_377),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_250),
.Y(n_569)
);

CKINVDCx16_ASAP7_75t_R g570 ( 
.A(n_103),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_281),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_409),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_139),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_189),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_255),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_165),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_160),
.Y(n_577)
);

INVxp67_ASAP7_75t_SL g578 ( 
.A(n_155),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_55),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_301),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_299),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_239),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_268),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_207),
.Y(n_584)
);

BUFx10_ASAP7_75t_L g585 ( 
.A(n_392),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_79),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_290),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_260),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_73),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_364),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_175),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_154),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_4),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_79),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_336),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_179),
.Y(n_596)
);

CKINVDCx16_ASAP7_75t_R g597 ( 
.A(n_254),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_347),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_18),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_408),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_65),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_113),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_311),
.Y(n_603)
);

CKINVDCx20_ASAP7_75t_R g604 ( 
.A(n_29),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_1),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_41),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_167),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_300),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_205),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_58),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_77),
.Y(n_611)
);

INVx1_ASAP7_75t_SL g612 ( 
.A(n_354),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_121),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_362),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_293),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_88),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_247),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_22),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_5),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_63),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_339),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_204),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_251),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_161),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_14),
.Y(n_625)
);

CKINVDCx16_ASAP7_75t_R g626 ( 
.A(n_178),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_209),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_361),
.Y(n_628)
);

INVxp67_ASAP7_75t_L g629 ( 
.A(n_270),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_265),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_20),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_323),
.Y(n_632)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_222),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_48),
.Y(n_634)
);

CKINVDCx14_ASAP7_75t_R g635 ( 
.A(n_10),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_15),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_250),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_237),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_55),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_105),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_405),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_258),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_61),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_226),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_144),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_61),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_344),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_134),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_253),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_375),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_25),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_160),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_196),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_363),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_141),
.Y(n_655)
);

CKINVDCx20_ASAP7_75t_R g656 ( 
.A(n_353),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_400),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_8),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_34),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_274),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_252),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_277),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_83),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_98),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_136),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_225),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_286),
.Y(n_667)
);

INVx1_ASAP7_75t_SL g668 ( 
.A(n_373),
.Y(n_668)
);

BUFx5_ASAP7_75t_L g669 ( 
.A(n_33),
.Y(n_669)
);

BUFx10_ASAP7_75t_L g670 ( 
.A(n_282),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_341),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_64),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_228),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_381),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_334),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_125),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_113),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_141),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_393),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_272),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_103),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_206),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_229),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_96),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_372),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_161),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_403),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_1),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_416),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_67),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_359),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_107),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_215),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_157),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_179),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_233),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_105),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_213),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_29),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_130),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_315),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_247),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_211),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_374),
.Y(n_704)
);

CKINVDCx20_ASAP7_75t_R g705 ( 
.A(n_379),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_331),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_144),
.Y(n_707)
);

BUFx10_ASAP7_75t_L g708 ( 
.A(n_41),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_237),
.Y(n_709)
);

INVxp67_ASAP7_75t_SL g710 ( 
.A(n_383),
.Y(n_710)
);

CKINVDCx16_ASAP7_75t_R g711 ( 
.A(n_84),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_335),
.Y(n_712)
);

CKINVDCx14_ASAP7_75t_R g713 ( 
.A(n_366),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_152),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_255),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_370),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_122),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_200),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_59),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_310),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_91),
.Y(n_721)
);

CKINVDCx14_ASAP7_75t_R g722 ( 
.A(n_94),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_412),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_231),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_246),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_116),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_197),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_188),
.Y(n_728)
);

CKINVDCx14_ASAP7_75t_R g729 ( 
.A(n_74),
.Y(n_729)
);

INVx1_ASAP7_75t_SL g730 ( 
.A(n_238),
.Y(n_730)
);

CKINVDCx14_ASAP7_75t_R g731 ( 
.A(n_248),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_223),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_129),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_159),
.Y(n_734)
);

HB1xp67_ASAP7_75t_L g735 ( 
.A(n_371),
.Y(n_735)
);

BUFx8_ASAP7_75t_SL g736 ( 
.A(n_358),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_77),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_178),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_143),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_139),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_56),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_84),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_404),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_227),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_108),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_396),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_150),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_62),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_213),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_230),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_202),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_348),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_355),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_415),
.Y(n_754)
);

CKINVDCx16_ASAP7_75t_R g755 ( 
.A(n_16),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_253),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_245),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_721),
.Y(n_758)
);

CKINVDCx16_ASAP7_75t_R g759 ( 
.A(n_514),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_669),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_669),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_547),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_621),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_669),
.Y(n_764)
);

BUFx2_ASAP7_75t_L g765 ( 
.A(n_635),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_722),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_669),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_669),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_669),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_669),
.Y(n_770)
);

HB1xp67_ASAP7_75t_L g771 ( 
.A(n_532),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_669),
.Y(n_772)
);

INVxp33_ASAP7_75t_SL g773 ( 
.A(n_445),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_721),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_721),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_729),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_453),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_453),
.Y(n_778)
);

NOR2xp67_ASAP7_75t_L g779 ( 
.A(n_460),
.B(n_0),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_731),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_443),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_443),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_444),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_581),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_669),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_466),
.Y(n_786)
);

INVx1_ASAP7_75t_SL g787 ( 
.A(n_429),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_466),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_466),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_622),
.Y(n_790)
);

BUFx10_ASAP7_75t_L g791 ( 
.A(n_735),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_446),
.Y(n_792)
);

CKINVDCx16_ASAP7_75t_R g793 ( 
.A(n_532),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_434),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_466),
.Y(n_795)
);

INVxp67_ASAP7_75t_SL g796 ( 
.A(n_622),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_471),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_471),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_471),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_446),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_434),
.Y(n_801)
);

BUFx10_ASAP7_75t_L g802 ( 
.A(n_622),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_471),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_570),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_622),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_456),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_456),
.Y(n_807)
);

CKINVDCx16_ASAP7_75t_R g808 ( 
.A(n_570),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_457),
.Y(n_809)
);

CKINVDCx20_ASAP7_75t_R g810 ( 
.A(n_600),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_457),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_622),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_434),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_470),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_470),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_485),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_472),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_472),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_482),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_482),
.Y(n_820)
);

CKINVDCx14_ASAP7_75t_R g821 ( 
.A(n_713),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_622),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_485),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_603),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_485),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_505),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_485),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_656),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_585),
.Y(n_829)
);

CKINVDCx16_ASAP7_75t_R g830 ( 
.A(n_597),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_585),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_432),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_432),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_435),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_435),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_442),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_585),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_442),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_585),
.Y(n_839)
);

OR2x2_ASAP7_75t_L g840 ( 
.A(n_597),
.B(n_2),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_670),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_670),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_670),
.Y(n_843)
);

BUFx2_ASAP7_75t_L g844 ( 
.A(n_626),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_448),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_621),
.Y(n_846)
);

BUFx2_ASAP7_75t_L g847 ( 
.A(n_626),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_448),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_455),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_455),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_513),
.Y(n_851)
);

CKINVDCx20_ASAP7_75t_R g852 ( 
.A(n_705),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_621),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_670),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_464),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_711),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_711),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_465),
.Y(n_858)
);

NOR2xp67_ASAP7_75t_L g859 ( 
.A(n_460),
.B(n_2),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_465),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_755),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_755),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_736),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_464),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_474),
.Y(n_865)
);

INVxp67_ASAP7_75t_L g866 ( 
.A(n_505),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_720),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_474),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_509),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_433),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_488),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_488),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_493),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_625),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_440),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_441),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_493),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_434),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_497),
.B(n_3),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_497),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_500),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_447),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_500),
.Y(n_883)
);

CKINVDCx14_ASAP7_75t_R g884 ( 
.A(n_513),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_449),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_501),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_501),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_523),
.B(n_4),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_523),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_509),
.Y(n_890)
);

CKINVDCx16_ASAP7_75t_R g891 ( 
.A(n_513),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_512),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_512),
.Y(n_893)
);

CKINVDCx20_ASAP7_75t_R g894 ( 
.A(n_604),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_517),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_454),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_625),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_517),
.Y(n_898)
);

INVxp33_ASAP7_75t_L g899 ( 
.A(n_522),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_522),
.Y(n_900)
);

CKINVDCx20_ASAP7_75t_R g901 ( 
.A(n_633),
.Y(n_901)
);

CKINVDCx20_ASAP7_75t_R g902 ( 
.A(n_646),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_463),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_528),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_528),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_473),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_529),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_529),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_475),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_535),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_476),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_535),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_537),
.Y(n_913)
);

CKINVDCx20_ASAP7_75t_R g914 ( 
.A(n_707),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_477),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_537),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_625),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_545),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_545),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_552),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_552),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_478),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_554),
.Y(n_923)
);

BUFx2_ASAP7_75t_L g924 ( 
.A(n_533),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_479),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_554),
.Y(n_926)
);

INVxp33_ASAP7_75t_L g927 ( 
.A(n_558),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_484),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_558),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_573),
.Y(n_930)
);

INVx1_ASAP7_75t_SL g931 ( 
.A(n_436),
.Y(n_931)
);

CKINVDCx20_ASAP7_75t_R g932 ( 
.A(n_487),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_573),
.Y(n_933)
);

CKINVDCx20_ASAP7_75t_R g934 ( 
.A(n_487),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_489),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_625),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_490),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_575),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_575),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_491),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_434),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_576),
.Y(n_942)
);

INVxp67_ASAP7_75t_SL g943 ( 
.A(n_625),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_499),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_495),
.Y(n_945)
);

INVxp67_ASAP7_75t_SL g946 ( 
.A(n_625),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_576),
.Y(n_947)
);

CKINVDCx20_ASAP7_75t_R g948 ( 
.A(n_499),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_526),
.B(n_6),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_599),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_496),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_599),
.Y(n_952)
);

BUFx3_ASAP7_75t_L g953 ( 
.A(n_687),
.Y(n_953)
);

INVxp67_ASAP7_75t_L g954 ( 
.A(n_602),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_602),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_605),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_498),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_605),
.Y(n_958)
);

CKINVDCx14_ASAP7_75t_R g959 ( 
.A(n_513),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_609),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_609),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_610),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_503),
.Y(n_963)
);

INVxp67_ASAP7_75t_SL g964 ( 
.A(n_610),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_618),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_618),
.Y(n_966)
);

CKINVDCx20_ASAP7_75t_R g967 ( 
.A(n_687),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_723),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_624),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_624),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_627),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_723),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_627),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_634),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_634),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_636),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_636),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_640),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_640),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_504),
.Y(n_980)
);

CKINVDCx14_ASAP7_75t_R g981 ( 
.A(n_527),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_643),
.Y(n_982)
);

HB1xp67_ASAP7_75t_L g983 ( 
.A(n_506),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_526),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_544),
.Y(n_985)
);

NOR2xp67_ASAP7_75t_L g986 ( 
.A(n_533),
.B(n_6),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_643),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_544),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_652),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_508),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_548),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_652),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_658),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_658),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_666),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_666),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_548),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_516),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_557),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_520),
.Y(n_1000)
);

NOR2xp67_ASAP7_75t_L g1001 ( 
.A(n_534),
.B(n_663),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_521),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_673),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_524),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_673),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_557),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_525),
.Y(n_1007)
);

CKINVDCx20_ASAP7_75t_R g1008 ( 
.A(n_527),
.Y(n_1008)
);

INVxp67_ASAP7_75t_SL g1009 ( 
.A(n_676),
.Y(n_1009)
);

CKINVDCx20_ASAP7_75t_R g1010 ( 
.A(n_527),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_530),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_531),
.Y(n_1012)
);

CKINVDCx16_ASAP7_75t_R g1013 ( 
.A(n_527),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_676),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_459),
.Y(n_1015)
);

INVx1_ASAP7_75t_SL g1016 ( 
.A(n_469),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_541),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_546),
.Y(n_1018)
);

BUFx3_ASAP7_75t_L g1019 ( 
.A(n_562),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_562),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_549),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_682),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_682),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_563),
.Y(n_1024)
);

INVx2_ASAP7_75t_SL g1025 ( 
.A(n_708),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_686),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_434),
.Y(n_1027)
);

CKINVDCx20_ASAP7_75t_R g1028 ( 
.A(n_708),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_686),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_690),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_550),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_690),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_563),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_697),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_583),
.B(n_588),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_583),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_553),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_697),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_715),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_715),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_725),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_588),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_561),
.Y(n_1043)
);

BUFx3_ASAP7_75t_L g1044 ( 
.A(n_614),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_564),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_725),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_732),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_732),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_699),
.Y(n_1049)
);

CKINVDCx14_ASAP7_75t_R g1050 ( 
.A(n_708),
.Y(n_1050)
);

INVxp67_ASAP7_75t_L g1051 ( 
.A(n_739),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_739),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_565),
.Y(n_1053)
);

NOR2xp67_ASAP7_75t_L g1054 ( 
.A(n_534),
.B(n_8),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_741),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_741),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_742),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_742),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_614),
.Y(n_1059)
);

NOR2xp67_ASAP7_75t_L g1060 ( 
.A(n_663),
.B(n_9),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_744),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_630),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_630),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_566),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_744),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_650),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_569),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_574),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_749),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_507),
.Y(n_1070)
);

HB1xp67_ASAP7_75t_L g1071 ( 
.A(n_577),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_749),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_579),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_750),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_750),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_751),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_751),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_582),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_584),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_586),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_589),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_756),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_650),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_756),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_480),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_480),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_657),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_591),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_657),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_679),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_679),
.B(n_9),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_754),
.Y(n_1092)
);

INVxp33_ASAP7_75t_SL g1093 ( 
.A(n_592),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_593),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_594),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_507),
.Y(n_1096)
);

INVxp67_ASAP7_75t_SL g1097 ( 
.A(n_567),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_596),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_507),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_754),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_518),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_601),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_606),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_607),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_567),
.Y(n_1105)
);

CKINVDCx20_ASAP7_75t_R g1106 ( 
.A(n_708),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_692),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_692),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_611),
.Y(n_1109)
);

INVx1_ASAP7_75t_SL g1110 ( 
.A(n_730),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_693),
.Y(n_1111)
);

CKINVDCx16_ASAP7_75t_R g1112 ( 
.A(n_536),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_693),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_613),
.Y(n_1114)
);

CKINVDCx20_ASAP7_75t_R g1115 ( 
.A(n_616),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_617),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_619),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_726),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_894),
.Y(n_1119)
);

CKINVDCx20_ASAP7_75t_R g1120 ( 
.A(n_901),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1112),
.B(n_511),
.Y(n_1121)
);

INVxp67_ASAP7_75t_L g1122 ( 
.A(n_931),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_867),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_790),
.Y(n_1124)
);

CKINVDCx20_ASAP7_75t_R g1125 ( 
.A(n_902),
.Y(n_1125)
);

INVxp33_ASAP7_75t_L g1126 ( 
.A(n_771),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_867),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_758),
.Y(n_1128)
);

CKINVDCx20_ASAP7_75t_R g1129 ( 
.A(n_914),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_774),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_775),
.Y(n_1131)
);

INVxp67_ASAP7_75t_SL g1132 ( 
.A(n_763),
.Y(n_1132)
);

CKINVDCx20_ASAP7_75t_R g1133 ( 
.A(n_784),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_790),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_821),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_810),
.Y(n_1136)
);

CKINVDCx20_ASAP7_75t_R g1137 ( 
.A(n_824),
.Y(n_1137)
);

HB1xp67_ASAP7_75t_L g1138 ( 
.A(n_1015),
.Y(n_1138)
);

CKINVDCx20_ASAP7_75t_R g1139 ( 
.A(n_828),
.Y(n_1139)
);

CKINVDCx20_ASAP7_75t_R g1140 ( 
.A(n_852),
.Y(n_1140)
);

INVxp67_ASAP7_75t_L g1141 ( 
.A(n_1016),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_884),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_786),
.B(n_629),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_796),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_943),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_946),
.Y(n_1146)
);

INVxp67_ASAP7_75t_L g1147 ( 
.A(n_1049),
.Y(n_1147)
);

HB1xp67_ASAP7_75t_L g1148 ( 
.A(n_1110),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_832),
.Y(n_1149)
);

CKINVDCx20_ASAP7_75t_R g1150 ( 
.A(n_1115),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_832),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_833),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_763),
.B(n_511),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_786),
.B(n_439),
.Y(n_1154)
);

CKINVDCx16_ASAP7_75t_R g1155 ( 
.A(n_759),
.Y(n_1155)
);

NOR2xp67_ASAP7_75t_L g1156 ( 
.A(n_863),
.B(n_430),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_833),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_805),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_959),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_844),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_981),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_834),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_1050),
.Y(n_1163)
);

CKINVDCx20_ASAP7_75t_R g1164 ( 
.A(n_932),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_834),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_835),
.Y(n_1166)
);

HB1xp67_ASAP7_75t_L g1167 ( 
.A(n_793),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_863),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_934),
.Y(n_1169)
);

CKINVDCx20_ASAP7_75t_R g1170 ( 
.A(n_944),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_788),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_835),
.Y(n_1172)
);

CKINVDCx20_ASAP7_75t_R g1173 ( 
.A(n_948),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_836),
.Y(n_1174)
);

CKINVDCx20_ASAP7_75t_R g1175 ( 
.A(n_967),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_808),
.Y(n_1176)
);

BUFx10_ASAP7_75t_L g1177 ( 
.A(n_788),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_789),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_844),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_789),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_760),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_795),
.B(n_797),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_795),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_760),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_797),
.Y(n_1185)
);

CKINVDCx16_ASAP7_75t_R g1186 ( 
.A(n_891),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_798),
.Y(n_1187)
);

CKINVDCx20_ASAP7_75t_R g1188 ( 
.A(n_787),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_798),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_761),
.Y(n_1190)
);

CKINVDCx20_ASAP7_75t_R g1191 ( 
.A(n_1008),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_799),
.Y(n_1192)
);

BUFx6f_ASAP7_75t_L g1193 ( 
.A(n_794),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_761),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_836),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_838),
.Y(n_1196)
);

CKINVDCx16_ASAP7_75t_R g1197 ( 
.A(n_1013),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_799),
.Y(n_1198)
);

INVxp67_ASAP7_75t_SL g1199 ( 
.A(n_846),
.Y(n_1199)
);

CKINVDCx16_ASAP7_75t_R g1200 ( 
.A(n_830),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_838),
.Y(n_1201)
);

INVxp67_ASAP7_75t_SL g1202 ( 
.A(n_846),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_803),
.B(n_458),
.Y(n_1203)
);

INVxp67_ASAP7_75t_SL g1204 ( 
.A(n_853),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_803),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_847),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_856),
.Y(n_1207)
);

BUFx2_ASAP7_75t_L g1208 ( 
.A(n_847),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_845),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_816),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_853),
.B(n_518),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_816),
.B(n_612),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_823),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_845),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_848),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_848),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_849),
.Y(n_1217)
);

INVxp67_ASAP7_75t_SL g1218 ( 
.A(n_858),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_1010),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_823),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_849),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_850),
.Y(n_1222)
);

INVxp67_ASAP7_75t_L g1223 ( 
.A(n_983),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_805),
.Y(n_1224)
);

NOR2xp67_ASAP7_75t_L g1225 ( 
.A(n_825),
.B(n_431),
.Y(n_1225)
);

CKINVDCx20_ASAP7_75t_R g1226 ( 
.A(n_1028),
.Y(n_1226)
);

INVxp67_ASAP7_75t_SL g1227 ( 
.A(n_858),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_850),
.Y(n_1228)
);

CKINVDCx20_ASAP7_75t_R g1229 ( 
.A(n_1106),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_855),
.Y(n_1230)
);

CKINVDCx20_ASAP7_75t_R g1231 ( 
.A(n_825),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_812),
.Y(n_1232)
);

CKINVDCx20_ASAP7_75t_R g1233 ( 
.A(n_827),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_855),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_864),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_864),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_827),
.B(n_829),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_865),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_865),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_829),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_868),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_868),
.Y(n_1242)
);

CKINVDCx20_ASAP7_75t_R g1243 ( 
.A(n_831),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_831),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_871),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_837),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_871),
.Y(n_1247)
);

CKINVDCx20_ASAP7_75t_R g1248 ( 
.A(n_837),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_872),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_839),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_872),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_839),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_841),
.Y(n_1253)
);

INVxp67_ASAP7_75t_L g1254 ( 
.A(n_1071),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_841),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_842),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_873),
.Y(n_1257)
);

CKINVDCx20_ASAP7_75t_R g1258 ( 
.A(n_842),
.Y(n_1258)
);

CKINVDCx20_ASAP7_75t_R g1259 ( 
.A(n_843),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_873),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_877),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_877),
.Y(n_1262)
);

CKINVDCx16_ASAP7_75t_R g1263 ( 
.A(n_765),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_880),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_880),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_843),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_854),
.B(n_654),
.Y(n_1267)
);

INVxp67_ASAP7_75t_SL g1268 ( 
.A(n_860),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_881),
.Y(n_1269)
);

INVxp67_ASAP7_75t_L g1270 ( 
.A(n_804),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_854),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_764),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_762),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_881),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_883),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_762),
.Y(n_1276)
);

INVx3_ASAP7_75t_L g1277 ( 
.A(n_802),
.Y(n_1277)
);

CKINVDCx20_ASAP7_75t_R g1278 ( 
.A(n_856),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_883),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_857),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_766),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_766),
.Y(n_1282)
);

CKINVDCx16_ASAP7_75t_R g1283 ( 
.A(n_765),
.Y(n_1283)
);

CKINVDCx20_ASAP7_75t_R g1284 ( 
.A(n_857),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_886),
.Y(n_1285)
);

CKINVDCx16_ASAP7_75t_R g1286 ( 
.A(n_791),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_861),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_776),
.Y(n_1288)
);

CKINVDCx20_ASAP7_75t_R g1289 ( 
.A(n_861),
.Y(n_1289)
);

CKINVDCx16_ASAP7_75t_R g1290 ( 
.A(n_791),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_776),
.Y(n_1291)
);

CKINVDCx16_ASAP7_75t_R g1292 ( 
.A(n_791),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_862),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_780),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_886),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_780),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_887),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_870),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_862),
.Y(n_1299)
);

NOR2xp67_ASAP7_75t_L g1300 ( 
.A(n_851),
.B(n_437),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_870),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_860),
.B(n_519),
.Y(n_1302)
);

CKINVDCx20_ASAP7_75t_R g1303 ( 
.A(n_875),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_887),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_953),
.B(n_519),
.Y(n_1305)
);

CKINVDCx20_ASAP7_75t_R g1306 ( 
.A(n_875),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_889),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_889),
.Y(n_1308)
);

CKINVDCx20_ASAP7_75t_R g1309 ( 
.A(n_876),
.Y(n_1309)
);

CKINVDCx16_ASAP7_75t_R g1310 ( 
.A(n_840),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_876),
.Y(n_1311)
);

BUFx10_ASAP7_75t_L g1312 ( 
.A(n_882),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_984),
.Y(n_1313)
);

INVxp33_ASAP7_75t_SL g1314 ( 
.A(n_882),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_885),
.Y(n_1315)
);

CKINVDCx20_ASAP7_75t_R g1316 ( 
.A(n_885),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_896),
.Y(n_1317)
);

NOR2xp67_ASAP7_75t_L g1318 ( 
.A(n_851),
.B(n_438),
.Y(n_1318)
);

BUFx10_ASAP7_75t_L g1319 ( 
.A(n_896),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_903),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_903),
.Y(n_1321)
);

NOR2xp67_ASAP7_75t_L g1322 ( 
.A(n_1025),
.B(n_906),
.Y(n_1322)
);

INVxp67_ASAP7_75t_L g1323 ( 
.A(n_1025),
.Y(n_1323)
);

CKINVDCx20_ASAP7_75t_R g1324 ( 
.A(n_906),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_984),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_909),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_909),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_911),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_911),
.Y(n_1329)
);

INVxp67_ASAP7_75t_SL g1330 ( 
.A(n_953),
.Y(n_1330)
);

INVxp33_ASAP7_75t_SL g1331 ( 
.A(n_915),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1093),
.B(n_668),
.Y(n_1332)
);

CKINVDCx20_ASAP7_75t_R g1333 ( 
.A(n_915),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1089),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1089),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1090),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1090),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1092),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1092),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_922),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_812),
.Y(n_1341)
);

CKINVDCx16_ASAP7_75t_R g1342 ( 
.A(n_840),
.Y(n_1342)
);

INVxp67_ASAP7_75t_SL g1343 ( 
.A(n_968),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_922),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_925),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_925),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_968),
.B(n_571),
.Y(n_1347)
);

CKINVDCx20_ASAP7_75t_R g1348 ( 
.A(n_928),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_781),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_782),
.Y(n_1350)
);

INVxp67_ASAP7_75t_SL g1351 ( 
.A(n_972),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_783),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_802),
.Y(n_1353)
);

INVxp67_ASAP7_75t_SL g1354 ( 
.A(n_972),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_928),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_935),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_935),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_792),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_937),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_800),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_937),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_806),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_807),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_764),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_940),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_767),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_940),
.Y(n_1367)
);

NOR2xp67_ASAP7_75t_L g1368 ( 
.A(n_945),
.B(n_450),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_945),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_809),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_964),
.B(n_571),
.Y(n_1371)
);

CKINVDCx20_ASAP7_75t_R g1372 ( 
.A(n_951),
.Y(n_1372)
);

BUFx2_ASAP7_75t_L g1373 ( 
.A(n_951),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_957),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_811),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_814),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_957),
.Y(n_1377)
);

CKINVDCx20_ASAP7_75t_R g1378 ( 
.A(n_963),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_815),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_817),
.Y(n_1380)
);

INVxp33_ASAP7_75t_SL g1381 ( 
.A(n_963),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_818),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_819),
.Y(n_1383)
);

CKINVDCx20_ASAP7_75t_R g1384 ( 
.A(n_980),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_R g1385 ( 
.A(n_980),
.B(n_451),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_990),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_990),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_998),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_820),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_826),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_890),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_892),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_893),
.Y(n_1393)
);

CKINVDCx16_ASAP7_75t_R g1394 ( 
.A(n_924),
.Y(n_1394)
);

CKINVDCx20_ASAP7_75t_R g1395 ( 
.A(n_998),
.Y(n_1395)
);

INVxp67_ASAP7_75t_L g1396 ( 
.A(n_1000),
.Y(n_1396)
);

INVxp67_ASAP7_75t_SL g1397 ( 
.A(n_1035),
.Y(n_1397)
);

CKINVDCx20_ASAP7_75t_R g1398 ( 
.A(n_1000),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1002),
.B(n_641),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1002),
.B(n_641),
.Y(n_1400)
);

CKINVDCx20_ASAP7_75t_R g1401 ( 
.A(n_1004),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_895),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_1004),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_802),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_1007),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_1007),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1011),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1011),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_1012),
.Y(n_1409)
);

INVxp67_ASAP7_75t_SL g1410 ( 
.A(n_988),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1012),
.Y(n_1411)
);

INVxp33_ASAP7_75t_L g1412 ( 
.A(n_899),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1017),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_898),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_1017),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_900),
.Y(n_1416)
);

NOR2xp67_ASAP7_75t_L g1417 ( 
.A(n_1018),
.B(n_452),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1018),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_904),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_905),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_907),
.Y(n_1421)
);

CKINVDCx20_ASAP7_75t_R g1422 ( 
.A(n_1021),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_1021),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1412),
.B(n_988),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1124),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1181),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1181),
.A2(n_785),
.B(n_768),
.Y(n_1427)
);

BUFx6f_ASAP7_75t_L g1428 ( 
.A(n_1193),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1410),
.B(n_1009),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_L g1430 ( 
.A(n_1193),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_1168),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1124),
.Y(n_1432)
);

AOI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1332),
.A2(n_773),
.B1(n_1037),
.B2(n_1031),
.Y(n_1433)
);

CKINVDCx16_ASAP7_75t_R g1434 ( 
.A(n_1200),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1397),
.A2(n_779),
.B1(n_986),
.B2(n_859),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1134),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1149),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1132),
.B(n_997),
.Y(n_1438)
);

AND2x6_ASAP7_75t_L g1439 ( 
.A(n_1151),
.B(n_743),
.Y(n_1439)
);

AND2x4_ASAP7_75t_L g1440 ( 
.A(n_1218),
.B(n_997),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1152),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1122),
.B(n_1019),
.Y(n_1442)
);

INVx1_ASAP7_75t_SL g1443 ( 
.A(n_1138),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1141),
.B(n_1019),
.Y(n_1444)
);

OAI22x1_ASAP7_75t_R g1445 ( 
.A1(n_1423),
.A2(n_1109),
.B1(n_1116),
.B2(n_1114),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1157),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1162),
.Y(n_1447)
);

AOI22x1_ASAP7_75t_R g1448 ( 
.A1(n_1301),
.A2(n_908),
.B1(n_912),
.B2(n_910),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1165),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1199),
.B(n_1033),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1166),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1193),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1184),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1184),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_1353),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1172),
.Y(n_1456)
);

AOI22x1_ASAP7_75t_SL g1457 ( 
.A1(n_1150),
.A2(n_620),
.B1(n_631),
.B2(n_623),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1174),
.Y(n_1458)
);

BUFx8_ASAP7_75t_L g1459 ( 
.A(n_1373),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1323),
.B(n_1031),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1195),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1147),
.B(n_1033),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1193),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1196),
.B(n_1044),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1182),
.A2(n_1060),
.B1(n_1054),
.B2(n_888),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_L g1466 ( 
.A(n_1193),
.Y(n_1466)
);

INVx3_ASAP7_75t_L g1467 ( 
.A(n_1190),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1202),
.B(n_1044),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1134),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1201),
.B(n_1083),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1204),
.B(n_1154),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1203),
.B(n_1212),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1190),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1194),
.Y(n_1474)
);

OAI22x1_ASAP7_75t_R g1475 ( 
.A1(n_1303),
.A2(n_1116),
.B1(n_1104),
.B2(n_1114),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1194),
.Y(n_1476)
);

INVx3_ASAP7_75t_L g1477 ( 
.A(n_1272),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1158),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1158),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1209),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1224),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1224),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1227),
.B(n_1083),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1214),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1353),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1232),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1272),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1232),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1215),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1267),
.B(n_1101),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1341),
.Y(n_1491)
);

CKINVDCx16_ASAP7_75t_R g1492 ( 
.A(n_1186),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1143),
.B(n_1144),
.Y(n_1493)
);

BUFx6f_ASAP7_75t_L g1494 ( 
.A(n_1364),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1341),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1145),
.B(n_1101),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1364),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1268),
.B(n_866),
.Y(n_1498)
);

AND2x6_ASAP7_75t_L g1499 ( 
.A(n_1216),
.B(n_743),
.Y(n_1499)
);

AOI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1399),
.A2(n_1043),
.B1(n_1045),
.B2(n_1037),
.Y(n_1500)
);

AOI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1400),
.A2(n_1322),
.B1(n_1121),
.B2(n_1237),
.Y(n_1501)
);

INVx3_ASAP7_75t_L g1502 ( 
.A(n_1366),
.Y(n_1502)
);

AOI22xp5_ASAP7_75t_SL g1503 ( 
.A1(n_1306),
.A2(n_1117),
.B1(n_1043),
.B2(n_1053),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1366),
.Y(n_1504)
);

BUFx6f_ASAP7_75t_L g1505 ( 
.A(n_1217),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1221),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1222),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_SL g1508 ( 
.A(n_1385),
.B(n_1045),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1228),
.Y(n_1509)
);

INVx4_ASAP7_75t_L g1510 ( 
.A(n_1277),
.Y(n_1510)
);

INVx6_ASAP7_75t_L g1511 ( 
.A(n_1404),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1277),
.Y(n_1512)
);

AOI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1223),
.A2(n_1064),
.B1(n_1067),
.B2(n_1053),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1230),
.Y(n_1514)
);

INVxp67_ASAP7_75t_L g1515 ( 
.A(n_1148),
.Y(n_1515)
);

INVx3_ASAP7_75t_L g1516 ( 
.A(n_1277),
.Y(n_1516)
);

INVx3_ASAP7_75t_L g1517 ( 
.A(n_1234),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1235),
.Y(n_1518)
);

INVx6_ASAP7_75t_L g1519 ( 
.A(n_1404),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1146),
.B(n_985),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1236),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1330),
.B(n_985),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_SL g1523 ( 
.A1(n_1119),
.A2(n_1064),
.B1(n_1068),
.B2(n_1067),
.Y(n_1523)
);

OAI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1153),
.A2(n_785),
.B(n_768),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1238),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_SL g1526 ( 
.A1(n_1120),
.A2(n_1068),
.B1(n_1078),
.B2(n_1073),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1239),
.Y(n_1527)
);

AOI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1254),
.A2(n_1178),
.B1(n_1180),
.B2(n_1171),
.Y(n_1528)
);

CKINVDCx16_ASAP7_75t_R g1529 ( 
.A(n_1197),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1241),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1242),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_L g1532 ( 
.A1(n_1245),
.A2(n_769),
.B(n_767),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1247),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1249),
.Y(n_1534)
);

OAI22x1_ASAP7_75t_R g1535 ( 
.A1(n_1309),
.A2(n_1078),
.B1(n_1079),
.B2(n_1073),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1343),
.B(n_991),
.Y(n_1536)
);

BUFx6f_ASAP7_75t_L g1537 ( 
.A(n_1251),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1257),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1260),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1261),
.Y(n_1540)
);

BUFx6f_ASAP7_75t_L g1541 ( 
.A(n_1262),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1394),
.Y(n_1542)
);

OAI21x1_ASAP7_75t_L g1543 ( 
.A1(n_1264),
.A2(n_770),
.B(n_769),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1265),
.B(n_927),
.Y(n_1544)
);

AOI22xp5_ASAP7_75t_SL g1545 ( 
.A1(n_1316),
.A2(n_1080),
.B1(n_1081),
.B2(n_1079),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1269),
.Y(n_1546)
);

BUFx6f_ASAP7_75t_L g1547 ( 
.A(n_1274),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1275),
.Y(n_1548)
);

BUFx6f_ASAP7_75t_L g1549 ( 
.A(n_1279),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1285),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1160),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1295),
.Y(n_1552)
);

BUFx8_ASAP7_75t_L g1553 ( 
.A(n_1373),
.Y(n_1553)
);

BUFx6f_ASAP7_75t_L g1554 ( 
.A(n_1297),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1304),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1307),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1351),
.B(n_869),
.Y(n_1557)
);

BUFx6f_ASAP7_75t_L g1558 ( 
.A(n_1308),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1313),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1354),
.B(n_991),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1171),
.A2(n_949),
.B1(n_1091),
.B2(n_879),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1178),
.A2(n_1081),
.B1(n_1088),
.B2(n_1080),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1325),
.B(n_1097),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1334),
.Y(n_1564)
);

AND2x4_ASAP7_75t_L g1565 ( 
.A(n_1371),
.B(n_954),
.Y(n_1565)
);

INVx3_ASAP7_75t_L g1566 ( 
.A(n_1335),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1336),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1337),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1338),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1339),
.Y(n_1570)
);

BUFx6f_ASAP7_75t_L g1571 ( 
.A(n_1128),
.Y(n_1571)
);

CKINVDCx11_ASAP7_75t_R g1572 ( 
.A(n_1317),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1349),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1350),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1352),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1130),
.Y(n_1576)
);

BUFx6f_ASAP7_75t_L g1577 ( 
.A(n_1131),
.Y(n_1577)
);

OA21x2_ASAP7_75t_L g1578 ( 
.A1(n_1211),
.A2(n_772),
.B(n_770),
.Y(n_1578)
);

BUFx3_ASAP7_75t_L g1579 ( 
.A(n_1358),
.Y(n_1579)
);

OAI22xp5_ASAP7_75t_SL g1580 ( 
.A1(n_1125),
.A2(n_1094),
.B1(n_1095),
.B2(n_1088),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1360),
.Y(n_1581)
);

AND2x4_ASAP7_75t_L g1582 ( 
.A(n_1362),
.B(n_1051),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1363),
.B(n_924),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1370),
.Y(n_1584)
);

BUFx8_ASAP7_75t_L g1585 ( 
.A(n_1160),
.Y(n_1585)
);

OAI21x1_ASAP7_75t_L g1586 ( 
.A1(n_1302),
.A2(n_772),
.B(n_999),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1375),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1376),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1379),
.Y(n_1589)
);

BUFx6f_ASAP7_75t_L g1590 ( 
.A(n_1380),
.Y(n_1590)
);

INVxp67_ASAP7_75t_L g1591 ( 
.A(n_1167),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1382),
.B(n_1001),
.Y(n_1592)
);

INVx3_ASAP7_75t_L g1593 ( 
.A(n_1383),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1389),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1390),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1179),
.Y(n_1596)
);

BUFx2_ASAP7_75t_L g1597 ( 
.A(n_1179),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1391),
.Y(n_1598)
);

INVx5_ASAP7_75t_L g1599 ( 
.A(n_1177),
.Y(n_1599)
);

BUFx3_ASAP7_75t_L g1600 ( 
.A(n_1392),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1393),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1402),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1177),
.B(n_1094),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1414),
.Y(n_1604)
);

OAI21x1_ASAP7_75t_L g1605 ( 
.A1(n_1305),
.A2(n_1006),
.B(n_999),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1416),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1300),
.B(n_1006),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1419),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1318),
.B(n_1020),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1420),
.Y(n_1610)
);

INVx2_ASAP7_75t_SL g1611 ( 
.A(n_1177),
.Y(n_1611)
);

INVx5_ASAP7_75t_L g1612 ( 
.A(n_1312),
.Y(n_1612)
);

INVx3_ASAP7_75t_L g1613 ( 
.A(n_1421),
.Y(n_1613)
);

INVx5_ASAP7_75t_L g1614 ( 
.A(n_1312),
.Y(n_1614)
);

AND2x4_ASAP7_75t_L g1615 ( 
.A(n_1347),
.B(n_1113),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1368),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1225),
.B(n_1020),
.Y(n_1617)
);

INVx5_ASAP7_75t_L g1618 ( 
.A(n_1312),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1417),
.Y(n_1619)
);

INVx3_ASAP7_75t_L g1620 ( 
.A(n_1319),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1320),
.Y(n_1621)
);

INVx3_ASAP7_75t_L g1622 ( 
.A(n_1319),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1180),
.B(n_1024),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1206),
.B(n_1113),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1206),
.B(n_1024),
.Y(n_1625)
);

AOI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1183),
.A2(n_1098),
.B1(n_1102),
.B2(n_1095),
.Y(n_1626)
);

INVx3_ASAP7_75t_L g1627 ( 
.A(n_1319),
.Y(n_1627)
);

BUFx6f_ASAP7_75t_L g1628 ( 
.A(n_1298),
.Y(n_1628)
);

OAI22xp5_ASAP7_75t_SL g1629 ( 
.A1(n_1129),
.A2(n_1102),
.B1(n_1103),
.B2(n_1098),
.Y(n_1629)
);

BUFx6f_ASAP7_75t_L g1630 ( 
.A(n_1298),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1355),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1408),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1208),
.Y(n_1633)
);

INVx5_ASAP7_75t_L g1634 ( 
.A(n_1155),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1263),
.Y(n_1635)
);

AOI22xp5_ASAP7_75t_SL g1636 ( 
.A1(n_1321),
.A2(n_1104),
.B1(n_1109),
.B2(n_1103),
.Y(n_1636)
);

INVx3_ASAP7_75t_L g1637 ( 
.A(n_1283),
.Y(n_1637)
);

BUFx6f_ASAP7_75t_L g1638 ( 
.A(n_1311),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1183),
.B(n_1036),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1411),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1185),
.B(n_1036),
.Y(n_1641)
);

INVx3_ASAP7_75t_L g1642 ( 
.A(n_1142),
.Y(n_1642)
);

AND2x2_ASAP7_75t_SL g1643 ( 
.A(n_1286),
.B(n_726),
.Y(n_1643)
);

OAI21x1_ASAP7_75t_L g1644 ( 
.A1(n_1156),
.A2(n_1059),
.B(n_1042),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1418),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1208),
.Y(n_1646)
);

INVx3_ASAP7_75t_L g1647 ( 
.A(n_1142),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1396),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1207),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1270),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1280),
.Y(n_1651)
);

INVxp33_ASAP7_75t_L g1652 ( 
.A(n_1126),
.Y(n_1652)
);

INVx3_ASAP7_75t_L g1653 ( 
.A(n_1159),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1185),
.B(n_1042),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1176),
.B(n_913),
.Y(n_1655)
);

OAI21x1_ASAP7_75t_L g1656 ( 
.A1(n_1293),
.A2(n_1062),
.B(n_1059),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1187),
.B(n_1062),
.Y(n_1657)
);

AND2x4_ASAP7_75t_L g1658 ( 
.A(n_1159),
.B(n_916),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1311),
.Y(n_1659)
);

AOI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1187),
.A2(n_1117),
.B1(n_638),
.B2(n_639),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1189),
.B(n_1063),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1161),
.B(n_1063),
.Y(n_1662)
);

INVx4_ASAP7_75t_L g1663 ( 
.A(n_1161),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1163),
.B(n_918),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1315),
.Y(n_1665)
);

BUFx6f_ASAP7_75t_L g1666 ( 
.A(n_1315),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1326),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1189),
.B(n_1066),
.Y(n_1668)
);

BUFx2_ASAP7_75t_L g1669 ( 
.A(n_1278),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1326),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1163),
.B(n_919),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1328),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1328),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1329),
.Y(n_1674)
);

NAND2xp33_ASAP7_75t_L g1675 ( 
.A(n_1192),
.B(n_507),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1329),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1340),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1192),
.B(n_1198),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_SL g1679 ( 
.A1(n_1310),
.A2(n_642),
.B1(n_644),
.B2(n_637),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1340),
.Y(n_1680)
);

BUFx2_ASAP7_75t_L g1681 ( 
.A(n_1284),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1344),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1198),
.A2(n_648),
.B1(n_649),
.B2(n_645),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_1168),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1344),
.Y(n_1685)
);

BUFx8_ASAP7_75t_L g1686 ( 
.A(n_1314),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1205),
.B(n_1066),
.Y(n_1687)
);

INVx4_ASAP7_75t_L g1688 ( 
.A(n_1135),
.Y(n_1688)
);

BUFx2_ASAP7_75t_L g1689 ( 
.A(n_1287),
.Y(n_1689)
);

INVx6_ASAP7_75t_L g1690 ( 
.A(n_1290),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1345),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1345),
.Y(n_1692)
);

OAI22xp5_ASAP7_75t_SL g1693 ( 
.A1(n_1342),
.A2(n_653),
.B1(n_655),
.B2(n_651),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1205),
.B(n_1087),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1346),
.Y(n_1695)
);

BUFx3_ASAP7_75t_L g1696 ( 
.A(n_1135),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1346),
.B(n_920),
.Y(n_1697)
);

OA21x2_ASAP7_75t_L g1698 ( 
.A1(n_1210),
.A2(n_1100),
.B(n_1087),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_1164),
.Y(n_1699)
);

NAND2xp33_ASAP7_75t_L g1700 ( 
.A(n_1210),
.B(n_1213),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1356),
.Y(n_1701)
);

AOI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1213),
.A2(n_661),
.B1(n_664),
.B2(n_659),
.Y(n_1702)
);

INVx6_ASAP7_75t_L g1703 ( 
.A(n_1292),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1356),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1220),
.B(n_1100),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1357),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1357),
.B(n_921),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1359),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1359),
.Y(n_1709)
);

NOR2x1_ASAP7_75t_L g1710 ( 
.A(n_1231),
.B(n_777),
.Y(n_1710)
);

BUFx6f_ASAP7_75t_L g1711 ( 
.A(n_1361),
.Y(n_1711)
);

AOI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1472),
.A2(n_1240),
.B1(n_1246),
.B2(n_1220),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1426),
.Y(n_1713)
);

OAI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1501),
.A2(n_1415),
.B1(n_1365),
.B2(n_1367),
.Y(n_1714)
);

AOI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1561),
.A2(n_1246),
.B1(n_1250),
.B2(n_1240),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_L g1716 ( 
.A(n_1515),
.B(n_1314),
.Y(n_1716)
);

INVx3_ASAP7_75t_L g1717 ( 
.A(n_1505),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1490),
.B(n_1250),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1424),
.B(n_1253),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1443),
.B(n_1136),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1424),
.B(n_1253),
.Y(n_1721)
);

NOR2xp33_ASAP7_75t_L g1722 ( 
.A(n_1652),
.B(n_1331),
.Y(n_1722)
);

AOI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1694),
.A2(n_1271),
.B1(n_1381),
.B2(n_1331),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1426),
.Y(n_1724)
);

OAI22xp33_ASAP7_75t_SL g1725 ( 
.A1(n_1623),
.A2(n_1381),
.B1(n_1123),
.B2(n_1127),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1453),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1497),
.Y(n_1727)
);

BUFx6f_ASAP7_75t_SL g1728 ( 
.A(n_1696),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1442),
.B(n_1271),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1442),
.B(n_1361),
.Y(n_1730)
);

AOI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1694),
.A2(n_1367),
.B1(n_1374),
.B2(n_1365),
.Y(n_1731)
);

OAI22xp33_ASAP7_75t_SL g1732 ( 
.A1(n_1639),
.A2(n_1123),
.B1(n_1127),
.B2(n_1374),
.Y(n_1732)
);

AOI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1698),
.A2(n_578),
.B1(n_1386),
.B2(n_1377),
.Y(n_1733)
);

OAI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1433),
.A2(n_1386),
.B1(n_1387),
.B2(n_1377),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1453),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1551),
.B(n_1136),
.Y(n_1736)
);

INVx1_ASAP7_75t_SL g1737 ( 
.A(n_1444),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1454),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1444),
.B(n_1387),
.Y(n_1739)
);

OAI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1528),
.A2(n_1405),
.B1(n_1406),
.B2(n_1388),
.Y(n_1740)
);

OAI22xp33_ASAP7_75t_SL g1741 ( 
.A1(n_1641),
.A2(n_1405),
.B1(n_1406),
.B2(n_1388),
.Y(n_1741)
);

OAI22xp33_ASAP7_75t_SL g1742 ( 
.A1(n_1654),
.A2(n_1413),
.B1(n_1415),
.B2(n_1407),
.Y(n_1742)
);

CKINVDCx6p67_ASAP7_75t_R g1743 ( 
.A(n_1634),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1497),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1504),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1493),
.B(n_1471),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1462),
.B(n_1407),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1462),
.B(n_1413),
.Y(n_1748)
);

INVx3_ASAP7_75t_L g1749 ( 
.A(n_1505),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1624),
.B(n_1273),
.Y(n_1750)
);

OR2x6_ASAP7_75t_L g1751 ( 
.A(n_1690),
.B(n_1133),
.Y(n_1751)
);

AOI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1698),
.A2(n_1233),
.B1(n_1244),
.B2(n_1243),
.Y(n_1752)
);

OAI22xp33_ASAP7_75t_SL g1753 ( 
.A1(n_1657),
.A2(n_1276),
.B1(n_1281),
.B2(n_1273),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1429),
.B(n_1276),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1504),
.Y(n_1755)
);

AO22x2_ASAP7_75t_L g1756 ( 
.A1(n_1457),
.A2(n_1170),
.B1(n_1173),
.B2(n_1169),
.Y(n_1756)
);

OAI22xp33_ASAP7_75t_SL g1757 ( 
.A1(n_1661),
.A2(n_1668),
.B1(n_1705),
.B2(n_1687),
.Y(n_1757)
);

AOI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1698),
.A2(n_1248),
.B1(n_1255),
.B2(n_1252),
.Y(n_1758)
);

OR2x6_ASAP7_75t_L g1759 ( 
.A(n_1690),
.B(n_1137),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1624),
.B(n_1281),
.Y(n_1760)
);

OAI22xp33_ASAP7_75t_R g1761 ( 
.A1(n_1682),
.A2(n_757),
.B1(n_926),
.B2(n_923),
.Y(n_1761)
);

OA22x2_ASAP7_75t_L g1762 ( 
.A1(n_1542),
.A2(n_1288),
.B1(n_1291),
.B2(n_1282),
.Y(n_1762)
);

AO22x2_ASAP7_75t_L g1763 ( 
.A1(n_1457),
.A2(n_1175),
.B1(n_1140),
.B2(n_1139),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1625),
.B(n_1282),
.Y(n_1764)
);

OAI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1628),
.A2(n_1291),
.B1(n_1294),
.B2(n_1288),
.Y(n_1765)
);

AO22x2_ASAP7_75t_L g1766 ( 
.A1(n_1435),
.A2(n_1191),
.B1(n_1226),
.B2(n_1219),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1625),
.B(n_1697),
.Y(n_1767)
);

AOI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1697),
.A2(n_1707),
.B1(n_1465),
.B2(n_1429),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1697),
.B(n_1294),
.Y(n_1769)
);

AOI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1707),
.A2(n_1429),
.B1(n_1557),
.B2(n_1498),
.Y(n_1770)
);

AOI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1707),
.A2(n_1258),
.B1(n_1259),
.B2(n_1256),
.Y(n_1771)
);

OR2x6_ASAP7_75t_L g1772 ( 
.A(n_1690),
.B(n_778),
.Y(n_1772)
);

OAI22xp5_ASAP7_75t_SL g1773 ( 
.A1(n_1699),
.A2(n_1327),
.B1(n_1333),
.B2(n_1324),
.Y(n_1773)
);

AO22x2_ASAP7_75t_L g1774 ( 
.A1(n_1633),
.A2(n_1229),
.B1(n_1188),
.B2(n_1348),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1551),
.B(n_1296),
.Y(n_1775)
);

OAI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1628),
.A2(n_1296),
.B1(n_1266),
.B2(n_1369),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1454),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1473),
.Y(n_1778)
);

INVx1_ASAP7_75t_SL g1779 ( 
.A(n_1597),
.Y(n_1779)
);

OAI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1628),
.A2(n_1378),
.B1(n_1384),
.B2(n_1372),
.Y(n_1780)
);

OAI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1628),
.A2(n_1398),
.B1(n_1401),
.B2(n_1395),
.Y(n_1781)
);

AOI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1498),
.A2(n_1299),
.B1(n_1289),
.B2(n_1403),
.Y(n_1782)
);

OAI22xp5_ASAP7_75t_SL g1783 ( 
.A1(n_1699),
.A2(n_1422),
.B1(n_1409),
.B2(n_1679),
.Y(n_1783)
);

AO22x2_ASAP7_75t_L g1784 ( 
.A1(n_1633),
.A2(n_757),
.B1(n_930),
.B2(n_929),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1494),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1597),
.B(n_933),
.Y(n_1786)
);

INVx1_ASAP7_75t_SL g1787 ( 
.A(n_1652),
.Y(n_1787)
);

INVx3_ASAP7_75t_L g1788 ( 
.A(n_1505),
.Y(n_1788)
);

OAI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1628),
.A2(n_1638),
.B1(n_1666),
.B2(n_1630),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1473),
.Y(n_1790)
);

AO22x2_ASAP7_75t_L g1791 ( 
.A1(n_1646),
.A2(n_938),
.B1(n_942),
.B2(n_939),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1498),
.A2(n_1557),
.B1(n_1565),
.B2(n_1662),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_L g1793 ( 
.A(n_1678),
.B(n_1648),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1650),
.B(n_947),
.Y(n_1794)
);

BUFx3_ASAP7_75t_L g1795 ( 
.A(n_1696),
.Y(n_1795)
);

OAI22xp33_ASAP7_75t_L g1796 ( 
.A1(n_1630),
.A2(n_672),
.B1(n_677),
.B2(n_665),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1494),
.Y(n_1797)
);

OAI22xp33_ASAP7_75t_R g1798 ( 
.A1(n_1682),
.A2(n_952),
.B1(n_955),
.B2(n_950),
.Y(n_1798)
);

OA22x2_ASAP7_75t_L g1799 ( 
.A1(n_1646),
.A2(n_958),
.B1(n_960),
.B2(n_956),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1494),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1494),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1650),
.B(n_961),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1655),
.B(n_962),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1494),
.Y(n_1804)
);

OAI22xp33_ASAP7_75t_L g1805 ( 
.A1(n_1630),
.A2(n_681),
.B1(n_683),
.B2(n_678),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1655),
.B(n_1544),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1655),
.B(n_965),
.Y(n_1807)
);

BUFx10_ASAP7_75t_L g1808 ( 
.A(n_1431),
.Y(n_1808)
);

AOI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1439),
.A2(n_536),
.B1(n_710),
.B2(n_688),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1460),
.B(n_684),
.Y(n_1810)
);

BUFx10_ASAP7_75t_L g1811 ( 
.A(n_1431),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1474),
.Y(n_1812)
);

OA22x2_ASAP7_75t_L g1813 ( 
.A1(n_1523),
.A2(n_969),
.B1(n_970),
.B2(n_966),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1544),
.B(n_971),
.Y(n_1814)
);

BUFx10_ASAP7_75t_L g1815 ( 
.A(n_1684),
.Y(n_1815)
);

AOI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1439),
.A2(n_695),
.B1(n_696),
.B2(n_694),
.Y(n_1816)
);

BUFx3_ASAP7_75t_L g1817 ( 
.A(n_1634),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_L g1818 ( 
.A(n_1620),
.B(n_698),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1662),
.B(n_973),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1565),
.B(n_974),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1565),
.B(n_1615),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1425),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1474),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1425),
.Y(n_1824)
);

INVx3_ASAP7_75t_L g1825 ( 
.A(n_1505),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1615),
.B(n_975),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1476),
.Y(n_1827)
);

BUFx6f_ASAP7_75t_L g1828 ( 
.A(n_1505),
.Y(n_1828)
);

AO22x2_ASAP7_75t_L g1829 ( 
.A1(n_1692),
.A2(n_977),
.B1(n_978),
.B2(n_976),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1432),
.Y(n_1830)
);

OAI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1620),
.A2(n_702),
.B1(n_703),
.B2(n_700),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1432),
.Y(n_1832)
);

OAI22xp33_ASAP7_75t_L g1833 ( 
.A1(n_1630),
.A2(n_714),
.B1(n_717),
.B2(n_709),
.Y(n_1833)
);

OAI22xp33_ASAP7_75t_SL g1834 ( 
.A1(n_1692),
.A2(n_719),
.B1(n_724),
.B2(n_718),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1436),
.Y(n_1835)
);

INVx3_ASAP7_75t_L g1836 ( 
.A(n_1525),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1476),
.Y(n_1837)
);

AOI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1439),
.A2(n_728),
.B1(n_733),
.B2(n_727),
.Y(n_1838)
);

CKINVDCx8_ASAP7_75t_R g1839 ( 
.A(n_1434),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1620),
.B(n_734),
.Y(n_1840)
);

OAI22xp33_ASAP7_75t_L g1841 ( 
.A1(n_1630),
.A2(n_738),
.B1(n_740),
.B2(n_737),
.Y(n_1841)
);

AOI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1557),
.A2(n_462),
.B1(n_467),
.B2(n_461),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1436),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1469),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1615),
.B(n_979),
.Y(n_1845)
);

AOI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1675),
.A2(n_481),
.B1(n_483),
.B2(n_468),
.Y(n_1846)
);

AOI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1675),
.A2(n_492),
.B1(n_494),
.B2(n_486),
.Y(n_1847)
);

AOI22xp5_ASAP7_75t_L g1848 ( 
.A1(n_1440),
.A2(n_510),
.B1(n_515),
.B2(n_502),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1487),
.Y(n_1849)
);

OAI22xp5_ASAP7_75t_SL g1850 ( 
.A1(n_1693),
.A2(n_747),
.B1(n_748),
.B2(n_745),
.Y(n_1850)
);

AO22x2_ASAP7_75t_L g1851 ( 
.A1(n_1704),
.A2(n_982),
.B1(n_989),
.B2(n_987),
.Y(n_1851)
);

AND2x6_ASAP7_75t_L g1852 ( 
.A(n_1622),
.B(n_507),
.Y(n_1852)
);

AOI22xp5_ASAP7_75t_L g1853 ( 
.A1(n_1440),
.A2(n_538),
.B1(n_540),
.B2(n_539),
.Y(n_1853)
);

AOI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1440),
.A2(n_542),
.B1(n_551),
.B2(n_543),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1469),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1478),
.Y(n_1856)
);

OAI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1622),
.A2(n_993),
.B1(n_994),
.B2(n_992),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1596),
.B(n_995),
.Y(n_1858)
);

NAND3x1_ASAP7_75t_L g1859 ( 
.A(n_1635),
.B(n_1003),
.C(n_996),
.Y(n_1859)
);

AOI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1483),
.A2(n_555),
.B1(n_559),
.B2(n_556),
.Y(n_1860)
);

AND2x2_ASAP7_75t_SL g1861 ( 
.A(n_1643),
.B(n_1005),
.Y(n_1861)
);

AO22x2_ASAP7_75t_L g1862 ( 
.A1(n_1704),
.A2(n_1022),
.B1(n_1023),
.B2(n_1014),
.Y(n_1862)
);

AO22x2_ASAP7_75t_L g1863 ( 
.A1(n_1706),
.A2(n_1029),
.B1(n_1030),
.B2(n_1026),
.Y(n_1863)
);

NAND3x1_ASAP7_75t_L g1864 ( 
.A(n_1635),
.B(n_1034),
.C(n_1032),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1637),
.B(n_1038),
.Y(n_1865)
);

OAI22xp33_ASAP7_75t_L g1866 ( 
.A1(n_1638),
.A2(n_1040),
.B1(n_1041),
.B2(n_1039),
.Y(n_1866)
);

OAI22xp5_ASAP7_75t_SL g1867 ( 
.A1(n_1643),
.A2(n_1047),
.B1(n_1048),
.B2(n_1046),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1478),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1487),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1479),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1483),
.B(n_1052),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1483),
.B(n_1055),
.Y(n_1872)
);

OAI22xp5_ASAP7_75t_SL g1873 ( 
.A1(n_1526),
.A2(n_1057),
.B1(n_1058),
.B2(n_1056),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1467),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1658),
.B(n_1061),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1467),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1479),
.Y(n_1877)
);

AOI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1500),
.A2(n_560),
.B1(n_572),
.B2(n_568),
.Y(n_1878)
);

AOI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1658),
.A2(n_580),
.B1(n_590),
.B2(n_587),
.Y(n_1879)
);

OAI22xp5_ASAP7_75t_SL g1880 ( 
.A1(n_1580),
.A2(n_1069),
.B1(n_1072),
.B2(n_1065),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1593),
.B(n_1074),
.Y(n_1881)
);

OA22x2_ASAP7_75t_L g1882 ( 
.A1(n_1629),
.A2(n_1076),
.B1(n_1077),
.B2(n_1075),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1658),
.B(n_1082),
.Y(n_1883)
);

NAND3x1_ASAP7_75t_L g1884 ( 
.A(n_1637),
.B(n_1084),
.C(n_1085),
.Y(n_1884)
);

AOI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1664),
.A2(n_595),
.B1(n_608),
.B2(n_598),
.Y(n_1885)
);

NOR2xp33_ASAP7_75t_L g1886 ( 
.A(n_1627),
.B(n_615),
.Y(n_1886)
);

OAI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1627),
.A2(n_628),
.B1(n_647),
.B2(n_632),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1664),
.B(n_1086),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1593),
.B(n_660),
.Y(n_1889)
);

AO22x2_ASAP7_75t_L g1890 ( 
.A1(n_1706),
.A2(n_1118),
.B1(n_1107),
.B2(n_1108),
.Y(n_1890)
);

OAI22xp5_ASAP7_75t_SL g1891 ( 
.A1(n_1684),
.A2(n_1529),
.B1(n_1492),
.B2(n_1669),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1481),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1481),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1467),
.Y(n_1894)
);

AO22x2_ASAP7_75t_L g1895 ( 
.A1(n_1709),
.A2(n_1107),
.B1(n_1108),
.B2(n_1105),
.Y(n_1895)
);

AO22x2_ASAP7_75t_L g1896 ( 
.A1(n_1709),
.A2(n_1111),
.B1(n_1105),
.B2(n_874),
.Y(n_1896)
);

AOI22xp5_ASAP7_75t_L g1897 ( 
.A1(n_1664),
.A2(n_662),
.B1(n_671),
.B2(n_667),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1671),
.B(n_1111),
.Y(n_1898)
);

OR2x6_ASAP7_75t_L g1899 ( 
.A(n_1690),
.B(n_822),
.Y(n_1899)
);

OAI22xp33_ASAP7_75t_L g1900 ( 
.A1(n_1638),
.A2(n_674),
.B1(n_680),
.B2(n_675),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1482),
.Y(n_1901)
);

BUFx2_ASAP7_75t_L g1902 ( 
.A(n_1637),
.Y(n_1902)
);

NAND3x1_ASAP7_75t_L g1903 ( 
.A(n_1626),
.B(n_10),
.C(n_11),
.Y(n_1903)
);

AO22x2_ASAP7_75t_L g1904 ( 
.A1(n_1665),
.A2(n_874),
.B1(n_897),
.B2(n_822),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1482),
.Y(n_1905)
);

OAI22xp33_ASAP7_75t_SL g1906 ( 
.A1(n_1665),
.A2(n_689),
.B1(n_691),
.B2(n_685),
.Y(n_1906)
);

INVx2_ASAP7_75t_SL g1907 ( 
.A(n_1634),
.Y(n_1907)
);

AOI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1671),
.A2(n_701),
.B1(n_706),
.B2(n_704),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1486),
.Y(n_1909)
);

OAI22xp33_ASAP7_75t_L g1910 ( 
.A1(n_1638),
.A2(n_712),
.B1(n_746),
.B2(n_716),
.Y(n_1910)
);

AO22x2_ASAP7_75t_L g1911 ( 
.A1(n_1672),
.A2(n_917),
.B1(n_936),
.B2(n_897),
.Y(n_1911)
);

INVx5_ASAP7_75t_L g1912 ( 
.A(n_1511),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1486),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1488),
.Y(n_1914)
);

AO22x2_ASAP7_75t_L g1915 ( 
.A1(n_1672),
.A2(n_936),
.B1(n_917),
.B2(n_13),
.Y(n_1915)
);

AO22x2_ASAP7_75t_L g1916 ( 
.A1(n_1674),
.A2(n_1680),
.B1(n_1685),
.B2(n_1677),
.Y(n_1916)
);

NOR2xp33_ASAP7_75t_L g1917 ( 
.A(n_1627),
.B(n_752),
.Y(n_1917)
);

OAI22xp33_ASAP7_75t_SL g1918 ( 
.A1(n_1674),
.A2(n_753),
.B1(n_13),
.B2(n_11),
.Y(n_1918)
);

AND2x2_ASAP7_75t_SL g1919 ( 
.A(n_1700),
.B(n_507),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1488),
.Y(n_1920)
);

AO22x2_ASAP7_75t_L g1921 ( 
.A1(n_1677),
.A2(n_15),
.B1(n_12),
.B2(n_14),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1671),
.B(n_12),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1491),
.Y(n_1923)
);

AOI22xp5_ASAP7_75t_L g1924 ( 
.A1(n_1582),
.A2(n_801),
.B1(n_813),
.B2(n_794),
.Y(n_1924)
);

INVx3_ASAP7_75t_L g1925 ( 
.A(n_1525),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1477),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1477),
.Y(n_1927)
);

AOI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1439),
.A2(n_801),
.B1(n_813),
.B2(n_794),
.Y(n_1928)
);

AOI22xp5_ASAP7_75t_L g1929 ( 
.A1(n_1439),
.A2(n_801),
.B1(n_813),
.B2(n_794),
.Y(n_1929)
);

OAI22xp5_ASAP7_75t_SL g1930 ( 
.A1(n_1669),
.A2(n_20),
.B1(n_17),
.B2(n_19),
.Y(n_1930)
);

OAI22xp33_ASAP7_75t_L g1931 ( 
.A1(n_1638),
.A2(n_22),
.B1(n_19),
.B2(n_21),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1513),
.B(n_21),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1477),
.Y(n_1933)
);

INVx3_ASAP7_75t_L g1934 ( 
.A(n_1525),
.Y(n_1934)
);

OR2x2_ASAP7_75t_L g1935 ( 
.A(n_1681),
.B(n_1689),
.Y(n_1935)
);

AO22x2_ASAP7_75t_L g1936 ( 
.A1(n_1680),
.A2(n_26),
.B1(n_23),
.B2(n_24),
.Y(n_1936)
);

AOI22xp5_ASAP7_75t_L g1937 ( 
.A1(n_1439),
.A2(n_1499),
.B1(n_1559),
.B2(n_1517),
.Y(n_1937)
);

AOI22xp5_ASAP7_75t_L g1938 ( 
.A1(n_1499),
.A2(n_801),
.B1(n_813),
.B2(n_794),
.Y(n_1938)
);

NOR2xp33_ASAP7_75t_L g1939 ( 
.A(n_1685),
.B(n_23),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1582),
.B(n_24),
.Y(n_1940)
);

OAI22xp5_ASAP7_75t_L g1941 ( 
.A1(n_1593),
.A2(n_30),
.B1(n_27),
.B2(n_28),
.Y(n_1941)
);

AOI22xp5_ASAP7_75t_L g1942 ( 
.A1(n_1499),
.A2(n_813),
.B1(n_878),
.B2(n_801),
.Y(n_1942)
);

NAND3x1_ASAP7_75t_L g1943 ( 
.A(n_1710),
.B(n_27),
.C(n_28),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1491),
.Y(n_1944)
);

INVx2_ASAP7_75t_SL g1945 ( 
.A(n_1634),
.Y(n_1945)
);

AOI22xp5_ASAP7_75t_L g1946 ( 
.A1(n_1499),
.A2(n_941),
.B1(n_1027),
.B2(n_878),
.Y(n_1946)
);

NOR2xp33_ASAP7_75t_L g1947 ( 
.A(n_1691),
.B(n_30),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1502),
.Y(n_1948)
);

AOI22xp5_ASAP7_75t_L g1949 ( 
.A1(n_1499),
.A2(n_941),
.B1(n_1027),
.B2(n_878),
.Y(n_1949)
);

NOR2xp33_ASAP7_75t_L g1950 ( 
.A(n_1691),
.B(n_1695),
.Y(n_1950)
);

AOI22xp5_ASAP7_75t_L g1951 ( 
.A1(n_1499),
.A2(n_941),
.B1(n_1027),
.B2(n_878),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1495),
.Y(n_1952)
);

INVx2_ASAP7_75t_SL g1953 ( 
.A(n_1634),
.Y(n_1953)
);

OAI22xp5_ASAP7_75t_SL g1954 ( 
.A1(n_1681),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_1954)
);

OR2x2_ASAP7_75t_L g1955 ( 
.A(n_1689),
.B(n_31),
.Y(n_1955)
);

AOI22xp5_ASAP7_75t_L g1956 ( 
.A1(n_1517),
.A2(n_1559),
.B1(n_1566),
.B2(n_1502),
.Y(n_1956)
);

AO22x2_ASAP7_75t_L g1957 ( 
.A1(n_1695),
.A2(n_35),
.B1(n_32),
.B2(n_34),
.Y(n_1957)
);

INVx2_ASAP7_75t_SL g1958 ( 
.A(n_1703),
.Y(n_1958)
);

OAI22xp5_ASAP7_75t_L g1959 ( 
.A1(n_1613),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_1959)
);

BUFx6f_ASAP7_75t_L g1960 ( 
.A(n_1525),
.Y(n_1960)
);

INVx3_ASAP7_75t_L g1961 ( 
.A(n_1525),
.Y(n_1961)
);

AOI22xp5_ASAP7_75t_L g1962 ( 
.A1(n_1517),
.A2(n_941),
.B1(n_1027),
.B2(n_878),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1502),
.Y(n_1963)
);

OAI22xp33_ASAP7_75t_L g1964 ( 
.A1(n_1666),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1495),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1537),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1537),
.Y(n_1967)
);

OAI22xp5_ASAP7_75t_SL g1968 ( 
.A1(n_1701),
.A2(n_1708),
.B1(n_1667),
.B2(n_1670),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1559),
.Y(n_1969)
);

AO22x2_ASAP7_75t_L g1970 ( 
.A1(n_1701),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_1970)
);

AOI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1582),
.A2(n_1027),
.B1(n_1070),
.B2(n_941),
.Y(n_1971)
);

INVx3_ASAP7_75t_L g1972 ( 
.A(n_1537),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1566),
.Y(n_1973)
);

AO22x2_ASAP7_75t_L g1974 ( 
.A1(n_1708),
.A2(n_42),
.B1(n_39),
.B2(n_40),
.Y(n_1974)
);

OR2x2_ASAP7_75t_L g1975 ( 
.A(n_1591),
.B(n_42),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1566),
.Y(n_1976)
);

OAI22xp33_ASAP7_75t_L g1977 ( 
.A1(n_1666),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_1977)
);

OAI22xp33_ASAP7_75t_L g1978 ( 
.A1(n_1666),
.A2(n_1711),
.B1(n_1683),
.B2(n_1702),
.Y(n_1978)
);

OAI22xp33_ASAP7_75t_L g1979 ( 
.A1(n_1666),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1503),
.B(n_1545),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1537),
.Y(n_1981)
);

AOI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1613),
.A2(n_1096),
.B1(n_1099),
.B2(n_1070),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1537),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1541),
.Y(n_1984)
);

AOI22xp5_ASAP7_75t_L g1985 ( 
.A1(n_1613),
.A2(n_1096),
.B1(n_1099),
.B2(n_1070),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1636),
.B(n_46),
.Y(n_1986)
);

AO22x2_ASAP7_75t_L g1987 ( 
.A1(n_1592),
.A2(n_1562),
.B1(n_1475),
.B2(n_1535),
.Y(n_1987)
);

AO22x2_ASAP7_75t_L g1988 ( 
.A1(n_1592),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1541),
.Y(n_1989)
);

AOI22xp5_ASAP7_75t_L g1990 ( 
.A1(n_1700),
.A2(n_1096),
.B1(n_1099),
.B2(n_1070),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1541),
.Y(n_1991)
);

OAI22xp33_ASAP7_75t_L g1992 ( 
.A1(n_1711),
.A2(n_50),
.B1(n_47),
.B2(n_49),
.Y(n_1992)
);

OAI22xp5_ASAP7_75t_SL g1993 ( 
.A1(n_1659),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1427),
.Y(n_1994)
);

OAI22xp33_ASAP7_75t_R g1995 ( 
.A1(n_1673),
.A2(n_54),
.B1(n_51),
.B2(n_53),
.Y(n_1995)
);

OAI22xp33_ASAP7_75t_L g1996 ( 
.A1(n_1711),
.A2(n_59),
.B1(n_54),
.B2(n_57),
.Y(n_1996)
);

OAI22xp33_ASAP7_75t_R g1997 ( 
.A1(n_1676),
.A2(n_66),
.B1(n_60),
.B2(n_65),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1583),
.B(n_60),
.Y(n_1998)
);

OAI22xp5_ASAP7_75t_L g1999 ( 
.A1(n_1599),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_1999)
);

AOI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1541),
.A2(n_1096),
.B1(n_1099),
.B2(n_1070),
.Y(n_2000)
);

OAI22xp33_ASAP7_75t_L g2001 ( 
.A1(n_1711),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_2001)
);

AOI22xp5_ASAP7_75t_L g2002 ( 
.A1(n_1541),
.A2(n_1549),
.B1(n_1554),
.B2(n_1547),
.Y(n_2002)
);

OAI22xp33_ASAP7_75t_L g2003 ( 
.A1(n_1711),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_2003)
);

OR2x6_ASAP7_75t_L g2004 ( 
.A(n_1703),
.B(n_1096),
.Y(n_2004)
);

OR2x2_ASAP7_75t_L g2005 ( 
.A(n_1720),
.B(n_1649),
.Y(n_2005)
);

INVx2_ASAP7_75t_SL g2006 ( 
.A(n_2004),
.Y(n_2006)
);

INVx1_ASAP7_75t_SL g2007 ( 
.A(n_1779),
.Y(n_2007)
);

BUFx3_ASAP7_75t_L g2008 ( 
.A(n_1795),
.Y(n_2008)
);

INVx2_ASAP7_75t_SL g2009 ( 
.A(n_2004),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1822),
.Y(n_2010)
);

AND2x4_ASAP7_75t_L g2011 ( 
.A(n_1821),
.B(n_1579),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1824),
.Y(n_2012)
);

INVx3_ASAP7_75t_L g2013 ( 
.A(n_1828),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1830),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1832),
.Y(n_2015)
);

OAI21xp33_ASAP7_75t_SL g2016 ( 
.A1(n_1919),
.A2(n_1514),
.B(n_1507),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1835),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1746),
.B(n_1611),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1843),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1793),
.B(n_1611),
.Y(n_2020)
);

AOI22xp33_ASAP7_75t_L g2021 ( 
.A1(n_1861),
.A2(n_1600),
.B1(n_1579),
.B2(n_1592),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1844),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1855),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1713),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1856),
.Y(n_2025)
);

INVx3_ASAP7_75t_L g2026 ( 
.A(n_1828),
.Y(n_2026)
);

AOI22xp33_ASAP7_75t_L g2027 ( 
.A1(n_1867),
.A2(n_1600),
.B1(n_1590),
.B2(n_1588),
.Y(n_2027)
);

AOI22xp33_ASAP7_75t_L g2028 ( 
.A1(n_1798),
.A2(n_1590),
.B1(n_1588),
.B2(n_1589),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_SL g2029 ( 
.A(n_1770),
.B(n_1612),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_SL g2030 ( 
.A(n_1978),
.B(n_1612),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1713),
.Y(n_2031)
);

AOI22xp33_ASAP7_75t_L g2032 ( 
.A1(n_1767),
.A2(n_1590),
.B1(n_1589),
.B2(n_1581),
.Y(n_2032)
);

NOR3xp33_ASAP7_75t_L g2033 ( 
.A(n_1734),
.B(n_1714),
.C(n_1740),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1724),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1810),
.B(n_1612),
.Y(n_2035)
);

INVx4_ASAP7_75t_L g2036 ( 
.A(n_1912),
.Y(n_2036)
);

BUFx3_ASAP7_75t_L g2037 ( 
.A(n_1751),
.Y(n_2037)
);

INVx4_ASAP7_75t_L g2038 ( 
.A(n_1912),
.Y(n_2038)
);

INVx3_ASAP7_75t_L g2039 ( 
.A(n_1828),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1950),
.B(n_1612),
.Y(n_2040)
);

NOR2xp33_ASAP7_75t_L g2041 ( 
.A(n_1712),
.B(n_1703),
.Y(n_2041)
);

BUFx3_ASAP7_75t_L g2042 ( 
.A(n_1759),
.Y(n_2042)
);

OAI21xp33_ASAP7_75t_SL g2043 ( 
.A1(n_1956),
.A2(n_1514),
.B(n_1507),
.Y(n_2043)
);

XOR2xp5_ASAP7_75t_L g2044 ( 
.A(n_1773),
.B(n_1987),
.Y(n_2044)
);

BUFx6f_ASAP7_75t_L g2045 ( 
.A(n_1960),
.Y(n_2045)
);

INVxp67_ASAP7_75t_SL g2046 ( 
.A(n_2002),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1726),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1735),
.Y(n_2048)
);

OAI22xp33_ASAP7_75t_L g2049 ( 
.A1(n_1712),
.A2(n_1715),
.B1(n_1768),
.B2(n_1731),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1735),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1718),
.B(n_1612),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_1868),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1870),
.Y(n_2053)
);

INVx4_ASAP7_75t_L g2054 ( 
.A(n_1912),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1877),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1738),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1892),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1893),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1901),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_1806),
.B(n_1820),
.Y(n_2060)
);

NOR2xp33_ASAP7_75t_L g2061 ( 
.A(n_1716),
.B(n_1703),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1738),
.Y(n_2062)
);

BUFx3_ASAP7_75t_L g2063 ( 
.A(n_1759),
.Y(n_2063)
);

AND2x6_ASAP7_75t_L g2064 ( 
.A(n_1937),
.B(n_1642),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1905),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1819),
.B(n_1614),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1792),
.B(n_1614),
.Y(n_2067)
);

OAI22xp33_ASAP7_75t_L g2068 ( 
.A1(n_1715),
.A2(n_1723),
.B1(n_1754),
.B2(n_1775),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1909),
.Y(n_2069)
);

OAI22xp33_ASAP7_75t_L g2070 ( 
.A1(n_1736),
.A2(n_1737),
.B1(n_1865),
.B2(n_1758),
.Y(n_2070)
);

INVx2_ASAP7_75t_SL g2071 ( 
.A(n_1772),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1777),
.Y(n_2072)
);

BUFx6f_ASAP7_75t_L g2073 ( 
.A(n_1960),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1913),
.Y(n_2074)
);

INVx4_ASAP7_75t_L g2075 ( 
.A(n_1960),
.Y(n_2075)
);

INVx4_ASAP7_75t_L g2076 ( 
.A(n_1743),
.Y(n_2076)
);

INVx6_ASAP7_75t_L g2077 ( 
.A(n_1817),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_1826),
.B(n_1464),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1777),
.Y(n_2079)
);

INVx5_ASAP7_75t_L g2080 ( 
.A(n_1852),
.Y(n_2080)
);

BUFx10_ASAP7_75t_L g2081 ( 
.A(n_1728),
.Y(n_2081)
);

NOR2xp33_ASAP7_75t_L g2082 ( 
.A(n_1722),
.B(n_1621),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1778),
.Y(n_2083)
);

BUFx6f_ASAP7_75t_L g2084 ( 
.A(n_1717),
.Y(n_2084)
);

CKINVDCx20_ASAP7_75t_R g2085 ( 
.A(n_1839),
.Y(n_2085)
);

INVx6_ASAP7_75t_L g2086 ( 
.A(n_1899),
.Y(n_2086)
);

BUFx6f_ASAP7_75t_L g2087 ( 
.A(n_1717),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1778),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1790),
.Y(n_2089)
);

NAND3xp33_ASAP7_75t_L g2090 ( 
.A(n_1782),
.B(n_1686),
.C(n_1553),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1914),
.Y(n_2091)
);

INVx4_ASAP7_75t_L g2092 ( 
.A(n_1749),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_SL g2093 ( 
.A(n_1765),
.B(n_1614),
.Y(n_2093)
);

AND2x6_ASAP7_75t_L g2094 ( 
.A(n_1937),
.B(n_1642),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1814),
.B(n_1614),
.Y(n_2095)
);

AOI22xp33_ASAP7_75t_L g2096 ( 
.A1(n_1932),
.A2(n_1590),
.B1(n_1601),
.B2(n_1581),
.Y(n_2096)
);

XOR2x2_ASAP7_75t_L g2097 ( 
.A(n_1980),
.B(n_1660),
.Y(n_2097)
);

NOR2xp33_ASAP7_75t_L g2098 ( 
.A(n_1730),
.B(n_1631),
.Y(n_2098)
);

INVx4_ASAP7_75t_L g2099 ( 
.A(n_1749),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_SL g2100 ( 
.A(n_1789),
.B(n_1614),
.Y(n_2100)
);

INVx3_ASAP7_75t_L g2101 ( 
.A(n_1788),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_1920),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1923),
.Y(n_2103)
);

INVx3_ASAP7_75t_L g2104 ( 
.A(n_1788),
.Y(n_2104)
);

INVx2_ASAP7_75t_SL g2105 ( 
.A(n_1772),
.Y(n_2105)
);

NAND2xp33_ASAP7_75t_L g2106 ( 
.A(n_1956),
.B(n_1599),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1812),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_1845),
.B(n_1464),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1871),
.B(n_1618),
.Y(n_2109)
);

INVx11_ASAP7_75t_L g2110 ( 
.A(n_1728),
.Y(n_2110)
);

INVx3_ASAP7_75t_L g2111 ( 
.A(n_1825),
.Y(n_2111)
);

INVx2_ASAP7_75t_SL g2112 ( 
.A(n_1899),
.Y(n_2112)
);

INVx3_ASAP7_75t_L g2113 ( 
.A(n_1825),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_SL g2114 ( 
.A(n_1739),
.B(n_1618),
.Y(n_2114)
);

NAND2xp33_ASAP7_75t_R g2115 ( 
.A(n_1769),
.B(n_1642),
.Y(n_2115)
);

BUFx3_ASAP7_75t_L g2116 ( 
.A(n_1958),
.Y(n_2116)
);

INVx2_ASAP7_75t_SL g2117 ( 
.A(n_1902),
.Y(n_2117)
);

CKINVDCx5p33_ASAP7_75t_R g2118 ( 
.A(n_1808),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1944),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1823),
.Y(n_2120)
);

AND2x6_ASAP7_75t_L g2121 ( 
.A(n_2002),
.B(n_1647),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1952),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_1965),
.Y(n_2123)
);

BUFx6f_ASAP7_75t_L g2124 ( 
.A(n_1836),
.Y(n_2124)
);

BUFx2_ASAP7_75t_L g2125 ( 
.A(n_1935),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_1803),
.B(n_1470),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1823),
.Y(n_2127)
);

INVxp33_ASAP7_75t_SL g2128 ( 
.A(n_1771),
.Y(n_2128)
);

INVx2_ASAP7_75t_SL g2129 ( 
.A(n_1719),
.Y(n_2129)
);

INVx1_ASAP7_75t_SL g2130 ( 
.A(n_1787),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1827),
.Y(n_2131)
);

INVx2_ASAP7_75t_SL g2132 ( 
.A(n_1721),
.Y(n_2132)
);

NOR2xp33_ASAP7_75t_L g2133 ( 
.A(n_1747),
.B(n_1632),
.Y(n_2133)
);

INVx2_ASAP7_75t_SL g2134 ( 
.A(n_1807),
.Y(n_2134)
);

AND2x2_ASAP7_75t_SL g2135 ( 
.A(n_1809),
.B(n_1733),
.Y(n_2135)
);

INVx3_ASAP7_75t_L g2136 ( 
.A(n_1836),
.Y(n_2136)
);

OAI22xp5_ASAP7_75t_L g2137 ( 
.A1(n_1827),
.A2(n_1510),
.B1(n_1516),
.B2(n_1512),
.Y(n_2137)
);

CKINVDCx5p33_ASAP7_75t_R g2138 ( 
.A(n_1808),
.Y(n_2138)
);

INVx3_ASAP7_75t_L g2139 ( 
.A(n_1925),
.Y(n_2139)
);

BUFx3_ASAP7_75t_L g2140 ( 
.A(n_1811),
.Y(n_2140)
);

INVxp67_ASAP7_75t_L g2141 ( 
.A(n_1748),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_SL g2142 ( 
.A(n_1729),
.B(n_1618),
.Y(n_2142)
);

INVx5_ASAP7_75t_L g2143 ( 
.A(n_1852),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1727),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_1744),
.Y(n_2145)
);

NOR2xp33_ASAP7_75t_L g2146 ( 
.A(n_1776),
.B(n_1640),
.Y(n_2146)
);

OAI22xp5_ASAP7_75t_L g2147 ( 
.A1(n_1837),
.A2(n_1510),
.B1(n_1516),
.B2(n_1512),
.Y(n_2147)
);

BUFx10_ASAP7_75t_L g2148 ( 
.A(n_1818),
.Y(n_2148)
);

INVx3_ASAP7_75t_L g2149 ( 
.A(n_1925),
.Y(n_2149)
);

BUFx6f_ASAP7_75t_L g2150 ( 
.A(n_1934),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1837),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_1745),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1849),
.Y(n_2153)
);

OR2x6_ASAP7_75t_L g2154 ( 
.A(n_1907),
.B(n_1688),
.Y(n_2154)
);

BUFx3_ASAP7_75t_L g2155 ( 
.A(n_1811),
.Y(n_2155)
);

INVx2_ASAP7_75t_SL g2156 ( 
.A(n_1875),
.Y(n_2156)
);

INVx4_ASAP7_75t_L g2157 ( 
.A(n_1934),
.Y(n_2157)
);

CKINVDCx5p33_ASAP7_75t_R g2158 ( 
.A(n_1815),
.Y(n_2158)
);

BUFx3_ASAP7_75t_L g2159 ( 
.A(n_1815),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_SL g2160 ( 
.A(n_1757),
.B(n_1618),
.Y(n_2160)
);

AOI22xp33_ASAP7_75t_L g2161 ( 
.A1(n_1761),
.A2(n_1733),
.B1(n_1851),
.B2(n_1829),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_1755),
.Y(n_2162)
);

BUFx3_ASAP7_75t_L g2163 ( 
.A(n_1961),
.Y(n_2163)
);

AND2x2_ASAP7_75t_SL g2164 ( 
.A(n_1809),
.B(n_1663),
.Y(n_2164)
);

INVx3_ASAP7_75t_L g2165 ( 
.A(n_1961),
.Y(n_2165)
);

AOI22xp33_ASAP7_75t_L g2166 ( 
.A1(n_1829),
.A2(n_1590),
.B1(n_1602),
.B2(n_1601),
.Y(n_2166)
);

INVxp33_ASAP7_75t_L g2167 ( 
.A(n_1750),
.Y(n_2167)
);

INVx3_ASAP7_75t_L g2168 ( 
.A(n_1972),
.Y(n_2168)
);

INVx2_ASAP7_75t_SL g2169 ( 
.A(n_1883),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_1872),
.B(n_1618),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_1874),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1874),
.Y(n_2172)
);

INVx3_ASAP7_75t_L g2173 ( 
.A(n_1972),
.Y(n_2173)
);

BUFx6f_ASAP7_75t_L g2174 ( 
.A(n_1785),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1869),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1876),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_SL g2177 ( 
.A(n_1968),
.B(n_1599),
.Y(n_2177)
);

INVxp33_ASAP7_75t_L g2178 ( 
.A(n_1760),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_1876),
.Y(n_2179)
);

BUFx10_ASAP7_75t_L g2180 ( 
.A(n_1840),
.Y(n_2180)
);

INVx2_ASAP7_75t_SL g2181 ( 
.A(n_1898),
.Y(n_2181)
);

BUFx6f_ASAP7_75t_L g2182 ( 
.A(n_1797),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_1894),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_1894),
.Y(n_2184)
);

AND2x4_ASAP7_75t_L g2185 ( 
.A(n_1940),
.B(n_1922),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_1926),
.Y(n_2186)
);

AOI22xp33_ASAP7_75t_L g2187 ( 
.A1(n_1851),
.A2(n_1608),
.B1(n_1610),
.B2(n_1602),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1926),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_1927),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_1927),
.Y(n_2190)
);

OAI22x1_ASAP7_75t_L g2191 ( 
.A1(n_1752),
.A2(n_1651),
.B1(n_1645),
.B2(n_1688),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_1933),
.Y(n_2192)
);

AOI22xp33_ASAP7_75t_L g2193 ( 
.A1(n_1862),
.A2(n_1610),
.B1(n_1608),
.B2(n_1549),
.Y(n_2193)
);

NOR2xp33_ASAP7_75t_L g2194 ( 
.A(n_1764),
.B(n_1688),
.Y(n_2194)
);

BUFx3_ASAP7_75t_L g2195 ( 
.A(n_1945),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_1933),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_1794),
.B(n_1470),
.Y(n_2197)
);

OR2x6_ASAP7_75t_L g2198 ( 
.A(n_1953),
.B(n_1663),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_1948),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_1802),
.B(n_1599),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_1948),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_1963),
.Y(n_2202)
);

INVx1_ASAP7_75t_SL g2203 ( 
.A(n_1786),
.Y(n_2203)
);

INVx3_ASAP7_75t_L g2204 ( 
.A(n_1800),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1963),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1969),
.Y(n_2206)
);

BUFx2_ASAP7_75t_L g2207 ( 
.A(n_1858),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_1998),
.B(n_1599),
.Y(n_2208)
);

AOI22xp5_ASAP7_75t_L g2209 ( 
.A1(n_1916),
.A2(n_1603),
.B1(n_1508),
.B2(n_1647),
.Y(n_2209)
);

INVx2_ASAP7_75t_SL g2210 ( 
.A(n_1888),
.Y(n_2210)
);

AOI22xp5_ASAP7_75t_L g2211 ( 
.A1(n_1916),
.A2(n_1653),
.B1(n_1647),
.B2(n_1609),
.Y(n_2211)
);

INVx3_ASAP7_75t_L g2212 ( 
.A(n_1801),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_1969),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1973),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_1791),
.B(n_1563),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1973),
.Y(n_2216)
);

AOI22xp33_ASAP7_75t_L g2217 ( 
.A1(n_1862),
.A2(n_1549),
.B1(n_1554),
.B2(n_1547),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_1976),
.Y(n_2218)
);

INVx2_ASAP7_75t_L g2219 ( 
.A(n_1976),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_1791),
.B(n_1563),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1881),
.Y(n_2221)
);

INVx2_ASAP7_75t_SL g2222 ( 
.A(n_1896),
.Y(n_2222)
);

INVx1_ASAP7_75t_SL g2223 ( 
.A(n_1955),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1994),
.Y(n_2224)
);

BUFx6f_ASAP7_75t_L g2225 ( 
.A(n_1804),
.Y(n_2225)
);

XNOR2xp5_ASAP7_75t_L g2226 ( 
.A(n_1987),
.B(n_1445),
.Y(n_2226)
);

BUFx3_ASAP7_75t_L g2227 ( 
.A(n_1966),
.Y(n_2227)
);

AOI22xp33_ASAP7_75t_SL g2228 ( 
.A1(n_1766),
.A2(n_1459),
.B1(n_1553),
.B2(n_1585),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_1895),
.B(n_1583),
.Y(n_2229)
);

INVx3_ASAP7_75t_L g2230 ( 
.A(n_1967),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_SL g2231 ( 
.A(n_1796),
.B(n_1653),
.Y(n_2231)
);

AND3x2_ASAP7_75t_L g2232 ( 
.A(n_1986),
.B(n_1572),
.C(n_1686),
.Y(n_2232)
);

BUFx6f_ASAP7_75t_L g2233 ( 
.A(n_1981),
.Y(n_2233)
);

INVx6_ASAP7_75t_L g2234 ( 
.A(n_1852),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_1886),
.B(n_1522),
.Y(n_2235)
);

INVx4_ASAP7_75t_L g2236 ( 
.A(n_1852),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1994),
.Y(n_2237)
);

NOR2xp33_ASAP7_75t_L g2238 ( 
.A(n_1780),
.B(n_1663),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1983),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1799),
.Y(n_2240)
);

BUFx6f_ASAP7_75t_L g2241 ( 
.A(n_1984),
.Y(n_2241)
);

AOI22xp5_ASAP7_75t_L g2242 ( 
.A1(n_1873),
.A2(n_1653),
.B1(n_1607),
.B2(n_1686),
.Y(n_2242)
);

INVx3_ASAP7_75t_L g2243 ( 
.A(n_1989),
.Y(n_2243)
);

AND2x6_ASAP7_75t_L g2244 ( 
.A(n_1928),
.B(n_1584),
.Y(n_2244)
);

OR2x2_ASAP7_75t_L g2245 ( 
.A(n_1781),
.B(n_1536),
.Y(n_2245)
);

CKINVDCx20_ASAP7_75t_R g2246 ( 
.A(n_1783),
.Y(n_2246)
);

INVx1_ASAP7_75t_SL g2247 ( 
.A(n_1774),
.Y(n_2247)
);

NAND2xp33_ASAP7_75t_L g2248 ( 
.A(n_1889),
.B(n_1512),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_1991),
.Y(n_2249)
);

INVx1_ASAP7_75t_SL g2250 ( 
.A(n_1774),
.Y(n_2250)
);

NOR2xp33_ASAP7_75t_L g2251 ( 
.A(n_1752),
.B(n_1758),
.Y(n_2251)
);

NOR2xp33_ASAP7_75t_SL g2252 ( 
.A(n_1891),
.B(n_1459),
.Y(n_2252)
);

NOR2xp33_ASAP7_75t_L g2253 ( 
.A(n_1842),
.B(n_1459),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_1917),
.B(n_1560),
.Y(n_2254)
);

INVx1_ASAP7_75t_SL g2255 ( 
.A(n_1880),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1896),
.Y(n_2256)
);

NOR2xp33_ASAP7_75t_L g2257 ( 
.A(n_1753),
.B(n_1553),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1904),
.Y(n_2258)
);

OAI22xp33_ASAP7_75t_SL g2259 ( 
.A1(n_1995),
.A2(n_1997),
.B1(n_1975),
.B2(n_1838),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_1784),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_1904),
.Y(n_2261)
);

INVx2_ASAP7_75t_SL g2262 ( 
.A(n_1895),
.Y(n_2262)
);

INVx4_ASAP7_75t_L g2263 ( 
.A(n_1915),
.Y(n_2263)
);

AOI21x1_ASAP7_75t_L g2264 ( 
.A1(n_1911),
.A2(n_1605),
.B(n_1586),
.Y(n_2264)
);

OR2x6_ASAP7_75t_L g2265 ( 
.A(n_1859),
.B(n_1584),
.Y(n_2265)
);

OR2x2_ASAP7_75t_L g2266 ( 
.A(n_1831),
.B(n_1438),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_1784),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1890),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_SL g2269 ( 
.A(n_1805),
.B(n_1455),
.Y(n_2269)
);

OAI22xp5_ASAP7_75t_SL g2270 ( 
.A1(n_1850),
.A2(n_1572),
.B1(n_1448),
.B2(n_1585),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_1939),
.B(n_1450),
.Y(n_2271)
);

INVx2_ASAP7_75t_SL g2272 ( 
.A(n_1890),
.Y(n_2272)
);

INVxp33_ASAP7_75t_SL g2273 ( 
.A(n_1762),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_1911),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_SL g2275 ( 
.A(n_1833),
.B(n_1455),
.Y(n_2275)
);

INVx3_ASAP7_75t_L g2276 ( 
.A(n_1915),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_1863),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1962),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2000),
.Y(n_2279)
);

OR2x2_ASAP7_75t_L g2280 ( 
.A(n_1857),
.B(n_1468),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_1962),
.Y(n_2281)
);

AOI22xp33_ASAP7_75t_L g2282 ( 
.A1(n_1863),
.A2(n_1549),
.B1(n_1554),
.B2(n_1547),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2000),
.Y(n_2283)
);

CKINVDCx11_ASAP7_75t_R g2284 ( 
.A(n_1941),
.Y(n_2284)
);

INVx4_ASAP7_75t_L g2285 ( 
.A(n_1988),
.Y(n_2285)
);

BUFx3_ASAP7_75t_L g2286 ( 
.A(n_1813),
.Y(n_2286)
);

OR2x2_ASAP7_75t_L g2287 ( 
.A(n_1879),
.B(n_1587),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_1947),
.B(n_1587),
.Y(n_2288)
);

INVx3_ASAP7_75t_L g2289 ( 
.A(n_1864),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_2171),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_SL g2291 ( 
.A(n_2049),
.B(n_1510),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2171),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2060),
.Y(n_2293)
);

AOI22xp5_ASAP7_75t_L g2294 ( 
.A1(n_2255),
.A2(n_1585),
.B1(n_1841),
.B2(n_1878),
.Y(n_2294)
);

AND2x4_ASAP7_75t_L g2295 ( 
.A(n_2011),
.B(n_2060),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_2172),
.Y(n_2296)
);

OR2x6_ASAP7_75t_L g2297 ( 
.A(n_2086),
.B(n_1766),
.Y(n_2297)
);

INVx2_ASAP7_75t_SL g2298 ( 
.A(n_2081),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2126),
.Y(n_2299)
);

NAND2x1p5_ASAP7_75t_L g2300 ( 
.A(n_2036),
.B(n_1547),
.Y(n_2300)
);

NOR2xp33_ASAP7_75t_L g2301 ( 
.A(n_2167),
.B(n_1725),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2126),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_2172),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2078),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_L g2305 ( 
.A(n_2020),
.B(n_1866),
.Y(n_2305)
);

NOR2xp33_ASAP7_75t_L g2306 ( 
.A(n_2167),
.B(n_2178),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2078),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2108),
.Y(n_2308)
);

AND2x4_ASAP7_75t_L g2309 ( 
.A(n_2011),
.B(n_1594),
.Y(n_2309)
);

AND2x4_ASAP7_75t_L g2310 ( 
.A(n_2008),
.B(n_1595),
.Y(n_2310)
);

AND2x2_ASAP7_75t_L g2311 ( 
.A(n_2203),
.B(n_2207),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2179),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2179),
.Y(n_2313)
);

NOR2xp33_ASAP7_75t_L g2314 ( 
.A(n_2178),
.B(n_2128),
.Y(n_2314)
);

HB1xp67_ASAP7_75t_L g2315 ( 
.A(n_2207),
.Y(n_2315)
);

CKINVDCx16_ASAP7_75t_R g2316 ( 
.A(n_2085),
.Y(n_2316)
);

OAI21xp33_ASAP7_75t_L g2317 ( 
.A1(n_2082),
.A2(n_1897),
.B(n_1885),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2108),
.Y(n_2318)
);

NOR2xp33_ASAP7_75t_L g2319 ( 
.A(n_2128),
.B(n_2018),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2024),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2031),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2183),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_2183),
.Y(n_2323)
);

AND2x4_ASAP7_75t_L g2324 ( 
.A(n_2008),
.B(n_1595),
.Y(n_2324)
);

OR2x2_ASAP7_75t_L g2325 ( 
.A(n_2125),
.B(n_1598),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_2184),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2034),
.Y(n_2327)
);

NOR2x1p5_ASAP7_75t_L g2328 ( 
.A(n_2140),
.B(n_1485),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_2184),
.Y(n_2329)
);

INVx2_ASAP7_75t_SL g2330 ( 
.A(n_2081),
.Y(n_2330)
);

HB1xp67_ASAP7_75t_L g2331 ( 
.A(n_2007),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_2194),
.B(n_1598),
.Y(n_2332)
);

AND2x4_ASAP7_75t_L g2333 ( 
.A(n_2156),
.B(n_1573),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2197),
.B(n_1521),
.Y(n_2334)
);

INVx4_ASAP7_75t_L g2335 ( 
.A(n_2110),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_2186),
.Y(n_2336)
);

BUFx6f_ASAP7_75t_L g2337 ( 
.A(n_2045),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2083),
.Y(n_2338)
);

NOR2xp33_ASAP7_75t_L g2339 ( 
.A(n_2068),
.B(n_1616),
.Y(n_2339)
);

INVx3_ASAP7_75t_L g2340 ( 
.A(n_2036),
.Y(n_2340)
);

INVxp67_ASAP7_75t_L g2341 ( 
.A(n_2125),
.Y(n_2341)
);

AOI22x1_ASAP7_75t_L g2342 ( 
.A1(n_2092),
.A2(n_1516),
.B1(n_1619),
.B2(n_1568),
.Y(n_2342)
);

NOR2xp33_ASAP7_75t_L g2343 ( 
.A(n_2041),
.B(n_1741),
.Y(n_2343)
);

INVx2_ASAP7_75t_SL g2344 ( 
.A(n_2081),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2088),
.Y(n_2345)
);

BUFx3_ASAP7_75t_L g2346 ( 
.A(n_2085),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2229),
.B(n_1882),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2061),
.B(n_1908),
.Y(n_2348)
);

OAI221xp5_ASAP7_75t_L g2349 ( 
.A1(n_2146),
.A2(n_1954),
.B1(n_1930),
.B2(n_1993),
.C(n_1816),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_2186),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_2098),
.B(n_1485),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_2188),
.Y(n_2352)
);

AND2x2_ASAP7_75t_L g2353 ( 
.A(n_2229),
.B(n_1763),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2133),
.B(n_1848),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2089),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2188),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2156),
.B(n_1853),
.Y(n_2357)
);

INVx2_ASAP7_75t_SL g2358 ( 
.A(n_2110),
.Y(n_2358)
);

BUFx6f_ASAP7_75t_L g2359 ( 
.A(n_2045),
.Y(n_2359)
);

INVx3_ASAP7_75t_L g2360 ( 
.A(n_2036),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_2189),
.Y(n_2361)
);

NOR2xp33_ASAP7_75t_L g2362 ( 
.A(n_2141),
.B(n_1742),
.Y(n_2362)
);

CKINVDCx5p33_ASAP7_75t_R g2363 ( 
.A(n_2118),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2107),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2127),
.Y(n_2365)
);

BUFx6f_ASAP7_75t_L g2366 ( 
.A(n_2045),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2151),
.Y(n_2367)
);

AND2x4_ASAP7_75t_L g2368 ( 
.A(n_2169),
.B(n_1574),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2169),
.B(n_1854),
.Y(n_2369)
);

AOI22xp5_ASAP7_75t_L g2370 ( 
.A1(n_2238),
.A2(n_1884),
.B1(n_1988),
.B2(n_1903),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_2189),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2190),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2153),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2047),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2190),
.Y(n_2375)
);

INVx3_ASAP7_75t_L g2376 ( 
.A(n_2038),
.Y(n_2376)
);

AND2x6_ASAP7_75t_L g2377 ( 
.A(n_2276),
.B(n_1928),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2047),
.Y(n_2378)
);

BUFx6f_ASAP7_75t_L g2379 ( 
.A(n_2045),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_2192),
.Y(n_2380)
);

OR2x2_ASAP7_75t_L g2381 ( 
.A(n_2005),
.B(n_1575),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2048),
.Y(n_2382)
);

INVx4_ASAP7_75t_L g2383 ( 
.A(n_2086),
.Y(n_2383)
);

AND2x6_ASAP7_75t_L g2384 ( 
.A(n_2276),
.B(n_1929),
.Y(n_2384)
);

OAI22xp5_ASAP7_75t_L g2385 ( 
.A1(n_2164),
.A2(n_1838),
.B1(n_1816),
.B2(n_1860),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2048),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_2192),
.Y(n_2387)
);

AND2x6_ASAP7_75t_L g2388 ( 
.A(n_2276),
.B(n_2289),
.Y(n_2388)
);

CKINVDCx20_ASAP7_75t_R g2389 ( 
.A(n_2246),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_2196),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2050),
.Y(n_2391)
);

INVxp67_ASAP7_75t_L g2392 ( 
.A(n_2134),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2050),
.Y(n_2393)
);

BUFx2_ASAP7_75t_L g2394 ( 
.A(n_2037),
.Y(n_2394)
);

INVx6_ASAP7_75t_L g2395 ( 
.A(n_2086),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2056),
.Y(n_2396)
);

AO22x2_ASAP7_75t_L g2397 ( 
.A1(n_2285),
.A2(n_1763),
.B1(n_1756),
.B2(n_1921),
.Y(n_2397)
);

INVxp67_ASAP7_75t_L g2398 ( 
.A(n_2130),
.Y(n_2398)
);

BUFx6f_ASAP7_75t_L g2399 ( 
.A(n_2045),
.Y(n_2399)
);

INVx3_ASAP7_75t_L g2400 ( 
.A(n_2038),
.Y(n_2400)
);

INVx3_ASAP7_75t_L g2401 ( 
.A(n_2038),
.Y(n_2401)
);

AND2x6_ASAP7_75t_L g2402 ( 
.A(n_2289),
.B(n_1929),
.Y(n_2402)
);

BUFx6f_ASAP7_75t_L g2403 ( 
.A(n_2073),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_SL g2404 ( 
.A(n_2164),
.B(n_1547),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_2196),
.Y(n_2405)
);

AND2x4_ASAP7_75t_L g2406 ( 
.A(n_2076),
.B(n_1604),
.Y(n_2406)
);

NAND2x1p5_ASAP7_75t_L g2407 ( 
.A(n_2054),
.B(n_1549),
.Y(n_2407)
);

INVx2_ASAP7_75t_L g2408 ( 
.A(n_2199),
.Y(n_2408)
);

HB1xp67_ASAP7_75t_L g2409 ( 
.A(n_2210),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_2181),
.B(n_2210),
.Y(n_2410)
);

INVx4_ASAP7_75t_L g2411 ( 
.A(n_2086),
.Y(n_2411)
);

CKINVDCx5p33_ASAP7_75t_R g2412 ( 
.A(n_2118),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_2161),
.B(n_1606),
.Y(n_2413)
);

BUFx6f_ASAP7_75t_L g2414 ( 
.A(n_2073),
.Y(n_2414)
);

INVx2_ASAP7_75t_L g2415 ( 
.A(n_2199),
.Y(n_2415)
);

BUFx3_ASAP7_75t_L g2416 ( 
.A(n_2037),
.Y(n_2416)
);

AND2x4_ASAP7_75t_L g2417 ( 
.A(n_2076),
.B(n_1437),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2062),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2072),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2201),
.Y(n_2420)
);

INVx6_ASAP7_75t_L g2421 ( 
.A(n_2076),
.Y(n_2421)
);

OAI22xp5_ASAP7_75t_L g2422 ( 
.A1(n_2288),
.A2(n_1519),
.B1(n_1511),
.B2(n_1931),
.Y(n_2422)
);

BUFx6f_ASAP7_75t_L g2423 ( 
.A(n_2073),
.Y(n_2423)
);

AND2x4_ASAP7_75t_L g2424 ( 
.A(n_2112),
.B(n_2071),
.Y(n_2424)
);

BUFx6f_ASAP7_75t_L g2425 ( 
.A(n_2073),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_SL g2426 ( 
.A(n_2043),
.B(n_1554),
.Y(n_2426)
);

BUFx6f_ASAP7_75t_L g2427 ( 
.A(n_2073),
.Y(n_2427)
);

AND2x4_ASAP7_75t_L g2428 ( 
.A(n_2112),
.B(n_1441),
.Y(n_2428)
);

BUFx6f_ASAP7_75t_L g2429 ( 
.A(n_2084),
.Y(n_2429)
);

INVx3_ASAP7_75t_L g2430 ( 
.A(n_2054),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_2201),
.Y(n_2431)
);

INVx4_ASAP7_75t_SL g2432 ( 
.A(n_2064),
.Y(n_2432)
);

BUFx10_ASAP7_75t_L g2433 ( 
.A(n_2253),
.Y(n_2433)
);

INVx4_ASAP7_75t_L g2434 ( 
.A(n_2054),
.Y(n_2434)
);

BUFx6f_ASAP7_75t_L g2435 ( 
.A(n_2084),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2072),
.Y(n_2436)
);

AND2x4_ASAP7_75t_L g2437 ( 
.A(n_2071),
.B(n_1446),
.Y(n_2437)
);

AND2x4_ASAP7_75t_L g2438 ( 
.A(n_2105),
.B(n_1447),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2079),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_2202),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_2202),
.Y(n_2441)
);

INVx3_ASAP7_75t_L g2442 ( 
.A(n_2075),
.Y(n_2442)
);

AND2x2_ASAP7_75t_L g2443 ( 
.A(n_2223),
.B(n_1756),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2079),
.Y(n_2444)
);

AND2x2_ASAP7_75t_L g2445 ( 
.A(n_2097),
.B(n_1921),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2251),
.B(n_1449),
.Y(n_2446)
);

NOR2xp33_ASAP7_75t_L g2447 ( 
.A(n_2070),
.B(n_1732),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2245),
.B(n_1451),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2213),
.Y(n_2449)
);

CKINVDCx5p33_ASAP7_75t_R g2450 ( 
.A(n_2138),
.Y(n_2450)
);

INVx2_ASAP7_75t_L g2451 ( 
.A(n_2213),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2120),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2120),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2131),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_2218),
.Y(n_2455)
);

BUFx6f_ASAP7_75t_L g2456 ( 
.A(n_2084),
.Y(n_2456)
);

AND2x4_ASAP7_75t_L g2457 ( 
.A(n_2105),
.B(n_1456),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_2218),
.Y(n_2458)
);

BUFx3_ASAP7_75t_L g2459 ( 
.A(n_2042),
.Y(n_2459)
);

NAND2x1p5_ASAP7_75t_L g2460 ( 
.A(n_2075),
.B(n_1554),
.Y(n_2460)
);

BUFx6f_ASAP7_75t_L g2461 ( 
.A(n_2084),
.Y(n_2461)
);

XOR2x2_ASAP7_75t_L g2462 ( 
.A(n_2226),
.B(n_2044),
.Y(n_2462)
);

BUFx6f_ASAP7_75t_L g2463 ( 
.A(n_2084),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2131),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2175),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2245),
.B(n_1458),
.Y(n_2466)
);

BUFx2_ASAP7_75t_L g2467 ( 
.A(n_2042),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2097),
.B(n_1936),
.Y(n_2468)
);

INVx6_ASAP7_75t_L g2469 ( 
.A(n_2077),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2175),
.Y(n_2470)
);

CKINVDCx5p33_ASAP7_75t_R g2471 ( 
.A(n_2138),
.Y(n_2471)
);

INVx3_ASAP7_75t_L g2472 ( 
.A(n_2075),
.Y(n_2472)
);

INVx2_ASAP7_75t_SL g2473 ( 
.A(n_2063),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2144),
.Y(n_2474)
);

AND2x2_ASAP7_75t_L g2475 ( 
.A(n_2286),
.B(n_1936),
.Y(n_2475)
);

NAND2x1p5_ASAP7_75t_L g2476 ( 
.A(n_2163),
.B(n_1558),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_2021),
.B(n_1461),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_2219),
.Y(n_2478)
);

INVx2_ASAP7_75t_SL g2479 ( 
.A(n_2063),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2144),
.Y(n_2480)
);

BUFx2_ASAP7_75t_L g2481 ( 
.A(n_2117),
.Y(n_2481)
);

AND2x4_ASAP7_75t_L g2482 ( 
.A(n_2286),
.B(n_2129),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2129),
.B(n_1480),
.Y(n_2483)
);

INVx3_ASAP7_75t_L g2484 ( 
.A(n_2092),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_2219),
.Y(n_2485)
);

INVx3_ASAP7_75t_L g2486 ( 
.A(n_2092),
.Y(n_2486)
);

BUFx3_ASAP7_75t_L g2487 ( 
.A(n_2140),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2176),
.Y(n_2488)
);

NAND2x1p5_ASAP7_75t_L g2489 ( 
.A(n_2163),
.B(n_1558),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_SL g2490 ( 
.A(n_2148),
.B(n_1558),
.Y(n_2490)
);

INVx3_ASAP7_75t_L g2491 ( 
.A(n_2099),
.Y(n_2491)
);

NOR2xp33_ASAP7_75t_L g2492 ( 
.A(n_2132),
.B(n_1617),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2132),
.B(n_1484),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2145),
.Y(n_2494)
);

BUFx2_ASAP7_75t_L g2495 ( 
.A(n_2117),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2145),
.Y(n_2496)
);

INVx4_ASAP7_75t_L g2497 ( 
.A(n_2077),
.Y(n_2497)
);

HB1xp67_ASAP7_75t_L g2498 ( 
.A(n_2046),
.Y(n_2498)
);

INVx3_ASAP7_75t_L g2499 ( 
.A(n_2099),
.Y(n_2499)
);

AO22x2_ASAP7_75t_L g2500 ( 
.A1(n_2285),
.A2(n_1970),
.B1(n_1974),
.B2(n_1957),
.Y(n_2500)
);

NOR2xp33_ASAP7_75t_L g2501 ( 
.A(n_2287),
.B(n_1489),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_2176),
.Y(n_2502)
);

AND2x2_ASAP7_75t_L g2503 ( 
.A(n_2185),
.B(n_1957),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2152),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2152),
.Y(n_2505)
);

AO22x2_ASAP7_75t_L g2506 ( 
.A1(n_2285),
.A2(n_1970),
.B1(n_1974),
.B2(n_1999),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2162),
.Y(n_2507)
);

BUFx2_ASAP7_75t_L g2508 ( 
.A(n_2155),
.Y(n_2508)
);

NOR2xp33_ASAP7_75t_L g2509 ( 
.A(n_2287),
.B(n_1527),
.Y(n_2509)
);

INVx1_ASAP7_75t_SL g2510 ( 
.A(n_2155),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2205),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2162),
.Y(n_2512)
);

AND2x4_ASAP7_75t_L g2513 ( 
.A(n_2289),
.B(n_1531),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2240),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2206),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2221),
.B(n_1538),
.Y(n_2516)
);

O2A1O1Ixp5_ASAP7_75t_L g2517 ( 
.A1(n_2385),
.A2(n_2160),
.B(n_2030),
.C(n_2231),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2319),
.B(n_2033),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2320),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2321),
.Y(n_2520)
);

NOR2xp67_ASAP7_75t_L g2521 ( 
.A(n_2335),
.B(n_2358),
.Y(n_2521)
);

NAND2xp5_ASAP7_75t_SL g2522 ( 
.A(n_2319),
.B(n_2148),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2501),
.B(n_2277),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2501),
.B(n_2185),
.Y(n_2524)
);

NAND2x1p5_ASAP7_75t_L g2525 ( 
.A(n_2383),
.B(n_2013),
.Y(n_2525)
);

OR2x2_ASAP7_75t_L g2526 ( 
.A(n_2325),
.B(n_2090),
.Y(n_2526)
);

AND2x4_ASAP7_75t_L g2527 ( 
.A(n_2383),
.B(n_2159),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2509),
.B(n_2185),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_SL g2529 ( 
.A(n_2332),
.B(n_2148),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2509),
.B(n_2242),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2327),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_L g2532 ( 
.A(n_2446),
.B(n_2268),
.Y(n_2532)
);

INVxp33_ASAP7_75t_L g2533 ( 
.A(n_2331),
.Y(n_2533)
);

AOI22xp33_ASAP7_75t_L g2534 ( 
.A1(n_2445),
.A2(n_2135),
.B1(n_2259),
.B2(n_2044),
.Y(n_2534)
);

BUFx6f_ASAP7_75t_L g2535 ( 
.A(n_2395),
.Y(n_2535)
);

AOI22xp5_ASAP7_75t_L g2536 ( 
.A1(n_2349),
.A2(n_2115),
.B1(n_2284),
.B2(n_2226),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2488),
.Y(n_2537)
);

INVx2_ASAP7_75t_SL g2538 ( 
.A(n_2487),
.Y(n_2538)
);

NOR2xp33_ASAP7_75t_L g2539 ( 
.A(n_2317),
.B(n_2135),
.Y(n_2539)
);

INVx2_ASAP7_75t_L g2540 ( 
.A(n_2488),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2502),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2502),
.Y(n_2542)
);

AOI22xp33_ASAP7_75t_L g2543 ( 
.A1(n_2468),
.A2(n_2228),
.B1(n_2284),
.B2(n_2263),
.Y(n_2543)
);

OAI221xp5_ASAP7_75t_L g2544 ( 
.A1(n_2447),
.A2(n_2028),
.B1(n_2270),
.B2(n_2016),
.C(n_2027),
.Y(n_2544)
);

AND2x2_ASAP7_75t_L g2545 ( 
.A(n_2311),
.B(n_2191),
.Y(n_2545)
);

NAND2xp33_ASAP7_75t_L g2546 ( 
.A(n_2354),
.B(n_2064),
.Y(n_2546)
);

AND2x6_ASAP7_75t_SL g2547 ( 
.A(n_2314),
.B(n_2257),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2511),
.Y(n_2548)
);

AND2x2_ASAP7_75t_L g2549 ( 
.A(n_2314),
.B(n_2315),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2381),
.B(n_2272),
.Y(n_2550)
);

BUFx12f_ASAP7_75t_L g2551 ( 
.A(n_2335),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2341),
.B(n_2272),
.Y(n_2552)
);

AND2x2_ASAP7_75t_L g2553 ( 
.A(n_2315),
.B(n_2191),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_SL g2554 ( 
.A(n_2348),
.B(n_2180),
.Y(n_2554)
);

AND2x6_ASAP7_75t_SL g2555 ( 
.A(n_2343),
.B(n_2232),
.Y(n_2555)
);

BUFx3_ASAP7_75t_L g2556 ( 
.A(n_2487),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_L g2557 ( 
.A(n_2341),
.B(n_2293),
.Y(n_2557)
);

AOI22xp5_ASAP7_75t_L g2558 ( 
.A1(n_2343),
.A2(n_2246),
.B1(n_2252),
.B2(n_2273),
.Y(n_2558)
);

AOI22xp5_ASAP7_75t_L g2559 ( 
.A1(n_2447),
.A2(n_2370),
.B1(n_2339),
.B2(n_2294),
.Y(n_2559)
);

OAI22xp33_ASAP7_75t_L g2560 ( 
.A1(n_2448),
.A2(n_2263),
.B1(n_2265),
.B2(n_2262),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2338),
.Y(n_2561)
);

INVxp67_ASAP7_75t_L g2562 ( 
.A(n_2331),
.Y(n_2562)
);

BUFx6f_ASAP7_75t_L g2563 ( 
.A(n_2395),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_SL g2564 ( 
.A(n_2351),
.B(n_2180),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_SL g2565 ( 
.A(n_2513),
.B(n_2180),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_L g2566 ( 
.A(n_2299),
.B(n_2158),
.Y(n_2566)
);

INVxp67_ASAP7_75t_SL g2567 ( 
.A(n_2498),
.Y(n_2567)
);

A2O1A1Ixp33_ASAP7_75t_L g2568 ( 
.A1(n_2339),
.A2(n_2266),
.B(n_2271),
.C(n_2209),
.Y(n_2568)
);

NAND2xp33_ASAP7_75t_L g2569 ( 
.A(n_2484),
.B(n_2064),
.Y(n_2569)
);

AOI22xp33_ASAP7_75t_L g2570 ( 
.A1(n_2500),
.A2(n_2263),
.B1(n_2262),
.B2(n_2260),
.Y(n_2570)
);

NAND2xp33_ASAP7_75t_L g2571 ( 
.A(n_2484),
.B(n_2064),
.Y(n_2571)
);

NOR2xp33_ASAP7_75t_L g2572 ( 
.A(n_2295),
.B(n_2306),
.Y(n_2572)
);

INVx2_ASAP7_75t_SL g2573 ( 
.A(n_2328),
.Y(n_2573)
);

AND2x2_ASAP7_75t_L g2574 ( 
.A(n_2347),
.B(n_2159),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2345),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_2511),
.Y(n_2576)
);

NOR2xp33_ASAP7_75t_L g2577 ( 
.A(n_2306),
.B(n_2273),
.Y(n_2577)
);

BUFx10_ASAP7_75t_L g2578 ( 
.A(n_2363),
.Y(n_2578)
);

A2O1A1Ixp33_ASAP7_75t_L g2579 ( 
.A1(n_2305),
.A2(n_2266),
.B(n_2211),
.C(n_2254),
.Y(n_2579)
);

NAND2xp33_ASAP7_75t_L g2580 ( 
.A(n_2486),
.B(n_2064),
.Y(n_2580)
);

INVx2_ASAP7_75t_L g2581 ( 
.A(n_2290),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2355),
.Y(n_2582)
);

BUFx5_ASAP7_75t_L g2583 ( 
.A(n_2388),
.Y(n_2583)
);

AOI21xp5_ASAP7_75t_L g2584 ( 
.A1(n_2291),
.A2(n_2106),
.B(n_2035),
.Y(n_2584)
);

NAND2xp33_ASAP7_75t_L g2585 ( 
.A(n_2486),
.B(n_2064),
.Y(n_2585)
);

AND2x2_ASAP7_75t_L g2586 ( 
.A(n_2475),
.B(n_2158),
.Y(n_2586)
);

NOR2xp33_ASAP7_75t_L g2587 ( 
.A(n_2295),
.B(n_2116),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_L g2588 ( 
.A(n_2302),
.B(n_2215),
.Y(n_2588)
);

INVx2_ASAP7_75t_L g2589 ( 
.A(n_2290),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_L g2590 ( 
.A(n_2304),
.B(n_2220),
.Y(n_2590)
);

OR2x6_ASAP7_75t_SL g2591 ( 
.A(n_2363),
.B(n_1959),
.Y(n_2591)
);

AND2x2_ASAP7_75t_L g2592 ( 
.A(n_2503),
.B(n_2116),
.Y(n_2592)
);

AND2x6_ASAP7_75t_SL g2593 ( 
.A(n_2362),
.B(n_2265),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_L g2594 ( 
.A(n_2307),
.B(n_2267),
.Y(n_2594)
);

OAI22xp33_ASAP7_75t_L g2595 ( 
.A1(n_2466),
.A2(n_2265),
.B1(n_2280),
.B2(n_1977),
.Y(n_2595)
);

AOI22xp33_ASAP7_75t_L g2596 ( 
.A1(n_2500),
.A2(n_2187),
.B1(n_2250),
.B2(n_2247),
.Y(n_2596)
);

HB1xp67_ASAP7_75t_L g2597 ( 
.A(n_2498),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2364),
.Y(n_2598)
);

NOR2xp67_ASAP7_75t_L g2599 ( 
.A(n_2398),
.B(n_2013),
.Y(n_2599)
);

AND2x2_ASAP7_75t_L g2600 ( 
.A(n_2308),
.B(n_2265),
.Y(n_2600)
);

OAI22xp5_ASAP7_75t_L g2601 ( 
.A1(n_2291),
.A2(n_2235),
.B1(n_2280),
.B2(n_2198),
.Y(n_2601)
);

OAI22xp5_ASAP7_75t_L g2602 ( 
.A1(n_2334),
.A2(n_2198),
.B1(n_2154),
.B2(n_2066),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_2292),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2292),
.Y(n_2604)
);

OR2x6_ASAP7_75t_L g2605 ( 
.A(n_2411),
.B(n_2222),
.Y(n_2605)
);

INVxp67_ASAP7_75t_L g2606 ( 
.A(n_2409),
.Y(n_2606)
);

AOI22xp33_ASAP7_75t_L g2607 ( 
.A1(n_2500),
.A2(n_2166),
.B1(n_2193),
.B2(n_2222),
.Y(n_2607)
);

NOR2xp33_ASAP7_75t_L g2608 ( 
.A(n_2309),
.B(n_2095),
.Y(n_2608)
);

NOR2xp33_ASAP7_75t_L g2609 ( 
.A(n_2309),
.B(n_2221),
.Y(n_2609)
);

INVxp67_ASAP7_75t_L g2610 ( 
.A(n_2409),
.Y(n_2610)
);

BUFx3_ASAP7_75t_L g2611 ( 
.A(n_2508),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2318),
.B(n_2121),
.Y(n_2612)
);

INVx2_ASAP7_75t_SL g2613 ( 
.A(n_2395),
.Y(n_2613)
);

OR2x6_ASAP7_75t_L g2614 ( 
.A(n_2411),
.B(n_2006),
.Y(n_2614)
);

NOR2xp33_ASAP7_75t_L g2615 ( 
.A(n_2357),
.B(n_2067),
.Y(n_2615)
);

NOR2xp33_ASAP7_75t_L g2616 ( 
.A(n_2481),
.B(n_1906),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_SL g2617 ( 
.A(n_2495),
.B(n_2099),
.Y(n_2617)
);

AOI22xp33_ASAP7_75t_L g2618 ( 
.A1(n_2397),
.A2(n_2094),
.B1(n_1964),
.B2(n_1992),
.Y(n_2618)
);

AND2x4_ASAP7_75t_L g2619 ( 
.A(n_2432),
.B(n_2006),
.Y(n_2619)
);

AND2x4_ASAP7_75t_L g2620 ( 
.A(n_2432),
.B(n_2009),
.Y(n_2620)
);

INVx2_ASAP7_75t_L g2621 ( 
.A(n_2296),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_SL g2622 ( 
.A(n_2310),
.B(n_2157),
.Y(n_2622)
);

AND2x2_ASAP7_75t_L g2623 ( 
.A(n_2482),
.B(n_2009),
.Y(n_2623)
);

AOI22xp33_ASAP7_75t_L g2624 ( 
.A1(n_2397),
.A2(n_2094),
.B1(n_1979),
.B2(n_2001),
.Y(n_2624)
);

A2O1A1Ixp33_ASAP7_75t_L g2625 ( 
.A1(n_2492),
.A2(n_2362),
.B(n_2301),
.C(n_2369),
.Y(n_2625)
);

AND2x2_ASAP7_75t_L g2626 ( 
.A(n_2482),
.B(n_1546),
.Y(n_2626)
);

NOR3xp33_ASAP7_75t_L g2627 ( 
.A(n_2301),
.B(n_2003),
.C(n_1996),
.Y(n_2627)
);

AOI22xp5_ASAP7_75t_L g2628 ( 
.A1(n_2506),
.A2(n_2094),
.B1(n_2121),
.B2(n_2269),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_L g2629 ( 
.A(n_2398),
.B(n_2121),
.Y(n_2629)
);

OAI22xp5_ASAP7_75t_L g2630 ( 
.A1(n_2483),
.A2(n_2154),
.B1(n_2198),
.B2(n_2217),
.Y(n_2630)
);

INVx2_ASAP7_75t_L g2631 ( 
.A(n_2296),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_L g2632 ( 
.A(n_2413),
.B(n_2121),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_2516),
.B(n_2121),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_2392),
.B(n_2121),
.Y(n_2634)
);

INVx4_ASAP7_75t_L g2635 ( 
.A(n_2469),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_2303),
.Y(n_2636)
);

INVxp67_ASAP7_75t_L g2637 ( 
.A(n_2310),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2303),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_SL g2639 ( 
.A(n_2324),
.B(n_2157),
.Y(n_2639)
);

NOR2xp33_ASAP7_75t_L g2640 ( 
.A(n_2316),
.B(n_1834),
.Y(n_2640)
);

INVx2_ASAP7_75t_SL g2641 ( 
.A(n_2346),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_L g2642 ( 
.A(n_2392),
.B(n_2094),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_L g2643 ( 
.A(n_2333),
.B(n_2094),
.Y(n_2643)
);

NAND2x1p5_ASAP7_75t_L g2644 ( 
.A(n_2497),
.B(n_2013),
.Y(n_2644)
);

NAND2x1p5_ASAP7_75t_L g2645 ( 
.A(n_2497),
.B(n_2026),
.Y(n_2645)
);

INVx2_ASAP7_75t_L g2646 ( 
.A(n_2312),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2365),
.Y(n_2647)
);

AND2x2_ASAP7_75t_L g2648 ( 
.A(n_2394),
.B(n_1548),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2367),
.Y(n_2649)
);

AOI21xp5_ASAP7_75t_L g2650 ( 
.A1(n_2426),
.A2(n_2106),
.B(n_2040),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_L g2651 ( 
.A(n_2333),
.B(n_2368),
.Y(n_2651)
);

NOR2x1p5_ASAP7_75t_L g2652 ( 
.A(n_2346),
.B(n_2412),
.Y(n_2652)
);

BUFx12f_ASAP7_75t_L g2653 ( 
.A(n_2412),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_2368),
.B(n_2094),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2373),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2514),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2312),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2324),
.B(n_2096),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_SL g2659 ( 
.A(n_2433),
.B(n_2157),
.Y(n_2659)
);

AOI22xp5_ASAP7_75t_L g2660 ( 
.A1(n_2506),
.A2(n_2275),
.B1(n_2029),
.B2(n_2244),
.Y(n_2660)
);

AO221x1_ASAP7_75t_L g2661 ( 
.A1(n_2506),
.A2(n_1910),
.B1(n_1900),
.B2(n_2039),
.C(n_2026),
.Y(n_2661)
);

OR2x2_ASAP7_75t_L g2662 ( 
.A(n_2467),
.B(n_1506),
.Y(n_2662)
);

AND2x2_ASAP7_75t_SL g2663 ( 
.A(n_2432),
.B(n_2282),
.Y(n_2663)
);

NOR2xp33_ASAP7_75t_L g2664 ( 
.A(n_2450),
.B(n_1887),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2374),
.Y(n_2665)
);

AOI22xp33_ASAP7_75t_L g2666 ( 
.A1(n_2397),
.A2(n_2256),
.B1(n_2244),
.B2(n_1918),
.Y(n_2666)
);

AOI22x1_ASAP7_75t_SL g2667 ( 
.A1(n_2450),
.A2(n_2471),
.B1(n_2389),
.B2(n_2510),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_2378),
.B(n_1555),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_L g2669 ( 
.A(n_2382),
.B(n_1567),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2386),
.B(n_1569),
.Y(n_2670)
);

INVxp67_ASAP7_75t_L g2671 ( 
.A(n_2410),
.Y(n_2671)
);

NOR2xp33_ASAP7_75t_L g2672 ( 
.A(n_2471),
.B(n_2077),
.Y(n_2672)
);

AND2x6_ASAP7_75t_L g2673 ( 
.A(n_2429),
.B(n_2258),
.Y(n_2673)
);

AOI22xp5_ASAP7_75t_L g2674 ( 
.A1(n_2388),
.A2(n_2244),
.B1(n_2177),
.B2(n_2032),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_2391),
.B(n_1570),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_SL g2676 ( 
.A(n_2433),
.B(n_2087),
.Y(n_2676)
);

A2O1A1Ixp33_ASAP7_75t_L g2677 ( 
.A1(n_2492),
.A2(n_2200),
.B(n_2051),
.C(n_2208),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2393),
.B(n_1506),
.Y(n_2678)
);

AOI22xp5_ASAP7_75t_L g2679 ( 
.A1(n_2388),
.A2(n_2244),
.B1(n_1943),
.B2(n_2142),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_L g2680 ( 
.A(n_2396),
.B(n_1509),
.Y(n_2680)
);

AND2x2_ASAP7_75t_L g2681 ( 
.A(n_2437),
.B(n_1509),
.Y(n_2681)
);

NOR2x1p5_ASAP7_75t_L g2682 ( 
.A(n_2416),
.B(n_2195),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2313),
.Y(n_2683)
);

NOR2xp33_ASAP7_75t_L g2684 ( 
.A(n_2404),
.B(n_2477),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2418),
.B(n_1518),
.Y(n_2685)
);

INVx2_ASAP7_75t_L g2686 ( 
.A(n_2313),
.Y(n_2686)
);

INVx2_ASAP7_75t_L g2687 ( 
.A(n_2322),
.Y(n_2687)
);

NOR2xp33_ASAP7_75t_L g2688 ( 
.A(n_2406),
.B(n_2417),
.Y(n_2688)
);

AOI22xp33_ASAP7_75t_L g2689 ( 
.A1(n_2297),
.A2(n_2244),
.B1(n_1533),
.B2(n_1534),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_2419),
.B(n_1530),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2436),
.B(n_1530),
.Y(n_2691)
);

AOI22xp33_ASAP7_75t_L g2692 ( 
.A1(n_2297),
.A2(n_2244),
.B1(n_1534),
.B2(n_1539),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2439),
.B(n_1533),
.Y(n_2693)
);

INVx2_ASAP7_75t_L g2694 ( 
.A(n_2322),
.Y(n_2694)
);

AOI22xp5_ASAP7_75t_L g2695 ( 
.A1(n_2388),
.A2(n_2114),
.B1(n_2198),
.B2(n_2154),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2444),
.B(n_1539),
.Y(n_2696)
);

INVx5_ASAP7_75t_L g2697 ( 
.A(n_2388),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2452),
.Y(n_2698)
);

INVx4_ASAP7_75t_L g2699 ( 
.A(n_2697),
.Y(n_2699)
);

INVx2_ASAP7_75t_L g2700 ( 
.A(n_2581),
.Y(n_2700)
);

BUFx3_ASAP7_75t_L g2701 ( 
.A(n_2551),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_SL g2702 ( 
.A(n_2601),
.B(n_2404),
.Y(n_2702)
);

INVx4_ASAP7_75t_L g2703 ( 
.A(n_2527),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2519),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2520),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_2518),
.B(n_2424),
.Y(n_2706)
);

INVx1_ASAP7_75t_SL g2707 ( 
.A(n_2556),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2523),
.B(n_2524),
.Y(n_2708)
);

NOR2xp33_ASAP7_75t_L g2709 ( 
.A(n_2530),
.B(n_2469),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2531),
.Y(n_2710)
);

OR2x2_ASAP7_75t_L g2711 ( 
.A(n_2549),
.B(n_2353),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2589),
.Y(n_2712)
);

INVx2_ASAP7_75t_L g2713 ( 
.A(n_2603),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2604),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2621),
.Y(n_2715)
);

INVx3_ASAP7_75t_L g2716 ( 
.A(n_2697),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2631),
.Y(n_2717)
);

HB1xp67_ASAP7_75t_L g2718 ( 
.A(n_2597),
.Y(n_2718)
);

AND3x1_ASAP7_75t_SL g2719 ( 
.A(n_2652),
.B(n_2454),
.C(n_2453),
.Y(n_2719)
);

OR2x2_ASAP7_75t_L g2720 ( 
.A(n_2550),
.B(n_2297),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_L g2721 ( 
.A(n_2528),
.B(n_2424),
.Y(n_2721)
);

OR2x2_ASAP7_75t_L g2722 ( 
.A(n_2562),
.B(n_2597),
.Y(n_2722)
);

NAND2xp33_ASAP7_75t_SL g2723 ( 
.A(n_2618),
.B(n_2093),
.Y(n_2723)
);

NOR2xp33_ASAP7_75t_L g2724 ( 
.A(n_2559),
.B(n_2469),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2636),
.Y(n_2725)
);

AND2x2_ASAP7_75t_L g2726 ( 
.A(n_2586),
.B(n_2416),
.Y(n_2726)
);

AND2x4_ASAP7_75t_L g2727 ( 
.A(n_2697),
.B(n_2429),
.Y(n_2727)
);

NOR2xp33_ASAP7_75t_L g2728 ( 
.A(n_2544),
.B(n_2406),
.Y(n_2728)
);

INVxp67_ASAP7_75t_L g2729 ( 
.A(n_2566),
.Y(n_2729)
);

BUFx4f_ASAP7_75t_L g2730 ( 
.A(n_2653),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_L g2731 ( 
.A(n_2625),
.B(n_2464),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2561),
.Y(n_2732)
);

INVx2_ASAP7_75t_L g2733 ( 
.A(n_2638),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2646),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_2609),
.B(n_2465),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2609),
.B(n_2470),
.Y(n_2736)
);

BUFx6f_ASAP7_75t_L g2737 ( 
.A(n_2697),
.Y(n_2737)
);

INVx3_ASAP7_75t_L g2738 ( 
.A(n_2635),
.Y(n_2738)
);

NOR2xp33_ASAP7_75t_L g2739 ( 
.A(n_2544),
.B(n_2417),
.Y(n_2739)
);

INVx2_ASAP7_75t_L g2740 ( 
.A(n_2657),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2615),
.B(n_2437),
.Y(n_2741)
);

BUFx3_ASAP7_75t_L g2742 ( 
.A(n_2527),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2575),
.Y(n_2743)
);

INVx5_ASAP7_75t_L g2744 ( 
.A(n_2673),
.Y(n_2744)
);

INVx1_ASAP7_75t_SL g2745 ( 
.A(n_2611),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2615),
.B(n_2438),
.Y(n_2746)
);

INVx6_ASAP7_75t_L g2747 ( 
.A(n_2635),
.Y(n_2747)
);

INVx1_ASAP7_75t_SL g2748 ( 
.A(n_2578),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_SL g2749 ( 
.A(n_2595),
.B(n_2422),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2683),
.Y(n_2750)
);

INVx3_ASAP7_75t_L g2751 ( 
.A(n_2535),
.Y(n_2751)
);

INVx3_ASAP7_75t_L g2752 ( 
.A(n_2535),
.Y(n_2752)
);

INVx2_ASAP7_75t_SL g2753 ( 
.A(n_2682),
.Y(n_2753)
);

INVx2_ASAP7_75t_L g2754 ( 
.A(n_2686),
.Y(n_2754)
);

HB1xp67_ASAP7_75t_L g2755 ( 
.A(n_2567),
.Y(n_2755)
);

INVx3_ASAP7_75t_L g2756 ( 
.A(n_2535),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2582),
.Y(n_2757)
);

OR2x2_ASAP7_75t_L g2758 ( 
.A(n_2562),
.B(n_2459),
.Y(n_2758)
);

BUFx3_ASAP7_75t_L g2759 ( 
.A(n_2563),
.Y(n_2759)
);

HB1xp67_ASAP7_75t_L g2760 ( 
.A(n_2567),
.Y(n_2760)
);

INVxp67_ASAP7_75t_L g2761 ( 
.A(n_2577),
.Y(n_2761)
);

AND3x2_ASAP7_75t_SL g2762 ( 
.A(n_2593),
.B(n_2261),
.C(n_2258),
.Y(n_2762)
);

BUFx2_ASAP7_75t_L g2763 ( 
.A(n_2637),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_2671),
.B(n_2438),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2598),
.Y(n_2765)
);

A2O1A1Ixp33_ASAP7_75t_SL g2766 ( 
.A1(n_2664),
.A2(n_2491),
.B(n_2499),
.C(n_2248),
.Y(n_2766)
);

INVx3_ASAP7_75t_L g2767 ( 
.A(n_2563),
.Y(n_2767)
);

AND2x6_ASAP7_75t_L g2768 ( 
.A(n_2628),
.B(n_2261),
.Y(n_2768)
);

AOI22xp33_ASAP7_75t_SL g2769 ( 
.A1(n_2539),
.A2(n_2443),
.B1(n_2389),
.B2(n_2402),
.Y(n_2769)
);

INVx2_ASAP7_75t_L g2770 ( 
.A(n_2687),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2647),
.Y(n_2771)
);

NOR2xp33_ASAP7_75t_L g2772 ( 
.A(n_2539),
.B(n_2421),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2649),
.Y(n_2773)
);

INVx2_ASAP7_75t_L g2774 ( 
.A(n_2694),
.Y(n_2774)
);

BUFx6f_ASAP7_75t_L g2775 ( 
.A(n_2619),
.Y(n_2775)
);

OR2x4_ASAP7_75t_L g2776 ( 
.A(n_2640),
.B(n_2429),
.Y(n_2776)
);

BUFx8_ASAP7_75t_L g2777 ( 
.A(n_2574),
.Y(n_2777)
);

AND2x4_ASAP7_75t_L g2778 ( 
.A(n_2619),
.B(n_2429),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2655),
.Y(n_2779)
);

NOR2xp33_ASAP7_75t_L g2780 ( 
.A(n_2522),
.B(n_2421),
.Y(n_2780)
);

INVx2_ASAP7_75t_SL g2781 ( 
.A(n_2578),
.Y(n_2781)
);

BUFx6f_ASAP7_75t_L g2782 ( 
.A(n_2620),
.Y(n_2782)
);

BUFx2_ASAP7_75t_L g2783 ( 
.A(n_2637),
.Y(n_2783)
);

INVx3_ASAP7_75t_L g2784 ( 
.A(n_2563),
.Y(n_2784)
);

INVx2_ASAP7_75t_L g2785 ( 
.A(n_2537),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_SL g2786 ( 
.A(n_2595),
.B(n_2490),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2540),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2665),
.Y(n_2788)
);

INVx4_ASAP7_75t_L g2789 ( 
.A(n_2614),
.Y(n_2789)
);

AOI22xp5_ASAP7_75t_L g2790 ( 
.A1(n_2536),
.A2(n_2402),
.B1(n_2457),
.B2(n_2428),
.Y(n_2790)
);

INVx4_ASAP7_75t_L g2791 ( 
.A(n_2614),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2541),
.Y(n_2792)
);

INVx3_ASAP7_75t_L g2793 ( 
.A(n_2525),
.Y(n_2793)
);

INVx2_ASAP7_75t_L g2794 ( 
.A(n_2542),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_SL g2795 ( 
.A(n_2568),
.B(n_2490),
.Y(n_2795)
);

BUFx3_ASAP7_75t_L g2796 ( 
.A(n_2688),
.Y(n_2796)
);

BUFx2_ASAP7_75t_L g2797 ( 
.A(n_2592),
.Y(n_2797)
);

INVx2_ASAP7_75t_L g2798 ( 
.A(n_2548),
.Y(n_2798)
);

AOI22xp5_ASAP7_75t_L g2799 ( 
.A1(n_2534),
.A2(n_2402),
.B1(n_2428),
.B2(n_2384),
.Y(n_2799)
);

INVx2_ASAP7_75t_SL g2800 ( 
.A(n_2538),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2698),
.Y(n_2801)
);

NOR2xp33_ASAP7_75t_L g2802 ( 
.A(n_2608),
.B(n_2421),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2532),
.B(n_2515),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2656),
.Y(n_2804)
);

AND2x4_ASAP7_75t_L g2805 ( 
.A(n_2620),
.B(n_2435),
.Y(n_2805)
);

INVx2_ASAP7_75t_SL g2806 ( 
.A(n_2613),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_2576),
.Y(n_2807)
);

INVx2_ASAP7_75t_SL g2808 ( 
.A(n_2573),
.Y(n_2808)
);

INVx5_ASAP7_75t_L g2809 ( 
.A(n_2673),
.Y(n_2809)
);

AND2x4_ASAP7_75t_L g2810 ( 
.A(n_2605),
.B(n_2435),
.Y(n_2810)
);

BUFx2_ASAP7_75t_L g2811 ( 
.A(n_2641),
.Y(n_2811)
);

BUFx6f_ASAP7_75t_L g2812 ( 
.A(n_2605),
.Y(n_2812)
);

AND2x2_ASAP7_75t_L g2813 ( 
.A(n_2534),
.B(n_2459),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2594),
.Y(n_2814)
);

BUFx6f_ASAP7_75t_L g2815 ( 
.A(n_2605),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2552),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2557),
.Y(n_2817)
);

NOR2xp33_ASAP7_75t_R g2818 ( 
.A(n_2569),
.B(n_2298),
.Y(n_2818)
);

INVx2_ASAP7_75t_SL g2819 ( 
.A(n_2648),
.Y(n_2819)
);

INVx3_ASAP7_75t_L g2820 ( 
.A(n_2525),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2606),
.Y(n_2821)
);

CKINVDCx20_ASAP7_75t_R g2822 ( 
.A(n_2667),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2606),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2610),
.Y(n_2824)
);

NOR2xp33_ASAP7_75t_R g2825 ( 
.A(n_2571),
.B(n_2330),
.Y(n_2825)
);

NOR2xp33_ASAP7_75t_L g2826 ( 
.A(n_2608),
.B(n_2493),
.Y(n_2826)
);

INVx3_ASAP7_75t_L g2827 ( 
.A(n_2644),
.Y(n_2827)
);

BUFx3_ASAP7_75t_L g2828 ( 
.A(n_2587),
.Y(n_2828)
);

INVx3_ASAP7_75t_L g2829 ( 
.A(n_2644),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_SL g2830 ( 
.A(n_2602),
.B(n_2426),
.Y(n_2830)
);

HB1xp67_ASAP7_75t_L g2831 ( 
.A(n_2610),
.Y(n_2831)
);

BUFx6f_ASAP7_75t_L g2832 ( 
.A(n_2673),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2588),
.Y(n_2833)
);

INVx3_ASAP7_75t_L g2834 ( 
.A(n_2645),
.Y(n_2834)
);

INVx3_ASAP7_75t_L g2835 ( 
.A(n_2645),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2632),
.Y(n_2836)
);

INVx5_ASAP7_75t_L g2837 ( 
.A(n_2673),
.Y(n_2837)
);

INVx2_ASAP7_75t_L g2838 ( 
.A(n_2673),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2590),
.Y(n_2839)
);

AND2x2_ASAP7_75t_L g2840 ( 
.A(n_2572),
.B(n_2473),
.Y(n_2840)
);

INVx3_ASAP7_75t_L g2841 ( 
.A(n_2614),
.Y(n_2841)
);

INVx4_ASAP7_75t_L g2842 ( 
.A(n_2626),
.Y(n_2842)
);

CKINVDCx5p33_ASAP7_75t_R g2843 ( 
.A(n_2547),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_L g2844 ( 
.A(n_2572),
.B(n_2479),
.Y(n_2844)
);

INVx2_ASAP7_75t_L g2845 ( 
.A(n_2612),
.Y(n_2845)
);

BUFx3_ASAP7_75t_L g2846 ( 
.A(n_2672),
.Y(n_2846)
);

INVx2_ASAP7_75t_SL g2847 ( 
.A(n_2662),
.Y(n_2847)
);

INVxp67_ASAP7_75t_SL g2848 ( 
.A(n_2580),
.Y(n_2848)
);

OR2x6_ASAP7_75t_L g2849 ( 
.A(n_2643),
.B(n_2274),
.Y(n_2849)
);

HB1xp67_ASAP7_75t_L g2850 ( 
.A(n_2553),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2678),
.Y(n_2851)
);

BUFx4f_ASAP7_75t_L g2852 ( 
.A(n_2526),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_2651),
.B(n_2323),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2680),
.Y(n_2854)
);

INVx1_ASAP7_75t_SL g2855 ( 
.A(n_2533),
.Y(n_2855)
);

AOI22xp33_ASAP7_75t_L g2856 ( 
.A1(n_2627),
.A2(n_2462),
.B1(n_2384),
.B2(n_2377),
.Y(n_2856)
);

INVx2_ASAP7_75t_SL g2857 ( 
.A(n_2623),
.Y(n_2857)
);

INVx1_ASAP7_75t_SL g2858 ( 
.A(n_2565),
.Y(n_2858)
);

AND2x4_ASAP7_75t_SL g2859 ( 
.A(n_2681),
.B(n_2435),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2685),
.Y(n_2860)
);

AOI22xp33_ASAP7_75t_L g2861 ( 
.A1(n_2543),
.A2(n_2384),
.B1(n_2377),
.B2(n_2402),
.Y(n_2861)
);

BUFx6f_ASAP7_75t_L g2862 ( 
.A(n_2663),
.Y(n_2862)
);

CKINVDCx5p33_ASAP7_75t_R g2863 ( 
.A(n_2555),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2690),
.Y(n_2864)
);

CKINVDCx8_ASAP7_75t_R g2865 ( 
.A(n_2616),
.Y(n_2865)
);

CKINVDCx16_ASAP7_75t_R g2866 ( 
.A(n_2591),
.Y(n_2866)
);

INVxp67_ASAP7_75t_L g2867 ( 
.A(n_2545),
.Y(n_2867)
);

INVx5_ASAP7_75t_L g2868 ( 
.A(n_2600),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2691),
.Y(n_2869)
);

BUFx3_ASAP7_75t_L g2870 ( 
.A(n_2629),
.Y(n_2870)
);

AND2x2_ASAP7_75t_L g2871 ( 
.A(n_2558),
.B(n_2344),
.Y(n_2871)
);

INVx2_ASAP7_75t_L g2872 ( 
.A(n_2693),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2554),
.B(n_2323),
.Y(n_2873)
);

BUFx2_ASAP7_75t_L g2874 ( 
.A(n_2634),
.Y(n_2874)
);

INVx2_ASAP7_75t_L g2875 ( 
.A(n_2696),
.Y(n_2875)
);

INVx3_ASAP7_75t_L g2876 ( 
.A(n_2583),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_2579),
.B(n_2529),
.Y(n_2877)
);

INVx2_ASAP7_75t_L g2878 ( 
.A(n_2633),
.Y(n_2878)
);

AND2x2_ASAP7_75t_L g2879 ( 
.A(n_2543),
.B(n_2326),
.Y(n_2879)
);

A2O1A1Ixp33_ASAP7_75t_L g2880 ( 
.A1(n_2728),
.A2(n_2517),
.B(n_2624),
.C(n_2618),
.Y(n_2880)
);

HB1xp67_ASAP7_75t_L g2881 ( 
.A(n_2718),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_SL g2882 ( 
.A(n_2852),
.B(n_2583),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2708),
.B(n_2684),
.Y(n_2883)
);

CKINVDCx8_ASAP7_75t_R g2884 ( 
.A(n_2863),
.Y(n_2884)
);

AOI21x1_ASAP7_75t_L g2885 ( 
.A1(n_2795),
.A2(n_2564),
.B(n_2676),
.Y(n_2885)
);

INVx2_ASAP7_75t_L g2886 ( 
.A(n_2785),
.Y(n_2886)
);

AOI21xp5_ASAP7_75t_L g2887 ( 
.A1(n_2848),
.A2(n_2585),
.B(n_2584),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2826),
.B(n_2684),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_L g2889 ( 
.A(n_2826),
.B(n_2666),
.Y(n_2889)
);

AOI22x1_ASAP7_75t_L g2890 ( 
.A1(n_2748),
.A2(n_2434),
.B1(n_2499),
.B2(n_2491),
.Y(n_2890)
);

AOI21xp5_ASAP7_75t_L g2891 ( 
.A1(n_2848),
.A2(n_2584),
.B(n_2546),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_SL g2892 ( 
.A(n_2852),
.B(n_2583),
.Y(n_2892)
);

AOI22xp33_ASAP7_75t_L g2893 ( 
.A1(n_2862),
.A2(n_2689),
.B1(n_2692),
.B2(n_2624),
.Y(n_2893)
);

BUFx12f_ASAP7_75t_L g2894 ( 
.A(n_2843),
.Y(n_2894)
);

AOI21xp5_ASAP7_75t_L g2895 ( 
.A1(n_2749),
.A2(n_2650),
.B(n_2677),
.Y(n_2895)
);

AND2x2_ASAP7_75t_L g2896 ( 
.A(n_2797),
.B(n_2666),
.Y(n_2896)
);

A2O1A1Ixp33_ASAP7_75t_L g2897 ( 
.A1(n_2728),
.A2(n_2517),
.B(n_2660),
.C(n_2679),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2831),
.Y(n_2898)
);

OAI22xp5_ASAP7_75t_L g2899 ( 
.A1(n_2856),
.A2(n_2692),
.B1(n_2689),
.B2(n_2674),
.Y(n_2899)
);

AOI22xp33_ASAP7_75t_L g2900 ( 
.A1(n_2862),
.A2(n_2661),
.B1(n_2663),
.B2(n_2560),
.Y(n_2900)
);

NOR2xp33_ASAP7_75t_L g2901 ( 
.A(n_2846),
.B(n_2659),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2831),
.Y(n_2902)
);

CKINVDCx11_ASAP7_75t_R g2903 ( 
.A(n_2822),
.Y(n_2903)
);

INVx3_ASAP7_75t_L g2904 ( 
.A(n_2789),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_SL g2905 ( 
.A(n_2818),
.B(n_2583),
.Y(n_2905)
);

NOR2xp33_ASAP7_75t_L g2906 ( 
.A(n_2846),
.B(n_2521),
.Y(n_2906)
);

AOI21xp5_ASAP7_75t_L g2907 ( 
.A1(n_2749),
.A2(n_2650),
.B(n_2100),
.Y(n_2907)
);

INVx2_ASAP7_75t_L g2908 ( 
.A(n_2787),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2718),
.Y(n_2909)
);

A2O1A1Ixp33_ASAP7_75t_L g2910 ( 
.A1(n_2739),
.A2(n_2695),
.B(n_2599),
.C(n_2630),
.Y(n_2910)
);

CKINVDCx16_ASAP7_75t_R g2911 ( 
.A(n_2822),
.Y(n_2911)
);

CKINVDCx20_ASAP7_75t_R g2912 ( 
.A(n_2701),
.Y(n_2912)
);

AOI21xp5_ASAP7_75t_L g2913 ( 
.A1(n_2795),
.A2(n_2560),
.B(n_2237),
.Y(n_2913)
);

OAI22xp5_ASAP7_75t_L g2914 ( 
.A1(n_2856),
.A2(n_2607),
.B1(n_2570),
.B2(n_2654),
.Y(n_2914)
);

AO32x1_ASAP7_75t_L g2915 ( 
.A1(n_2847),
.A2(n_2274),
.A3(n_2224),
.B1(n_2237),
.B2(n_2326),
.Y(n_2915)
);

A2O1A1Ixp33_ASAP7_75t_L g2916 ( 
.A1(n_2739),
.A2(n_2607),
.B(n_2596),
.C(n_2658),
.Y(n_2916)
);

AOI21xp5_ASAP7_75t_L g2917 ( 
.A1(n_2723),
.A2(n_2224),
.B(n_2248),
.Y(n_2917)
);

HB1xp67_ASAP7_75t_L g2918 ( 
.A(n_2755),
.Y(n_2918)
);

AND2x2_ASAP7_75t_SL g2919 ( 
.A(n_2862),
.B(n_2570),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_L g2920 ( 
.A(n_2817),
.B(n_2642),
.Y(n_2920)
);

OAI22xp5_ASAP7_75t_L g2921 ( 
.A1(n_2861),
.A2(n_2596),
.B1(n_2669),
.B2(n_2668),
.Y(n_2921)
);

O2A1O1Ixp33_ASAP7_75t_L g2922 ( 
.A1(n_2877),
.A2(n_2622),
.B(n_2639),
.C(n_2617),
.Y(n_2922)
);

OAI22xp5_ASAP7_75t_L g2923 ( 
.A1(n_2861),
.A2(n_2670),
.B1(n_2675),
.B2(n_2154),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2788),
.Y(n_2924)
);

AOI21xp33_ASAP7_75t_L g2925 ( 
.A1(n_2786),
.A2(n_2830),
.B(n_2799),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_2735),
.B(n_2329),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2736),
.B(n_2329),
.Y(n_2927)
);

OAI22xp5_ASAP7_75t_L g2928 ( 
.A1(n_2866),
.A2(n_2214),
.B1(n_2216),
.B2(n_2205),
.Y(n_2928)
);

OAI21xp5_ASAP7_75t_L g2929 ( 
.A1(n_2786),
.A2(n_2170),
.B(n_2109),
.Y(n_2929)
);

INVxp67_ASAP7_75t_L g2930 ( 
.A(n_2840),
.Y(n_2930)
);

A2O1A1Ixp33_ASAP7_75t_L g2931 ( 
.A1(n_2723),
.A2(n_2195),
.B(n_1847),
.C(n_1846),
.Y(n_2931)
);

OAI21xp33_ASAP7_75t_L g2932 ( 
.A1(n_2731),
.A2(n_1550),
.B(n_1540),
.Y(n_2932)
);

O2A1O1Ixp33_ASAP7_75t_L g2933 ( 
.A1(n_2729),
.A2(n_1550),
.B(n_1552),
.C(n_1540),
.Y(n_2933)
);

OAI22xp5_ASAP7_75t_L g2934 ( 
.A1(n_2790),
.A2(n_2216),
.B1(n_2214),
.B2(n_2342),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2833),
.B(n_2839),
.Y(n_2935)
);

AND2x2_ASAP7_75t_L g2936 ( 
.A(n_2726),
.B(n_2435),
.Y(n_2936)
);

AOI21xp5_ASAP7_75t_L g2937 ( 
.A1(n_2830),
.A2(n_2236),
.B(n_2147),
.Y(n_2937)
);

OR2x2_ASAP7_75t_L g2938 ( 
.A(n_2722),
.B(n_2711),
.Y(n_2938)
);

OAI22xp5_ASAP7_75t_L g2939 ( 
.A1(n_2865),
.A2(n_2350),
.B1(n_2352),
.B2(n_2336),
.Y(n_2939)
);

O2A1O1Ixp33_ASAP7_75t_L g2940 ( 
.A1(n_2766),
.A2(n_1564),
.B(n_1556),
.C(n_1520),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_SL g2941 ( 
.A(n_2818),
.B(n_2583),
.Y(n_2941)
);

INVx3_ASAP7_75t_L g2942 ( 
.A(n_2789),
.Y(n_2942)
);

A2O1A1Ixp33_ASAP7_75t_SL g2943 ( 
.A1(n_2738),
.A2(n_1564),
.B(n_2104),
.C(n_2101),
.Y(n_2943)
);

CKINVDCx20_ASAP7_75t_R g2944 ( 
.A(n_2701),
.Y(n_2944)
);

OA21x2_ASAP7_75t_L g2945 ( 
.A1(n_2702),
.A2(n_1605),
.B(n_2264),
.Y(n_2945)
);

AND2x2_ASAP7_75t_L g2946 ( 
.A(n_2819),
.B(n_2456),
.Y(n_2946)
);

NOR2xp67_ASAP7_75t_L g2947 ( 
.A(n_2744),
.B(n_2434),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_2755),
.B(n_2760),
.Y(n_2948)
);

HB1xp67_ASAP7_75t_L g2949 ( 
.A(n_2760),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2787),
.Y(n_2950)
);

BUFx4f_ASAP7_75t_L g2951 ( 
.A(n_2737),
.Y(n_2951)
);

AOI21xp5_ASAP7_75t_L g2952 ( 
.A1(n_2766),
.A2(n_2236),
.B(n_2137),
.Y(n_2952)
);

NOR2xp33_ASAP7_75t_L g2953 ( 
.A(n_2761),
.B(n_71),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_L g2954 ( 
.A(n_2816),
.B(n_2350),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_L g2955 ( 
.A(n_2741),
.B(n_2352),
.Y(n_2955)
);

O2A1O1Ixp5_ASAP7_75t_SL g2956 ( 
.A1(n_2821),
.A2(n_2239),
.B(n_2472),
.C(n_2442),
.Y(n_2956)
);

OA22x2_ASAP7_75t_L g2957 ( 
.A1(n_2813),
.A2(n_2361),
.B1(n_2371),
.B2(n_2356),
.Y(n_2957)
);

NOR2xp67_ASAP7_75t_SL g2958 ( 
.A(n_2843),
.B(n_2337),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2801),
.Y(n_2959)
);

BUFx3_ASAP7_75t_L g2960 ( 
.A(n_2730),
.Y(n_2960)
);

CKINVDCx10_ASAP7_75t_R g2961 ( 
.A(n_2730),
.Y(n_2961)
);

NOR2xp33_ASAP7_75t_L g2962 ( 
.A(n_2745),
.B(n_72),
.Y(n_2962)
);

BUFx6f_ASAP7_75t_L g2963 ( 
.A(n_2828),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2704),
.Y(n_2964)
);

AOI21x1_ASAP7_75t_L g2965 ( 
.A1(n_2871),
.A2(n_2264),
.B(n_1644),
.Y(n_2965)
);

AND2x2_ASAP7_75t_L g2966 ( 
.A(n_2857),
.B(n_2828),
.Y(n_2966)
);

AOI21xp5_ASAP7_75t_L g2967 ( 
.A1(n_2702),
.A2(n_2236),
.B(n_2143),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_L g2968 ( 
.A(n_2746),
.B(n_2356),
.Y(n_2968)
);

OAI21xp5_ASAP7_75t_L g2969 ( 
.A1(n_2724),
.A2(n_1644),
.B(n_2377),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2706),
.B(n_2361),
.Y(n_2970)
);

AOI22xp33_ASAP7_75t_L g2971 ( 
.A1(n_2862),
.A2(n_2402),
.B1(n_2384),
.B2(n_2377),
.Y(n_2971)
);

AND2x2_ASAP7_75t_L g2972 ( 
.A(n_2796),
.B(n_2456),
.Y(n_2972)
);

AOI21xp5_ASAP7_75t_L g2973 ( 
.A1(n_2744),
.A2(n_2143),
.B(n_2080),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_SL g2974 ( 
.A(n_2825),
.B(n_2583),
.Y(n_2974)
);

O2A1O1Ixp33_ASAP7_75t_L g2975 ( 
.A1(n_2709),
.A2(n_2472),
.B(n_2442),
.C(n_2360),
.Y(n_2975)
);

BUFx12f_ASAP7_75t_L g2976 ( 
.A(n_2863),
.Y(n_2976)
);

NOR2xp33_ASAP7_75t_L g2977 ( 
.A(n_2842),
.B(n_72),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_L g2978 ( 
.A(n_2803),
.B(n_2371),
.Y(n_2978)
);

OAI21xp33_ASAP7_75t_L g2979 ( 
.A1(n_2823),
.A2(n_1990),
.B(n_1656),
.Y(n_2979)
);

OR2x6_ASAP7_75t_SL g2980 ( 
.A(n_2844),
.B(n_2372),
.Y(n_2980)
);

AO21x1_ASAP7_75t_L g2981 ( 
.A1(n_2873),
.A2(n_2489),
.B(n_2476),
.Y(n_2981)
);

NOR2xp33_ASAP7_75t_L g2982 ( 
.A(n_2842),
.B(n_75),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2705),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_2814),
.B(n_2372),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2764),
.B(n_2375),
.Y(n_2985)
);

OAI22xp5_ASAP7_75t_L g2986 ( 
.A1(n_2769),
.A2(n_2375),
.B1(n_2387),
.B2(n_2380),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2710),
.Y(n_2987)
);

AO21x1_ASAP7_75t_L g2988 ( 
.A1(n_2709),
.A2(n_2489),
.B(n_2476),
.Y(n_2988)
);

AOI21xp5_ASAP7_75t_L g2989 ( 
.A1(n_2744),
.A2(n_2143),
.B(n_2080),
.Y(n_2989)
);

OAI22xp5_ASAP7_75t_L g2990 ( 
.A1(n_2824),
.A2(n_2387),
.B1(n_2405),
.B2(n_2390),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2732),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2743),
.Y(n_2992)
);

AOI21xp5_ASAP7_75t_L g2993 ( 
.A1(n_2744),
.A2(n_2143),
.B(n_2080),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_2792),
.Y(n_2994)
);

INVx2_ASAP7_75t_L g2995 ( 
.A(n_2794),
.Y(n_2995)
);

OAI22x1_ASAP7_75t_L g2996 ( 
.A1(n_2867),
.A2(n_2405),
.B1(n_2408),
.B2(n_2390),
.Y(n_2996)
);

NOR2xp33_ASAP7_75t_L g2997 ( 
.A(n_2707),
.B(n_75),
.Y(n_2997)
);

XOR2xp5_ASAP7_75t_L g2998 ( 
.A(n_2720),
.B(n_2337),
.Y(n_2998)
);

AOI22xp33_ASAP7_75t_L g2999 ( 
.A1(n_2879),
.A2(n_2384),
.B1(n_2377),
.B2(n_2474),
.Y(n_2999)
);

BUFx6f_ASAP7_75t_L g3000 ( 
.A(n_2759),
.Y(n_3000)
);

CKINVDCx5p33_ASAP7_75t_R g3001 ( 
.A(n_2781),
.Y(n_3001)
);

AOI21xp5_ASAP7_75t_L g3002 ( 
.A1(n_2809),
.A2(n_2837),
.B(n_2699),
.Y(n_3002)
);

A2O1A1Ixp33_ASAP7_75t_L g3003 ( 
.A1(n_2772),
.A2(n_2408),
.B(n_2420),
.C(n_2415),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_L g3004 ( 
.A(n_2721),
.B(n_2415),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_2763),
.B(n_2420),
.Y(n_3005)
);

BUFx3_ASAP7_75t_L g3006 ( 
.A(n_2811),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2783),
.B(n_2431),
.Y(n_3007)
);

NOR2xp33_ASAP7_75t_L g3008 ( 
.A(n_2703),
.B(n_76),
.Y(n_3008)
);

AO32x2_ASAP7_75t_L g3009 ( 
.A1(n_2791),
.A2(n_2440),
.A3(n_2449),
.B1(n_2441),
.B2(n_2431),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_SL g3010 ( 
.A(n_2825),
.B(n_2456),
.Y(n_3010)
);

NOR2xp33_ASAP7_75t_L g3011 ( 
.A(n_2703),
.B(n_76),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_L g3012 ( 
.A(n_2851),
.B(n_2440),
.Y(n_3012)
);

AOI22xp5_ASAP7_75t_L g3013 ( 
.A1(n_2772),
.A2(n_2077),
.B1(n_2234),
.B2(n_2039),
.Y(n_3013)
);

INVx2_ASAP7_75t_L g3014 ( 
.A(n_2794),
.Y(n_3014)
);

AOI21xp5_ASAP7_75t_L g3015 ( 
.A1(n_2809),
.A2(n_2143),
.B(n_2080),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_L g3016 ( 
.A(n_2854),
.B(n_2441),
.Y(n_3016)
);

INVx2_ASAP7_75t_L g3017 ( 
.A(n_2798),
.Y(n_3017)
);

OAI21xp5_ASAP7_75t_L g3018 ( 
.A1(n_2802),
.A2(n_1656),
.B(n_1524),
.Y(n_3018)
);

OR2x2_ASAP7_75t_L g3019 ( 
.A(n_2850),
.B(n_2449),
.Y(n_3019)
);

CKINVDCx16_ASAP7_75t_R g3020 ( 
.A(n_2796),
.Y(n_3020)
);

OAI21xp5_ASAP7_75t_L g3021 ( 
.A1(n_2802),
.A2(n_1524),
.B(n_1586),
.Y(n_3021)
);

AOI21xp5_ASAP7_75t_L g3022 ( 
.A1(n_2809),
.A2(n_2080),
.B(n_2337),
.Y(n_3022)
);

OAI22xp5_ASAP7_75t_L g3023 ( 
.A1(n_2809),
.A2(n_2451),
.B1(n_2458),
.B2(n_2455),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2757),
.Y(n_3024)
);

AO32x1_ASAP7_75t_L g3025 ( 
.A1(n_2791),
.A2(n_2455),
.A3(n_2478),
.B1(n_2458),
.B2(n_2451),
.Y(n_3025)
);

AOI21xp5_ASAP7_75t_L g3026 ( 
.A1(n_2837),
.A2(n_2359),
.B(n_2337),
.Y(n_3026)
);

NOR2xp33_ASAP7_75t_L g3027 ( 
.A(n_2806),
.B(n_78),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2836),
.B(n_2478),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_L g3029 ( 
.A(n_2836),
.B(n_2485),
.Y(n_3029)
);

AND2x2_ASAP7_75t_L g3030 ( 
.A(n_2850),
.B(n_2456),
.Y(n_3030)
);

XOR2xp5_ASAP7_75t_L g3031 ( 
.A(n_2758),
.B(n_2359),
.Y(n_3031)
);

AOI21xp5_ASAP7_75t_L g3032 ( 
.A1(n_2837),
.A2(n_2366),
.B(n_2359),
.Y(n_3032)
);

NAND2x1p5_ASAP7_75t_L g3033 ( 
.A(n_2837),
.B(n_2699),
.Y(n_3033)
);

NOR2x1_ASAP7_75t_L g3034 ( 
.A(n_2742),
.B(n_2759),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2878),
.B(n_2870),
.Y(n_3035)
);

NOR2xp33_ASAP7_75t_L g3036 ( 
.A(n_2808),
.B(n_78),
.Y(n_3036)
);

INVx2_ASAP7_75t_L g3037 ( 
.A(n_2798),
.Y(n_3037)
);

INVx2_ASAP7_75t_L g3038 ( 
.A(n_2807),
.Y(n_3038)
);

AOI21xp5_ASAP7_75t_L g3039 ( 
.A1(n_2699),
.A2(n_2366),
.B(n_2359),
.Y(n_3039)
);

A2O1A1Ixp33_ASAP7_75t_L g3040 ( 
.A1(n_2753),
.A2(n_2485),
.B(n_2227),
.C(n_2239),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_SL g3041 ( 
.A(n_2738),
.B(n_2461),
.Y(n_3041)
);

AOI21xp5_ASAP7_75t_L g3042 ( 
.A1(n_2780),
.A2(n_2379),
.B(n_2366),
.Y(n_3042)
);

NAND3xp33_ASAP7_75t_SL g3043 ( 
.A(n_2858),
.B(n_2780),
.C(n_2855),
.Y(n_3043)
);

OAI21x1_ASAP7_75t_L g3044 ( 
.A1(n_2716),
.A2(n_2460),
.B(n_2407),
.Y(n_3044)
);

NOR2xp33_ASAP7_75t_SL g3045 ( 
.A(n_2832),
.B(n_2461),
.Y(n_3045)
);

OAI22xp5_ASAP7_75t_L g3046 ( 
.A1(n_2776),
.A2(n_2283),
.B1(n_2281),
.B2(n_2278),
.Y(n_3046)
);

INVx2_ASAP7_75t_L g3047 ( 
.A(n_2807),
.Y(n_3047)
);

BUFx3_ASAP7_75t_L g3048 ( 
.A(n_2777),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_SL g3049 ( 
.A(n_2812),
.B(n_2461),
.Y(n_3049)
);

NOR2xp33_ASAP7_75t_L g3050 ( 
.A(n_2800),
.B(n_80),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_2860),
.B(n_2463),
.Y(n_3051)
);

NAND2xp5_ASAP7_75t_L g3052 ( 
.A(n_2864),
.B(n_2463),
.Y(n_3052)
);

BUFx2_ASAP7_75t_L g3053 ( 
.A(n_2777),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_SL g3054 ( 
.A(n_2812),
.B(n_2463),
.Y(n_3054)
);

O2A1O1Ixp5_ASAP7_75t_L g3055 ( 
.A1(n_2876),
.A2(n_2360),
.B(n_2376),
.C(n_2340),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_SL g3056 ( 
.A(n_2812),
.B(n_2463),
.Y(n_3056)
);

NAND2xp5_ASAP7_75t_SL g3057 ( 
.A(n_2812),
.B(n_2366),
.Y(n_3057)
);

NOR2xp33_ASAP7_75t_L g3058 ( 
.A(n_2751),
.B(n_80),
.Y(n_3058)
);

AND2x2_ASAP7_75t_L g3059 ( 
.A(n_2742),
.B(n_2765),
.Y(n_3059)
);

AOI22xp33_ASAP7_75t_L g3060 ( 
.A1(n_2768),
.A2(n_2494),
.B1(n_2496),
.B2(n_2480),
.Y(n_3060)
);

NAND2xp5_ASAP7_75t_L g3061 ( 
.A(n_2869),
.B(n_2504),
.Y(n_3061)
);

INVx4_ASAP7_75t_L g3062 ( 
.A(n_2747),
.Y(n_3062)
);

INVx2_ASAP7_75t_L g3063 ( 
.A(n_2771),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_L g3064 ( 
.A(n_2773),
.B(n_2505),
.Y(n_3064)
);

A2O1A1Ixp33_ASAP7_75t_SL g3065 ( 
.A1(n_2751),
.A2(n_2104),
.B(n_2111),
.C(n_2101),
.Y(n_3065)
);

OAI22xp5_ASAP7_75t_L g3066 ( 
.A1(n_2776),
.A2(n_2283),
.B1(n_2281),
.B2(n_2278),
.Y(n_3066)
);

AOI31xp67_ASAP7_75t_L g3067 ( 
.A1(n_3041),
.A2(n_2878),
.A3(n_2845),
.B(n_2875),
.Y(n_3067)
);

NOR2xp33_ASAP7_75t_L g3068 ( 
.A(n_2884),
.B(n_2747),
.Y(n_3068)
);

AOI21xp5_ASAP7_75t_L g3069 ( 
.A1(n_2895),
.A2(n_2876),
.B(n_2727),
.Y(n_3069)
);

OAI21xp5_ASAP7_75t_L g3070 ( 
.A1(n_2913),
.A2(n_2804),
.B(n_2779),
.Y(n_3070)
);

AOI21xp5_ASAP7_75t_L g3071 ( 
.A1(n_2887),
.A2(n_2891),
.B(n_2907),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2881),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2888),
.B(n_2874),
.Y(n_3073)
);

NOR2x1_ASAP7_75t_SL g3074 ( 
.A(n_2905),
.B(n_2832),
.Y(n_3074)
);

OAI22xp5_ASAP7_75t_L g3075 ( 
.A1(n_2880),
.A2(n_2868),
.B1(n_2832),
.B2(n_2849),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2909),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_L g3077 ( 
.A(n_2883),
.B(n_2845),
.Y(n_3077)
);

INVxp67_ASAP7_75t_L g3078 ( 
.A(n_2963),
.Y(n_3078)
);

OAI21x1_ASAP7_75t_L g3079 ( 
.A1(n_2956),
.A2(n_2716),
.B(n_2841),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2898),
.Y(n_3080)
);

OAI21x1_ASAP7_75t_L g3081 ( 
.A1(n_2917),
.A2(n_2841),
.B(n_2872),
.Y(n_3081)
);

BUFx3_ASAP7_75t_L g3082 ( 
.A(n_2912),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2948),
.B(n_2870),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_SL g3084 ( 
.A(n_3020),
.B(n_2737),
.Y(n_3084)
);

AND2x2_ASAP7_75t_L g3085 ( 
.A(n_2938),
.B(n_2868),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_2948),
.B(n_2872),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2902),
.Y(n_3087)
);

NAND3xp33_ASAP7_75t_L g3088 ( 
.A(n_2953),
.B(n_2925),
.C(n_2977),
.Y(n_3088)
);

INVx6_ASAP7_75t_L g3089 ( 
.A(n_2963),
.Y(n_3089)
);

CKINVDCx20_ASAP7_75t_R g3090 ( 
.A(n_2903),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_L g3091 ( 
.A(n_2918),
.B(n_2875),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_L g3092 ( 
.A(n_2949),
.B(n_2768),
.Y(n_3092)
);

AOI22x1_ASAP7_75t_L g3093 ( 
.A1(n_3001),
.A2(n_2719),
.B1(n_2756),
.B2(n_2752),
.Y(n_3093)
);

BUFx3_ASAP7_75t_L g3094 ( 
.A(n_2944),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_2924),
.B(n_2768),
.Y(n_3095)
);

NOR2x1_ASAP7_75t_SL g3096 ( 
.A(n_2941),
.B(n_2832),
.Y(n_3096)
);

HB1xp67_ASAP7_75t_L g3097 ( 
.A(n_3059),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_2959),
.B(n_2768),
.Y(n_3098)
);

NAND2xp5_ASAP7_75t_SL g3099 ( 
.A(n_2963),
.B(n_2815),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_2964),
.B(n_2768),
.Y(n_3100)
);

BUFx2_ASAP7_75t_L g3101 ( 
.A(n_3006),
.Y(n_3101)
);

OAI21x1_ASAP7_75t_L g3102 ( 
.A1(n_3002),
.A2(n_2838),
.B(n_2820),
.Y(n_3102)
);

OAI21xp5_ASAP7_75t_L g3103 ( 
.A1(n_2897),
.A2(n_2810),
.B(n_2853),
.Y(n_3103)
);

OAI21x1_ASAP7_75t_L g3104 ( 
.A1(n_2965),
.A2(n_2838),
.B(n_2820),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_L g3105 ( 
.A(n_2983),
.B(n_2700),
.Y(n_3105)
);

OAI21x1_ASAP7_75t_L g3106 ( 
.A1(n_2885),
.A2(n_2827),
.B(n_2793),
.Y(n_3106)
);

AOI221x1_ASAP7_75t_L g3107 ( 
.A1(n_3043),
.A2(n_2982),
.B1(n_3008),
.B2(n_3011),
.C(n_3058),
.Y(n_3107)
);

AOI21xp5_ASAP7_75t_L g3108 ( 
.A1(n_2934),
.A2(n_2810),
.B(n_2793),
.Y(n_3108)
);

OAI21x1_ASAP7_75t_L g3109 ( 
.A1(n_2952),
.A2(n_2929),
.B(n_2937),
.Y(n_3109)
);

INVx2_ASAP7_75t_L g3110 ( 
.A(n_3063),
.Y(n_3110)
);

AND2x4_ASAP7_75t_L g3111 ( 
.A(n_3030),
.B(n_2868),
.Y(n_3111)
);

BUFx12f_ASAP7_75t_L g3112 ( 
.A(n_2976),
.Y(n_3112)
);

INVx2_ASAP7_75t_L g3113 ( 
.A(n_2886),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_2920),
.B(n_2777),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_L g3115 ( 
.A(n_2987),
.B(n_2752),
.Y(n_3115)
);

INVx2_ASAP7_75t_SL g3116 ( 
.A(n_2966),
.Y(n_3116)
);

BUFx2_ASAP7_75t_L g3117 ( 
.A(n_3053),
.Y(n_3117)
);

NOR2xp33_ASAP7_75t_L g3118 ( 
.A(n_2894),
.B(n_2747),
.Y(n_3118)
);

OAI21x1_ASAP7_75t_L g3119 ( 
.A1(n_2929),
.A2(n_2829),
.B(n_2827),
.Y(n_3119)
);

O2A1O1Ixp5_ASAP7_75t_L g3120 ( 
.A1(n_2925),
.A2(n_2756),
.B(n_2784),
.C(n_2767),
.Y(n_3120)
);

O2A1O1Ixp5_ASAP7_75t_L g3121 ( 
.A1(n_2988),
.A2(n_2928),
.B(n_3050),
.C(n_3027),
.Y(n_3121)
);

AOI22xp5_ASAP7_75t_L g3122 ( 
.A1(n_2899),
.A2(n_2719),
.B1(n_2849),
.B2(n_2859),
.Y(n_3122)
);

AO21x1_ASAP7_75t_L g3123 ( 
.A1(n_2928),
.A2(n_2859),
.B(n_2805),
.Y(n_3123)
);

INVx5_ASAP7_75t_L g3124 ( 
.A(n_3000),
.Y(n_3124)
);

OAI21x1_ASAP7_75t_L g3125 ( 
.A1(n_3021),
.A2(n_2834),
.B(n_2829),
.Y(n_3125)
);

AO21x2_ASAP7_75t_L g3126 ( 
.A1(n_3023),
.A2(n_2712),
.B(n_2700),
.Y(n_3126)
);

BUFx5_ASAP7_75t_L g3127 ( 
.A(n_2972),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_L g3128 ( 
.A(n_2991),
.B(n_2712),
.Y(n_3128)
);

INVx3_ASAP7_75t_L g3129 ( 
.A(n_2904),
.Y(n_3129)
);

CKINVDCx14_ASAP7_75t_R g3130 ( 
.A(n_3048),
.Y(n_3130)
);

OAI21x1_ASAP7_75t_L g3131 ( 
.A1(n_3021),
.A2(n_2835),
.B(n_2834),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_L g3132 ( 
.A(n_2992),
.B(n_2713),
.Y(n_3132)
);

OA22x2_ASAP7_75t_L g3133 ( 
.A1(n_2889),
.A2(n_2849),
.B1(n_2778),
.B2(n_2805),
.Y(n_3133)
);

OAI21xp5_ASAP7_75t_L g3134 ( 
.A1(n_2931),
.A2(n_2835),
.B(n_2407),
.Y(n_3134)
);

OAI21x1_ASAP7_75t_L g3135 ( 
.A1(n_2969),
.A2(n_2714),
.B(n_2713),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_3024),
.B(n_2714),
.Y(n_3136)
);

AO21x1_ASAP7_75t_L g3137 ( 
.A1(n_2899),
.A2(n_2805),
.B(n_2778),
.Y(n_3137)
);

BUFx6f_ASAP7_75t_L g3138 ( 
.A(n_3000),
.Y(n_3138)
);

NAND3xp33_ASAP7_75t_L g3139 ( 
.A(n_2997),
.B(n_2784),
.C(n_2815),
.Y(n_3139)
);

AOI21xp5_ASAP7_75t_L g3140 ( 
.A1(n_3010),
.A2(n_2868),
.B(n_2778),
.Y(n_3140)
);

NAND3xp33_ASAP7_75t_L g3141 ( 
.A(n_2962),
.B(n_2815),
.C(n_2782),
.Y(n_3141)
);

AOI21x1_ASAP7_75t_L g3142 ( 
.A1(n_2958),
.A2(n_2717),
.B(n_2715),
.Y(n_3142)
);

NAND2x1_ASAP7_75t_L g3143 ( 
.A(n_2904),
.B(n_2942),
.Y(n_3143)
);

NOR2xp67_ASAP7_75t_L g3144 ( 
.A(n_3062),
.B(n_2815),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_3035),
.B(n_2715),
.Y(n_3145)
);

AOI21xp5_ASAP7_75t_L g3146 ( 
.A1(n_2923),
.A2(n_2399),
.B(n_2379),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_L g3147 ( 
.A(n_3035),
.B(n_2717),
.Y(n_3147)
);

BUFx6f_ASAP7_75t_L g3148 ( 
.A(n_3000),
.Y(n_3148)
);

OAI21x1_ASAP7_75t_L g3149 ( 
.A1(n_2969),
.A2(n_2733),
.B(n_2725),
.Y(n_3149)
);

AO31x2_ASAP7_75t_L g3150 ( 
.A1(n_3023),
.A2(n_2733),
.A3(n_2734),
.B(n_2725),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_3019),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_2935),
.B(n_2734),
.Y(n_3152)
);

AO22x2_ASAP7_75t_L g3153 ( 
.A1(n_2914),
.A2(n_2750),
.B1(n_2754),
.B2(n_2740),
.Y(n_3153)
);

OAI21x1_ASAP7_75t_L g3154 ( 
.A1(n_3026),
.A2(n_2750),
.B(n_2740),
.Y(n_3154)
);

OAI21x1_ASAP7_75t_L g3155 ( 
.A1(n_3032),
.A2(n_2967),
.B(n_3022),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_3064),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_SL g3157 ( 
.A(n_3062),
.B(n_2782),
.Y(n_3157)
);

OAI21x1_ASAP7_75t_L g3158 ( 
.A1(n_2973),
.A2(n_2770),
.B(n_2754),
.Y(n_3158)
);

NOR2xp67_ASAP7_75t_L g3159 ( 
.A(n_2906),
.B(n_2901),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_L g3160 ( 
.A(n_2930),
.B(n_2770),
.Y(n_3160)
);

OAI21x1_ASAP7_75t_L g3161 ( 
.A1(n_2989),
.A2(n_2774),
.B(n_2300),
.Y(n_3161)
);

AOI21x1_ASAP7_75t_L g3162 ( 
.A1(n_3042),
.A2(n_2774),
.B(n_2512),
.Y(n_3162)
);

AOI21x1_ASAP7_75t_L g3163 ( 
.A1(n_3057),
.A2(n_2507),
.B(n_1496),
.Y(n_3163)
);

OAI21x1_ASAP7_75t_L g3164 ( 
.A1(n_2993),
.A2(n_2376),
.B(n_2340),
.Y(n_3164)
);

OAI21xp5_ASAP7_75t_L g3165 ( 
.A1(n_2923),
.A2(n_1985),
.B(n_1982),
.Y(n_3165)
);

INVx2_ASAP7_75t_L g3166 ( 
.A(n_2908),
.Y(n_3166)
);

OR2x2_ASAP7_75t_L g3167 ( 
.A(n_3005),
.B(n_2775),
.Y(n_3167)
);

AO31x2_ASAP7_75t_L g3168 ( 
.A1(n_2996),
.A2(n_2762),
.A3(n_2279),
.B(n_2249),
.Y(n_3168)
);

AO21x1_ASAP7_75t_L g3169 ( 
.A1(n_2921),
.A2(n_2762),
.B(n_81),
.Y(n_3169)
);

AO31x2_ASAP7_75t_L g3170 ( 
.A1(n_2981),
.A2(n_2279),
.A3(n_2249),
.B(n_2010),
.Y(n_3170)
);

BUFx3_ASAP7_75t_L g3171 ( 
.A(n_2960),
.Y(n_3171)
);

OAI22xp5_ASAP7_75t_L g3172 ( 
.A1(n_2971),
.A2(n_2782),
.B1(n_2775),
.B2(n_2401),
.Y(n_3172)
);

OAI21x1_ASAP7_75t_L g3173 ( 
.A1(n_3015),
.A2(n_2401),
.B(n_2400),
.Y(n_3173)
);

AOI21xp5_ASAP7_75t_L g3174 ( 
.A1(n_2974),
.A2(n_2399),
.B(n_2379),
.Y(n_3174)
);

NAND3x1_ASAP7_75t_L g3175 ( 
.A(n_2911),
.B(n_2430),
.C(n_2400),
.Y(n_3175)
);

OAI21x1_ASAP7_75t_L g3176 ( 
.A1(n_3018),
.A2(n_2430),
.B(n_1427),
.Y(n_3176)
);

O2A1O1Ixp5_ASAP7_75t_SL g3177 ( 
.A1(n_3049),
.A2(n_2243),
.B(n_2230),
.C(n_2212),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_3028),
.Y(n_3178)
);

NAND2x1p5_ASAP7_75t_L g3179 ( 
.A(n_2951),
.B(n_2782),
.Y(n_3179)
);

INVx2_ASAP7_75t_L g3180 ( 
.A(n_2950),
.Y(n_3180)
);

OAI21x1_ASAP7_75t_L g3181 ( 
.A1(n_3018),
.A2(n_2243),
.B(n_2230),
.Y(n_3181)
);

INVx1_ASAP7_75t_SL g3182 ( 
.A(n_2980),
.Y(n_3182)
);

CKINVDCx5p33_ASAP7_75t_R g3183 ( 
.A(n_2961),
.Y(n_3183)
);

OAI21x1_ASAP7_75t_L g3184 ( 
.A1(n_3033),
.A2(n_2243),
.B(n_2230),
.Y(n_3184)
);

BUFx2_ASAP7_75t_L g3185 ( 
.A(n_2936),
.Y(n_3185)
);

OAI21x1_ASAP7_75t_L g3186 ( 
.A1(n_3033),
.A2(n_1543),
.B(n_1532),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_2926),
.B(n_2775),
.Y(n_3187)
);

OAI21x1_ASAP7_75t_L g3188 ( 
.A1(n_3039),
.A2(n_1543),
.B(n_1532),
.Y(n_3188)
);

AND2x2_ASAP7_75t_L g3189 ( 
.A(n_2946),
.B(n_2775),
.Y(n_3189)
);

BUFx2_ASAP7_75t_L g3190 ( 
.A(n_2942),
.Y(n_3190)
);

OAI21xp5_ASAP7_75t_L g3191 ( 
.A1(n_2921),
.A2(n_1971),
.B(n_1924),
.Y(n_3191)
);

A2O1A1Ixp33_ASAP7_75t_L g3192 ( 
.A1(n_2910),
.A2(n_1942),
.B(n_1946),
.C(n_1938),
.Y(n_3192)
);

HB1xp67_ASAP7_75t_L g3193 ( 
.A(n_3007),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_3028),
.Y(n_3194)
);

AND2x4_ASAP7_75t_L g3195 ( 
.A(n_3034),
.B(n_2379),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_L g3196 ( 
.A(n_2927),
.B(n_2399),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_L g3197 ( 
.A(n_2978),
.B(n_2399),
.Y(n_3197)
);

AOI21xp33_ASAP7_75t_L g3198 ( 
.A1(n_2939),
.A2(n_2427),
.B(n_2414),
.Y(n_3198)
);

NOR2x1_ASAP7_75t_SL g3199 ( 
.A(n_2882),
.B(n_2403),
.Y(n_3199)
);

OAI21x1_ASAP7_75t_L g3200 ( 
.A1(n_3044),
.A2(n_2212),
.B(n_2204),
.Y(n_3200)
);

INVx3_ASAP7_75t_L g3201 ( 
.A(n_2951),
.Y(n_3201)
);

INVxp67_ASAP7_75t_SL g3202 ( 
.A(n_3051),
.Y(n_3202)
);

INVx4_ASAP7_75t_L g3203 ( 
.A(n_2945),
.Y(n_3203)
);

OAI21x1_ASAP7_75t_L g3204 ( 
.A1(n_3055),
.A2(n_2212),
.B(n_2204),
.Y(n_3204)
);

OAI21x1_ASAP7_75t_L g3205 ( 
.A1(n_2939),
.A2(n_2204),
.B(n_2039),
.Y(n_3205)
);

AO31x2_ASAP7_75t_L g3206 ( 
.A1(n_2990),
.A2(n_2010),
.A3(n_2014),
.B(n_2012),
.Y(n_3206)
);

AO31x2_ASAP7_75t_L g3207 ( 
.A1(n_2990),
.A2(n_2012),
.A3(n_2015),
.B(n_2014),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_2970),
.B(n_81),
.Y(n_3208)
);

BUFx6f_ASAP7_75t_L g3209 ( 
.A(n_3054),
.Y(n_3209)
);

A2O1A1Ixp33_ASAP7_75t_L g3210 ( 
.A1(n_2916),
.A2(n_1942),
.B(n_1946),
.C(n_1938),
.Y(n_3210)
);

OR2x2_ASAP7_75t_L g3211 ( 
.A(n_2896),
.B(n_82),
.Y(n_3211)
);

OAI21x1_ASAP7_75t_L g3212 ( 
.A1(n_2890),
.A2(n_2026),
.B(n_2111),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_3029),
.Y(n_3213)
);

OAI21x1_ASAP7_75t_L g3214 ( 
.A1(n_2940),
.A2(n_2979),
.B(n_2932),
.Y(n_3214)
);

OAI21x1_ASAP7_75t_L g3215 ( 
.A1(n_2945),
.A2(n_2136),
.B(n_2113),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_L g3216 ( 
.A(n_2955),
.B(n_2414),
.Y(n_3216)
);

AOI21xp5_ASAP7_75t_L g3217 ( 
.A1(n_2943),
.A2(n_2423),
.B(n_2414),
.Y(n_3217)
);

OAI21x1_ASAP7_75t_L g3218 ( 
.A1(n_2922),
.A2(n_2136),
.B(n_2113),
.Y(n_3218)
);

OAI21x1_ASAP7_75t_L g3219 ( 
.A1(n_2892),
.A2(n_2136),
.B(n_2113),
.Y(n_3219)
);

HB1xp67_ASAP7_75t_L g3220 ( 
.A(n_3052),
.Y(n_3220)
);

OAI21x1_ASAP7_75t_L g3221 ( 
.A1(n_3056),
.A2(n_2975),
.B(n_3060),
.Y(n_3221)
);

OAI21xp5_ASAP7_75t_L g3222 ( 
.A1(n_2933),
.A2(n_1951),
.B(n_1949),
.Y(n_3222)
);

CKINVDCx12_ASAP7_75t_R g3223 ( 
.A(n_2994),
.Y(n_3223)
);

INVx2_ASAP7_75t_L g3224 ( 
.A(n_2995),
.Y(n_3224)
);

OAI21x1_ASAP7_75t_L g3225 ( 
.A1(n_3046),
.A2(n_3066),
.B(n_3061),
.Y(n_3225)
);

BUFx4_ASAP7_75t_SL g3226 ( 
.A(n_3031),
.Y(n_3226)
);

CKINVDCx14_ASAP7_75t_R g3227 ( 
.A(n_2998),
.Y(n_3227)
);

AOI21x1_ASAP7_75t_L g3228 ( 
.A1(n_2947),
.A2(n_2017),
.B(n_2015),
.Y(n_3228)
);

AOI21xp5_ASAP7_75t_L g3229 ( 
.A1(n_3065),
.A2(n_2423),
.B(n_2414),
.Y(n_3229)
);

OAI21xp5_ASAP7_75t_L g3230 ( 
.A1(n_2986),
.A2(n_1951),
.B(n_1949),
.Y(n_3230)
);

HB1xp67_ASAP7_75t_L g3231 ( 
.A(n_2968),
.Y(n_3231)
);

OAI21x1_ASAP7_75t_L g3232 ( 
.A1(n_3046),
.A2(n_2149),
.B(n_2139),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_3029),
.B(n_2423),
.Y(n_3233)
);

AND2x2_ASAP7_75t_L g3234 ( 
.A(n_2919),
.B(n_2423),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_2954),
.Y(n_3235)
);

INVxp67_ASAP7_75t_L g3236 ( 
.A(n_2985),
.Y(n_3236)
);

INVx3_ASAP7_75t_L g3237 ( 
.A(n_2957),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_3004),
.B(n_2425),
.Y(n_3238)
);

AND2x2_ASAP7_75t_L g3239 ( 
.A(n_3036),
.B(n_2425),
.Y(n_3239)
);

O2A1O1Ixp5_ASAP7_75t_L g3240 ( 
.A1(n_2986),
.A2(n_2149),
.B(n_2165),
.C(n_2139),
.Y(n_3240)
);

AO31x2_ASAP7_75t_L g3241 ( 
.A1(n_3066),
.A2(n_2017),
.A3(n_2022),
.B(n_2019),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_L g3242 ( 
.A(n_2984),
.B(n_3012),
.Y(n_3242)
);

AOI21xp5_ASAP7_75t_L g3243 ( 
.A1(n_3045),
.A2(n_2427),
.B(n_2425),
.Y(n_3243)
);

OAI21x1_ASAP7_75t_L g3244 ( 
.A1(n_2957),
.A2(n_2149),
.B(n_2139),
.Y(n_3244)
);

AND2x4_ASAP7_75t_L g3245 ( 
.A(n_3047),
.B(n_2427),
.Y(n_3245)
);

AND2x2_ASAP7_75t_L g3246 ( 
.A(n_2999),
.B(n_3014),
.Y(n_3246)
);

O2A1O1Ixp5_ASAP7_75t_L g3247 ( 
.A1(n_2914),
.A2(n_2168),
.B(n_2173),
.C(n_2165),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_3016),
.Y(n_3248)
);

AOI21xp5_ASAP7_75t_L g3249 ( 
.A1(n_3045),
.A2(n_2427),
.B(n_2168),
.Y(n_3249)
);

NOR2xp33_ASAP7_75t_L g3250 ( 
.A(n_3013),
.B(n_82),
.Y(n_3250)
);

NAND2xp33_ASAP7_75t_L g3251 ( 
.A(n_2900),
.B(n_3040),
.Y(n_3251)
);

AND2x2_ASAP7_75t_L g3252 ( 
.A(n_3017),
.B(n_83),
.Y(n_3252)
);

AND2x4_ASAP7_75t_L g3253 ( 
.A(n_3038),
.B(n_2233),
.Y(n_3253)
);

NOR2x1_ASAP7_75t_SL g3254 ( 
.A(n_3037),
.B(n_2087),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_L g3255 ( 
.A(n_3003),
.B(n_85),
.Y(n_3255)
);

AND2x2_ASAP7_75t_L g3256 ( 
.A(n_2893),
.B(n_85),
.Y(n_3256)
);

O2A1O1Ixp5_ASAP7_75t_L g3257 ( 
.A1(n_2915),
.A2(n_2168),
.B(n_2173),
.C(n_2165),
.Y(n_3257)
);

AOI21xp5_ASAP7_75t_L g3258 ( 
.A1(n_2915),
.A2(n_2173),
.B(n_2124),
.Y(n_3258)
);

OAI22xp5_ASAP7_75t_L g3259 ( 
.A1(n_2915),
.A2(n_2087),
.B1(n_2150),
.B2(n_2124),
.Y(n_3259)
);

NAND2xp5_ASAP7_75t_L g3260 ( 
.A(n_3009),
.B(n_86),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_L g3261 ( 
.A(n_3009),
.B(n_87),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_SL g3262 ( 
.A(n_3025),
.B(n_2233),
.Y(n_3262)
);

AOI21x1_ASAP7_75t_L g3263 ( 
.A1(n_3025),
.A2(n_2022),
.B(n_2019),
.Y(n_3263)
);

AND2x2_ASAP7_75t_L g3264 ( 
.A(n_3009),
.B(n_87),
.Y(n_3264)
);

NOR2xp67_ASAP7_75t_L g3265 ( 
.A(n_3139),
.B(n_88),
.Y(n_3265)
);

OAI21x1_ASAP7_75t_SL g3266 ( 
.A1(n_3123),
.A2(n_89),
.B(n_90),
.Y(n_3266)
);

NOR2xp33_ASAP7_75t_SL g3267 ( 
.A(n_3090),
.B(n_2234),
.Y(n_3267)
);

OAI21x1_ASAP7_75t_L g3268 ( 
.A1(n_3263),
.A2(n_3025),
.B(n_2025),
.Y(n_3268)
);

A2O1A1Ixp33_ASAP7_75t_L g3269 ( 
.A1(n_3121),
.A2(n_2227),
.B(n_91),
.C(n_89),
.Y(n_3269)
);

AOI21xp5_ASAP7_75t_L g3270 ( 
.A1(n_3071),
.A2(n_2182),
.B(n_2174),
.Y(n_3270)
);

NAND2x1p5_ASAP7_75t_L g3271 ( 
.A(n_3124),
.B(n_3201),
.Y(n_3271)
);

OAI21x1_ASAP7_75t_L g3272 ( 
.A1(n_3079),
.A2(n_2025),
.B(n_2023),
.Y(n_3272)
);

AO31x2_ASAP7_75t_L g3273 ( 
.A1(n_3169),
.A2(n_2052),
.A3(n_2053),
.B(n_2023),
.Y(n_3273)
);

OAI21x1_ASAP7_75t_L g3274 ( 
.A1(n_3155),
.A2(n_2053),
.B(n_2052),
.Y(n_3274)
);

OAI21x1_ASAP7_75t_L g3275 ( 
.A1(n_3109),
.A2(n_2057),
.B(n_2055),
.Y(n_3275)
);

AND2x2_ASAP7_75t_L g3276 ( 
.A(n_3097),
.B(n_90),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_L g3277 ( 
.A(n_3073),
.B(n_92),
.Y(n_3277)
);

OAI21xp5_ASAP7_75t_L g3278 ( 
.A1(n_3088),
.A2(n_92),
.B(n_93),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_3220),
.B(n_93),
.Y(n_3279)
);

OAI22xp5_ASAP7_75t_L g3280 ( 
.A1(n_3088),
.A2(n_2087),
.B1(n_2150),
.B2(n_2124),
.Y(n_3280)
);

NOR2xp33_ASAP7_75t_L g3281 ( 
.A(n_3171),
.B(n_94),
.Y(n_3281)
);

AND2x4_ASAP7_75t_L g3282 ( 
.A(n_3085),
.B(n_95),
.Y(n_3282)
);

AOI21xp5_ASAP7_75t_L g3283 ( 
.A1(n_3251),
.A2(n_2182),
.B(n_2174),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_3193),
.B(n_95),
.Y(n_3284)
);

NAND3x1_ASAP7_75t_L g3285 ( 
.A(n_3118),
.B(n_97),
.C(n_99),
.Y(n_3285)
);

OAI21xp5_ASAP7_75t_L g3286 ( 
.A1(n_3107),
.A2(n_99),
.B(n_100),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_SL g3287 ( 
.A(n_3159),
.B(n_2233),
.Y(n_3287)
);

AOI21xp5_ASAP7_75t_L g3288 ( 
.A1(n_3247),
.A2(n_2182),
.B(n_2174),
.Y(n_3288)
);

BUFx2_ASAP7_75t_L g3289 ( 
.A(n_3078),
.Y(n_3289)
);

AOI21xp5_ASAP7_75t_L g3290 ( 
.A1(n_3255),
.A2(n_2182),
.B(n_2174),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_L g3291 ( 
.A(n_3202),
.B(n_100),
.Y(n_3291)
);

OAI22xp5_ASAP7_75t_L g3292 ( 
.A1(n_3122),
.A2(n_2087),
.B1(n_2150),
.B2(n_2124),
.Y(n_3292)
);

AO31x2_ASAP7_75t_L g3293 ( 
.A1(n_3137),
.A2(n_2057),
.A3(n_2058),
.B(n_2055),
.Y(n_3293)
);

AO31x2_ASAP7_75t_L g3294 ( 
.A1(n_3260),
.A2(n_3261),
.A3(n_3254),
.B(n_3203),
.Y(n_3294)
);

AOI21xp33_ASAP7_75t_L g3295 ( 
.A1(n_3182),
.A2(n_2241),
.B(n_2233),
.Y(n_3295)
);

AOI21xp5_ASAP7_75t_L g3296 ( 
.A1(n_3255),
.A2(n_2182),
.B(n_2174),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_L g3297 ( 
.A(n_3083),
.B(n_3231),
.Y(n_3297)
);

BUFx3_ASAP7_75t_L g3298 ( 
.A(n_3082),
.Y(n_3298)
);

AOI31xp67_ASAP7_75t_L g3299 ( 
.A1(n_3262),
.A2(n_2059),
.A3(n_2065),
.B(n_2058),
.Y(n_3299)
);

OR2x2_ASAP7_75t_L g3300 ( 
.A(n_3083),
.B(n_3072),
.Y(n_3300)
);

AO31x2_ASAP7_75t_L g3301 ( 
.A1(n_3203),
.A2(n_2065),
.A3(n_2069),
.B(n_2059),
.Y(n_3301)
);

OAI21x1_ASAP7_75t_L g3302 ( 
.A1(n_3120),
.A2(n_2074),
.B(n_2069),
.Y(n_3302)
);

AOI21xp5_ASAP7_75t_L g3303 ( 
.A1(n_3240),
.A2(n_2225),
.B(n_2150),
.Y(n_3303)
);

AOI21xp5_ASAP7_75t_L g3304 ( 
.A1(n_3069),
.A2(n_2225),
.B(n_2150),
.Y(n_3304)
);

INVx3_ASAP7_75t_L g3305 ( 
.A(n_3089),
.Y(n_3305)
);

OAI22xp5_ASAP7_75t_L g3306 ( 
.A1(n_3250),
.A2(n_2124),
.B1(n_2225),
.B2(n_2233),
.Y(n_3306)
);

A2O1A1Ixp33_ASAP7_75t_L g3307 ( 
.A1(n_3256),
.A2(n_104),
.B(n_101),
.C(n_102),
.Y(n_3307)
);

O2A1O1Ixp33_ASAP7_75t_L g3308 ( 
.A1(n_3208),
.A2(n_108),
.B(n_101),
.C(n_106),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_3156),
.B(n_106),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_3086),
.B(n_109),
.Y(n_3310)
);

INVx2_ASAP7_75t_L g3311 ( 
.A(n_3110),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_L g3312 ( 
.A(n_3086),
.B(n_109),
.Y(n_3312)
);

OAI21xp5_ASAP7_75t_L g3313 ( 
.A1(n_3139),
.A2(n_3225),
.B(n_3070),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_3080),
.Y(n_3314)
);

AO21x2_ASAP7_75t_L g3315 ( 
.A1(n_3264),
.A2(n_2091),
.B(n_2074),
.Y(n_3315)
);

NOR2xp33_ASAP7_75t_L g3316 ( 
.A(n_3130),
.B(n_3094),
.Y(n_3316)
);

OA21x2_ASAP7_75t_L g3317 ( 
.A1(n_3257),
.A2(n_2102),
.B(n_2091),
.Y(n_3317)
);

NAND2x1p5_ASAP7_75t_L g3318 ( 
.A(n_3124),
.B(n_2241),
.Y(n_3318)
);

AOI21xp5_ASAP7_75t_L g3319 ( 
.A1(n_3108),
.A2(n_2225),
.B(n_2241),
.Y(n_3319)
);

AOI221x1_ASAP7_75t_L g3320 ( 
.A1(n_3141),
.A2(n_2241),
.B1(n_2225),
.B2(n_1099),
.C(n_2122),
.Y(n_3320)
);

BUFx6f_ASAP7_75t_L g3321 ( 
.A(n_3138),
.Y(n_3321)
);

BUFx3_ASAP7_75t_L g3322 ( 
.A(n_3112),
.Y(n_3322)
);

AOI21xp5_ASAP7_75t_L g3323 ( 
.A1(n_3229),
.A2(n_2241),
.B(n_2103),
.Y(n_3323)
);

NOR2xp67_ASAP7_75t_L g3324 ( 
.A(n_3141),
.B(n_110),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_3087),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_3076),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_3091),
.Y(n_3327)
);

AOI21xp5_ASAP7_75t_L g3328 ( 
.A1(n_3243),
.A2(n_3214),
.B(n_3146),
.Y(n_3328)
);

OAI21x1_ASAP7_75t_L g3329 ( 
.A1(n_3162),
.A2(n_2103),
.B(n_2102),
.Y(n_3329)
);

INVx5_ASAP7_75t_L g3330 ( 
.A(n_3138),
.Y(n_3330)
);

BUFx2_ASAP7_75t_L g3331 ( 
.A(n_3101),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_3236),
.B(n_110),
.Y(n_3332)
);

CKINVDCx11_ASAP7_75t_R g3333 ( 
.A(n_3117),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3145),
.Y(n_3334)
);

AOI21xp5_ASAP7_75t_L g3335 ( 
.A1(n_3134),
.A2(n_2122),
.B(n_2119),
.Y(n_3335)
);

NAND2x1p5_ASAP7_75t_L g3336 ( 
.A(n_3124),
.B(n_3201),
.Y(n_3336)
);

OAI21x1_ASAP7_75t_L g3337 ( 
.A1(n_3104),
.A2(n_2123),
.B(n_2119),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_3077),
.B(n_111),
.Y(n_3338)
);

INVx5_ASAP7_75t_L g3339 ( 
.A(n_3138),
.Y(n_3339)
);

O2A1O1Ixp33_ASAP7_75t_L g3340 ( 
.A1(n_3210),
.A2(n_115),
.B(n_112),
.C(n_114),
.Y(n_3340)
);

AOI21xp5_ASAP7_75t_SL g3341 ( 
.A1(n_3074),
.A2(n_1558),
.B(n_1571),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_3091),
.B(n_114),
.Y(n_3342)
);

AO31x2_ASAP7_75t_L g3343 ( 
.A1(n_3075),
.A2(n_2123),
.A3(n_118),
.B(n_115),
.Y(n_3343)
);

AO21x2_ASAP7_75t_L g3344 ( 
.A1(n_3145),
.A2(n_3147),
.B(n_3126),
.Y(n_3344)
);

AOI21xp5_ASAP7_75t_L g3345 ( 
.A1(n_3134),
.A2(n_1578),
.B(n_1558),
.Y(n_3345)
);

AND2x2_ASAP7_75t_L g3346 ( 
.A(n_3185),
.B(n_117),
.Y(n_3346)
);

NOR3xp33_ASAP7_75t_L g3347 ( 
.A(n_3221),
.B(n_117),
.C(n_118),
.Y(n_3347)
);

OAI21xp5_ASAP7_75t_L g3348 ( 
.A1(n_3175),
.A2(n_3182),
.B(n_3106),
.Y(n_3348)
);

OAI21x1_ASAP7_75t_L g3349 ( 
.A1(n_3228),
.A2(n_1578),
.B(n_2234),
.Y(n_3349)
);

INVx2_ASAP7_75t_L g3350 ( 
.A(n_3113),
.Y(n_3350)
);

INVx6_ASAP7_75t_L g3351 ( 
.A(n_3089),
.Y(n_3351)
);

AOI21xp5_ASAP7_75t_L g3352 ( 
.A1(n_3249),
.A2(n_1578),
.B(n_1576),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_3147),
.Y(n_3353)
);

OAI21x1_ASAP7_75t_L g3354 ( 
.A1(n_3142),
.A2(n_3081),
.B(n_3125),
.Y(n_3354)
);

A2O1A1Ixp33_ASAP7_75t_L g3355 ( 
.A1(n_3237),
.A2(n_119),
.B(n_120),
.C(n_122),
.Y(n_3355)
);

NAND3xp33_ASAP7_75t_L g3356 ( 
.A(n_3115),
.B(n_1576),
.C(n_1571),
.Y(n_3356)
);

AOI21xp5_ASAP7_75t_L g3357 ( 
.A1(n_3217),
.A2(n_1576),
.B(n_1571),
.Y(n_3357)
);

AOI21x1_ASAP7_75t_L g3358 ( 
.A1(n_3163),
.A2(n_119),
.B(n_123),
.Y(n_3358)
);

NOR2xp33_ASAP7_75t_L g3359 ( 
.A(n_3068),
.B(n_124),
.Y(n_3359)
);

OAI21x1_ASAP7_75t_L g3360 ( 
.A1(n_3131),
.A2(n_3215),
.B(n_3102),
.Y(n_3360)
);

AND2x4_ASAP7_75t_L g3361 ( 
.A(n_3111),
.B(n_124),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3105),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_3105),
.Y(n_3363)
);

NOR2xp33_ASAP7_75t_L g3364 ( 
.A(n_3114),
.B(n_126),
.Y(n_3364)
);

NOR2xp33_ASAP7_75t_L g3365 ( 
.A(n_3116),
.B(n_126),
.Y(n_3365)
);

A2O1A1Ixp33_ASAP7_75t_L g3366 ( 
.A1(n_3237),
.A2(n_128),
.B(n_129),
.C(n_131),
.Y(n_3366)
);

O2A1O1Ixp33_ASAP7_75t_SL g3367 ( 
.A1(n_3084),
.A2(n_128),
.B(n_131),
.C(n_132),
.Y(n_3367)
);

O2A1O1Ixp33_ASAP7_75t_SL g3368 ( 
.A1(n_3143),
.A2(n_132),
.B(n_133),
.C(n_134),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_SL g3369 ( 
.A(n_3148),
.B(n_1571),
.Y(n_3369)
);

AND2x4_ASAP7_75t_L g3370 ( 
.A(n_3111),
.B(n_133),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_3235),
.B(n_135),
.Y(n_3371)
);

BUFx10_ASAP7_75t_L g3372 ( 
.A(n_3183),
.Y(n_3372)
);

AO32x2_ASAP7_75t_L g3373 ( 
.A1(n_3075),
.A2(n_135),
.A3(n_136),
.B1(n_137),
.B2(n_140),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_3128),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_L g3375 ( 
.A(n_3248),
.B(n_137),
.Y(n_3375)
);

OAI21xp5_ASAP7_75t_L g3376 ( 
.A1(n_3192),
.A2(n_142),
.B(n_143),
.Y(n_3376)
);

AO21x1_ASAP7_75t_L g3377 ( 
.A1(n_3211),
.A2(n_3160),
.B(n_3098),
.Y(n_3377)
);

A2O1A1Ixp33_ASAP7_75t_L g3378 ( 
.A1(n_3103),
.A2(n_142),
.B(n_145),
.C(n_147),
.Y(n_3378)
);

BUFx10_ASAP7_75t_L g3379 ( 
.A(n_3148),
.Y(n_3379)
);

OR2x2_ASAP7_75t_L g3380 ( 
.A(n_3151),
.B(n_145),
.Y(n_3380)
);

OAI22x1_ASAP7_75t_L g3381 ( 
.A1(n_3093),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_3381)
);

AOI22xp33_ASAP7_75t_L g3382 ( 
.A1(n_3133),
.A2(n_3246),
.B1(n_3234),
.B2(n_3103),
.Y(n_3382)
);

BUFx12f_ASAP7_75t_L g3383 ( 
.A(n_3148),
.Y(n_3383)
);

INVx2_ASAP7_75t_L g3384 ( 
.A(n_3166),
.Y(n_3384)
);

OAI22xp5_ASAP7_75t_L g3385 ( 
.A1(n_3227),
.A2(n_2234),
.B1(n_1577),
.B2(n_1576),
.Y(n_3385)
);

NAND2x1p5_ASAP7_75t_L g3386 ( 
.A(n_3124),
.B(n_3144),
.Y(n_3386)
);

OAI21x1_ASAP7_75t_L g3387 ( 
.A1(n_3205),
.A2(n_148),
.B(n_149),
.Y(n_3387)
);

CKINVDCx16_ASAP7_75t_R g3388 ( 
.A(n_3189),
.Y(n_3388)
);

AO31x2_ASAP7_75t_L g3389 ( 
.A1(n_3096),
.A2(n_150),
.A3(n_151),
.B(n_152),
.Y(n_3389)
);

A2O1A1Ixp33_ASAP7_75t_L g3390 ( 
.A1(n_3095),
.A2(n_151),
.B(n_153),
.C(n_155),
.Y(n_3390)
);

A2O1A1Ixp33_ASAP7_75t_L g3391 ( 
.A1(n_3095),
.A2(n_153),
.B(n_156),
.C(n_157),
.Y(n_3391)
);

INVx1_ASAP7_75t_SL g3392 ( 
.A(n_3226),
.Y(n_3392)
);

INVx2_ASAP7_75t_L g3393 ( 
.A(n_3180),
.Y(n_3393)
);

OAI21x1_ASAP7_75t_L g3394 ( 
.A1(n_3119),
.A2(n_156),
.B(n_158),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_3128),
.Y(n_3395)
);

AO31x2_ASAP7_75t_L g3396 ( 
.A1(n_3259),
.A2(n_158),
.A3(n_159),
.B(n_162),
.Y(n_3396)
);

INVx8_ASAP7_75t_L g3397 ( 
.A(n_3239),
.Y(n_3397)
);

OAI22xp5_ASAP7_75t_L g3398 ( 
.A1(n_3092),
.A2(n_1577),
.B1(n_1519),
.B2(n_1511),
.Y(n_3398)
);

BUFx3_ASAP7_75t_L g3399 ( 
.A(n_3167),
.Y(n_3399)
);

OA21x2_ASAP7_75t_L g3400 ( 
.A1(n_3092),
.A2(n_163),
.B(n_164),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_3196),
.B(n_163),
.Y(n_3401)
);

OAI21xp5_ASAP7_75t_L g3402 ( 
.A1(n_3232),
.A2(n_164),
.B(n_166),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_3132),
.Y(n_3403)
);

AOI31xp67_ASAP7_75t_L g3404 ( 
.A1(n_3157),
.A2(n_166),
.A3(n_167),
.B(n_168),
.Y(n_3404)
);

AOI22xp5_ASAP7_75t_L g3405 ( 
.A1(n_3172),
.A2(n_1577),
.B1(n_1519),
.B2(n_1511),
.Y(n_3405)
);

NOR2xp33_ASAP7_75t_L g3406 ( 
.A(n_3129),
.B(n_168),
.Y(n_3406)
);

OAI21x1_ASAP7_75t_SL g3407 ( 
.A1(n_3199),
.A2(n_169),
.B(n_170),
.Y(n_3407)
);

OA21x2_ASAP7_75t_L g3408 ( 
.A1(n_3098),
.A2(n_169),
.B(n_170),
.Y(n_3408)
);

AO31x2_ASAP7_75t_L g3409 ( 
.A1(n_3259),
.A2(n_3172),
.A3(n_3100),
.B(n_3140),
.Y(n_3409)
);

AO31x2_ASAP7_75t_L g3410 ( 
.A1(n_3100),
.A2(n_171),
.A3(n_172),
.B(n_174),
.Y(n_3410)
);

BUFx12f_ASAP7_75t_L g3411 ( 
.A(n_3252),
.Y(n_3411)
);

AO21x1_ASAP7_75t_L g3412 ( 
.A1(n_3132),
.A2(n_171),
.B(n_172),
.Y(n_3412)
);

OAI21x1_ASAP7_75t_L g3413 ( 
.A1(n_3181),
.A2(n_175),
.B(n_176),
.Y(n_3413)
);

AOI21xp5_ASAP7_75t_L g3414 ( 
.A1(n_3174),
.A2(n_1577),
.B(n_1430),
.Y(n_3414)
);

A2O1A1Ixp33_ASAP7_75t_L g3415 ( 
.A1(n_3191),
.A2(n_176),
.B(n_177),
.C(n_180),
.Y(n_3415)
);

AOI21xp5_ASAP7_75t_L g3416 ( 
.A1(n_3258),
.A2(n_1577),
.B(n_1430),
.Y(n_3416)
);

OR2x2_ASAP7_75t_L g3417 ( 
.A(n_3136),
.B(n_177),
.Y(n_3417)
);

BUFx10_ASAP7_75t_L g3418 ( 
.A(n_3195),
.Y(n_3418)
);

NOR2xp33_ASAP7_75t_L g3419 ( 
.A(n_3129),
.B(n_180),
.Y(n_3419)
);

INVx3_ASAP7_75t_L g3420 ( 
.A(n_3190),
.Y(n_3420)
);

BUFx2_ASAP7_75t_L g3421 ( 
.A(n_3127),
.Y(n_3421)
);

INVx2_ASAP7_75t_L g3422 ( 
.A(n_3224),
.Y(n_3422)
);

OAI22x1_ASAP7_75t_L g3423 ( 
.A1(n_3099),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_3403),
.Y(n_3424)
);

OAI21x1_ASAP7_75t_L g3425 ( 
.A1(n_3328),
.A2(n_3154),
.B(n_3133),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3403),
.Y(n_3426)
);

AOI22xp33_ASAP7_75t_L g3427 ( 
.A1(n_3286),
.A2(n_3153),
.B1(n_3191),
.B2(n_3126),
.Y(n_3427)
);

AND2x2_ASAP7_75t_L g3428 ( 
.A(n_3388),
.B(n_3127),
.Y(n_3428)
);

NOR3xp33_ASAP7_75t_SL g3429 ( 
.A(n_3313),
.B(n_3196),
.C(n_3216),
.Y(n_3429)
);

NOR2xp33_ASAP7_75t_L g3430 ( 
.A(n_3392),
.B(n_3209),
.Y(n_3430)
);

OAI21x1_ASAP7_75t_L g3431 ( 
.A1(n_3348),
.A2(n_3149),
.B(n_3135),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_3327),
.Y(n_3432)
);

OAI21xp5_ASAP7_75t_L g3433 ( 
.A1(n_3269),
.A2(n_3230),
.B(n_3165),
.Y(n_3433)
);

INVx2_ASAP7_75t_SL g3434 ( 
.A(n_3397),
.Y(n_3434)
);

CKINVDCx11_ASAP7_75t_R g3435 ( 
.A(n_3372),
.Y(n_3435)
);

AND2x2_ASAP7_75t_SL g3436 ( 
.A(n_3282),
.B(n_3209),
.Y(n_3436)
);

OA21x2_ASAP7_75t_L g3437 ( 
.A1(n_3354),
.A2(n_3136),
.B(n_3152),
.Y(n_3437)
);

AND2x4_ASAP7_75t_L g3438 ( 
.A(n_3331),
.B(n_3216),
.Y(n_3438)
);

NOR2xp33_ASAP7_75t_SL g3439 ( 
.A(n_3265),
.B(n_3198),
.Y(n_3439)
);

INVx6_ASAP7_75t_L g3440 ( 
.A(n_3372),
.Y(n_3440)
);

OAI221xp5_ASAP7_75t_L g3441 ( 
.A1(n_3376),
.A2(n_3230),
.B1(n_3165),
.B2(n_3198),
.C(n_3187),
.Y(n_3441)
);

OAI21x1_ASAP7_75t_L g3442 ( 
.A1(n_3360),
.A2(n_3158),
.B(n_3161),
.Y(n_3442)
);

AOI22xp33_ASAP7_75t_SL g3443 ( 
.A1(n_3400),
.A2(n_3153),
.B1(n_3209),
.B2(n_3127),
.Y(n_3443)
);

NOR2xp33_ASAP7_75t_L g3444 ( 
.A(n_3333),
.B(n_3127),
.Y(n_3444)
);

OA21x2_ASAP7_75t_L g3445 ( 
.A1(n_3272),
.A2(n_3194),
.B(n_3178),
.Y(n_3445)
);

CKINVDCx14_ASAP7_75t_R g3446 ( 
.A(n_3316),
.Y(n_3446)
);

AND2x2_ASAP7_75t_L g3447 ( 
.A(n_3420),
.B(n_3127),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_L g3448 ( 
.A(n_3327),
.B(n_3213),
.Y(n_3448)
);

CKINVDCx20_ASAP7_75t_R g3449 ( 
.A(n_3298),
.Y(n_3449)
);

AOI22xp33_ASAP7_75t_L g3450 ( 
.A1(n_3382),
.A2(n_3253),
.B1(n_3187),
.B2(n_3242),
.Y(n_3450)
);

INVx8_ASAP7_75t_L g3451 ( 
.A(n_3361),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_3362),
.Y(n_3452)
);

OAI21x1_ASAP7_75t_L g3453 ( 
.A1(n_3270),
.A2(n_3197),
.B(n_3238),
.Y(n_3453)
);

OA21x2_ASAP7_75t_L g3454 ( 
.A1(n_3377),
.A2(n_3238),
.B(n_3197),
.Y(n_3454)
);

AND2x4_ASAP7_75t_L g3455 ( 
.A(n_3420),
.B(n_3195),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3363),
.Y(n_3456)
);

AOI22xp33_ASAP7_75t_L g3457 ( 
.A1(n_3347),
.A2(n_3253),
.B1(n_3245),
.B2(n_3244),
.Y(n_3457)
);

INVx2_ASAP7_75t_L g3458 ( 
.A(n_3344),
.Y(n_3458)
);

OAI221xp5_ASAP7_75t_L g3459 ( 
.A1(n_3278),
.A2(n_3222),
.B1(n_3233),
.B2(n_3179),
.C(n_3223),
.Y(n_3459)
);

OAI22xp5_ASAP7_75t_L g3460 ( 
.A1(n_3378),
.A2(n_3233),
.B1(n_3179),
.B2(n_3245),
.Y(n_3460)
);

AND2x4_ASAP7_75t_L g3461 ( 
.A(n_3421),
.B(n_3176),
.Y(n_3461)
);

AND2x4_ASAP7_75t_L g3462 ( 
.A(n_3289),
.B(n_3168),
.Y(n_3462)
);

OAI21xp5_ASAP7_75t_L g3463 ( 
.A1(n_3415),
.A2(n_3222),
.B(n_3067),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_L g3464 ( 
.A(n_3374),
.B(n_3241),
.Y(n_3464)
);

AOI21xp5_ASAP7_75t_L g3465 ( 
.A1(n_3345),
.A2(n_3218),
.B(n_3184),
.Y(n_3465)
);

OA21x2_ASAP7_75t_L g3466 ( 
.A1(n_3334),
.A2(n_3219),
.B(n_3200),
.Y(n_3466)
);

INVx3_ASAP7_75t_SL g3467 ( 
.A(n_3361),
.Y(n_3467)
);

AOI221xp5_ASAP7_75t_L g3468 ( 
.A1(n_3308),
.A2(n_181),
.B1(n_182),
.B2(n_186),
.C(n_187),
.Y(n_3468)
);

AO21x2_ASAP7_75t_L g3469 ( 
.A1(n_3310),
.A2(n_3204),
.B(n_3173),
.Y(n_3469)
);

BUFx2_ASAP7_75t_L g3470 ( 
.A(n_3305),
.Y(n_3470)
);

INVx2_ASAP7_75t_L g3471 ( 
.A(n_3395),
.Y(n_3471)
);

INVx2_ASAP7_75t_L g3472 ( 
.A(n_3353),
.Y(n_3472)
);

OAI21x1_ASAP7_75t_L g3473 ( 
.A1(n_3319),
.A2(n_3177),
.B(n_3164),
.Y(n_3473)
);

O2A1O1Ixp33_ASAP7_75t_SL g3474 ( 
.A1(n_3359),
.A2(n_186),
.B(n_187),
.C(n_190),
.Y(n_3474)
);

OAI21x1_ASAP7_75t_L g3475 ( 
.A1(n_3268),
.A2(n_3212),
.B(n_3188),
.Y(n_3475)
);

AO21x2_ASAP7_75t_L g3476 ( 
.A1(n_3312),
.A2(n_3170),
.B(n_3186),
.Y(n_3476)
);

AO21x2_ASAP7_75t_L g3477 ( 
.A1(n_3342),
.A2(n_3170),
.B(n_3241),
.Y(n_3477)
);

OA21x2_ASAP7_75t_L g3478 ( 
.A1(n_3297),
.A2(n_3150),
.B(n_3168),
.Y(n_3478)
);

OR2x6_ASAP7_75t_L g3479 ( 
.A(n_3341),
.B(n_3283),
.Y(n_3479)
);

AO21x2_ASAP7_75t_L g3480 ( 
.A1(n_3291),
.A2(n_3241),
.B(n_3207),
.Y(n_3480)
);

NAND2x1p5_ASAP7_75t_L g3481 ( 
.A(n_3330),
.B(n_3168),
.Y(n_3481)
);

O2A1O1Ixp33_ASAP7_75t_L g3482 ( 
.A1(n_3307),
.A2(n_192),
.B(n_193),
.C(n_194),
.Y(n_3482)
);

NOR2xp33_ASAP7_75t_L g3483 ( 
.A(n_3322),
.B(n_192),
.Y(n_3483)
);

OAI221xp5_ASAP7_75t_L g3484 ( 
.A1(n_3355),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.C(n_197),
.Y(n_3484)
);

INVxp67_ASAP7_75t_L g3485 ( 
.A(n_3300),
.Y(n_3485)
);

OAI22xp5_ASAP7_75t_L g3486 ( 
.A1(n_3390),
.A2(n_198),
.B1(n_199),
.B2(n_201),
.Y(n_3486)
);

OAI21x1_ASAP7_75t_L g3487 ( 
.A1(n_3416),
.A2(n_3274),
.B(n_3290),
.Y(n_3487)
);

OAI21xp33_ASAP7_75t_L g3488 ( 
.A1(n_3391),
.A2(n_198),
.B(n_199),
.Y(n_3488)
);

OAI21x1_ASAP7_75t_L g3489 ( 
.A1(n_3296),
.A2(n_3150),
.B(n_3207),
.Y(n_3489)
);

INVx2_ASAP7_75t_L g3490 ( 
.A(n_3311),
.Y(n_3490)
);

A2O1A1Ixp33_ASAP7_75t_L g3491 ( 
.A1(n_3340),
.A2(n_201),
.B(n_203),
.C(n_205),
.Y(n_3491)
);

AOI21xp33_ASAP7_75t_L g3492 ( 
.A1(n_3412),
.A2(n_203),
.B(n_206),
.Y(n_3492)
);

NAND2x1p5_ASAP7_75t_L g3493 ( 
.A(n_3330),
.B(n_3206),
.Y(n_3493)
);

OA21x2_ASAP7_75t_L g3494 ( 
.A1(n_3279),
.A2(n_3207),
.B(n_3206),
.Y(n_3494)
);

INVx2_ASAP7_75t_L g3495 ( 
.A(n_3350),
.Y(n_3495)
);

INVx1_ASAP7_75t_L g3496 ( 
.A(n_3314),
.Y(n_3496)
);

NAND2xp33_ASAP7_75t_SL g3497 ( 
.A(n_3276),
.B(n_207),
.Y(n_3497)
);

AND2x4_ASAP7_75t_L g3498 ( 
.A(n_3294),
.B(n_3206),
.Y(n_3498)
);

INVx1_ASAP7_75t_L g3499 ( 
.A(n_3325),
.Y(n_3499)
);

OA21x2_ASAP7_75t_L g3500 ( 
.A1(n_3284),
.A2(n_3401),
.B(n_3326),
.Y(n_3500)
);

NAND2x1p5_ASAP7_75t_L g3501 ( 
.A(n_3330),
.B(n_208),
.Y(n_3501)
);

OR2x2_ASAP7_75t_L g3502 ( 
.A(n_3399),
.B(n_208),
.Y(n_3502)
);

NAND2x1p5_ASAP7_75t_L g3503 ( 
.A(n_3339),
.B(n_209),
.Y(n_3503)
);

NOR2xp33_ASAP7_75t_L g3504 ( 
.A(n_3277),
.B(n_211),
.Y(n_3504)
);

AOI21xp5_ASAP7_75t_L g3505 ( 
.A1(n_3352),
.A2(n_1428),
.B(n_1430),
.Y(n_3505)
);

INVx3_ASAP7_75t_L g3506 ( 
.A(n_3418),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_3294),
.B(n_212),
.Y(n_3507)
);

AOI21xp5_ASAP7_75t_L g3508 ( 
.A1(n_3357),
.A2(n_1428),
.B(n_1430),
.Y(n_3508)
);

NOR2xp33_ASAP7_75t_L g3509 ( 
.A(n_3364),
.B(n_3332),
.Y(n_3509)
);

AO21x2_ASAP7_75t_L g3510 ( 
.A1(n_3295),
.A2(n_212),
.B(n_214),
.Y(n_3510)
);

BUFx8_ASAP7_75t_SL g3511 ( 
.A(n_3411),
.Y(n_3511)
);

OAI21x1_ASAP7_75t_L g3512 ( 
.A1(n_3304),
.A2(n_214),
.B(n_215),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_3417),
.Y(n_3513)
);

OAI222xp33_ASAP7_75t_L g3514 ( 
.A1(n_3380),
.A2(n_3282),
.B1(n_3346),
.B2(n_3292),
.C1(n_3306),
.C2(n_3384),
.Y(n_3514)
);

INVx4_ASAP7_75t_L g3515 ( 
.A(n_3383),
.Y(n_3515)
);

OR2x2_ASAP7_75t_L g3516 ( 
.A(n_3294),
.B(n_216),
.Y(n_3516)
);

NAND2x1p5_ASAP7_75t_L g3517 ( 
.A(n_3339),
.B(n_216),
.Y(n_3517)
);

INVx2_ASAP7_75t_L g3518 ( 
.A(n_3393),
.Y(n_3518)
);

OA21x2_ASAP7_75t_L g3519 ( 
.A1(n_3371),
.A2(n_3375),
.B(n_3320),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_3422),
.Y(n_3520)
);

NAND2x1p5_ASAP7_75t_L g3521 ( 
.A(n_3339),
.B(n_217),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_3409),
.B(n_217),
.Y(n_3522)
);

AOI22xp33_ASAP7_75t_L g3523 ( 
.A1(n_3315),
.A2(n_1519),
.B1(n_1466),
.B2(n_1463),
.Y(n_3523)
);

AOI22xp5_ASAP7_75t_L g3524 ( 
.A1(n_3285),
.A2(n_3324),
.B1(n_3366),
.B2(n_3423),
.Y(n_3524)
);

OAI211xp5_ASAP7_75t_L g3525 ( 
.A1(n_3368),
.A2(n_218),
.B(n_219),
.C(n_220),
.Y(n_3525)
);

OA21x2_ASAP7_75t_L g3526 ( 
.A1(n_3338),
.A2(n_218),
.B(n_219),
.Y(n_3526)
);

INVx1_ASAP7_75t_L g3527 ( 
.A(n_3410),
.Y(n_3527)
);

INVx3_ASAP7_75t_L g3528 ( 
.A(n_3418),
.Y(n_3528)
);

OAI21x1_ASAP7_75t_L g3529 ( 
.A1(n_3275),
.A2(n_220),
.B(n_221),
.Y(n_3529)
);

AO21x2_ASAP7_75t_L g3530 ( 
.A1(n_3266),
.A2(n_221),
.B(n_222),
.Y(n_3530)
);

O2A1O1Ixp33_ASAP7_75t_SL g3531 ( 
.A1(n_3281),
.A2(n_224),
.B(n_226),
.C(n_227),
.Y(n_3531)
);

OAI21x1_ASAP7_75t_SL g3532 ( 
.A1(n_3407),
.A2(n_224),
.B(n_228),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3410),
.Y(n_3533)
);

OAI21x1_ASAP7_75t_L g3534 ( 
.A1(n_3400),
.A2(n_229),
.B(n_230),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3410),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_L g3536 ( 
.A(n_3409),
.B(n_232),
.Y(n_3536)
);

AOI221xp5_ASAP7_75t_L g3537 ( 
.A1(n_3309),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.C(n_235),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_3408),
.Y(n_3538)
);

BUFx8_ASAP7_75t_L g3539 ( 
.A(n_3370),
.Y(n_3539)
);

OAI21x1_ASAP7_75t_L g3540 ( 
.A1(n_3287),
.A2(n_234),
.B(n_236),
.Y(n_3540)
);

OR2x2_ASAP7_75t_L g3541 ( 
.A(n_3409),
.B(n_236),
.Y(n_3541)
);

CKINVDCx5p33_ASAP7_75t_R g3542 ( 
.A(n_3351),
.Y(n_3542)
);

OAI22xp33_ASAP7_75t_L g3543 ( 
.A1(n_3381),
.A2(n_238),
.B1(n_241),
.B2(n_242),
.Y(n_3543)
);

OR2x2_ASAP7_75t_L g3544 ( 
.A(n_3305),
.B(n_241),
.Y(n_3544)
);

INVx2_ASAP7_75t_L g3545 ( 
.A(n_3293),
.Y(n_3545)
);

AOI22xp33_ASAP7_75t_L g3546 ( 
.A1(n_3433),
.A2(n_3385),
.B1(n_3402),
.B2(n_3280),
.Y(n_3546)
);

INVx6_ASAP7_75t_L g3547 ( 
.A(n_3539),
.Y(n_3547)
);

OR2x6_ASAP7_75t_L g3548 ( 
.A(n_3433),
.B(n_3370),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_3538),
.B(n_3396),
.Y(n_3549)
);

OA21x2_ASAP7_75t_L g3550 ( 
.A1(n_3458),
.A2(n_3323),
.B(n_3414),
.Y(n_3550)
);

OAI21xp5_ASAP7_75t_L g3551 ( 
.A1(n_3524),
.A2(n_3404),
.B(n_3365),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3452),
.Y(n_3552)
);

INVx2_ASAP7_75t_L g3553 ( 
.A(n_3516),
.Y(n_3553)
);

AO31x2_ASAP7_75t_L g3554 ( 
.A1(n_3522),
.A2(n_3419),
.A3(n_3406),
.B(n_3398),
.Y(n_3554)
);

INVx1_ASAP7_75t_L g3555 ( 
.A(n_3456),
.Y(n_3555)
);

AO21x2_ASAP7_75t_L g3556 ( 
.A1(n_3536),
.A2(n_3358),
.B(n_3356),
.Y(n_3556)
);

BUFx6f_ASAP7_75t_L g3557 ( 
.A(n_3435),
.Y(n_3557)
);

CKINVDCx20_ASAP7_75t_R g3558 ( 
.A(n_3449),
.Y(n_3558)
);

AO21x2_ASAP7_75t_L g3559 ( 
.A1(n_3536),
.A2(n_3394),
.B(n_3413),
.Y(n_3559)
);

INVx2_ASAP7_75t_L g3560 ( 
.A(n_3437),
.Y(n_3560)
);

CKINVDCx11_ASAP7_75t_R g3561 ( 
.A(n_3467),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_L g3562 ( 
.A(n_3432),
.B(n_3396),
.Y(n_3562)
);

OAI21x1_ASAP7_75t_SL g3563 ( 
.A1(n_3434),
.A2(n_3373),
.B(n_3303),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_3424),
.B(n_3396),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3448),
.Y(n_3565)
);

BUFx10_ASAP7_75t_L g3566 ( 
.A(n_3483),
.Y(n_3566)
);

INVx2_ASAP7_75t_L g3567 ( 
.A(n_3437),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_L g3568 ( 
.A(n_3426),
.B(n_3500),
.Y(n_3568)
);

INVx2_ASAP7_75t_L g3569 ( 
.A(n_3471),
.Y(n_3569)
);

INVx3_ASAP7_75t_L g3570 ( 
.A(n_3455),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_3500),
.B(n_3389),
.Y(n_3571)
);

INVx3_ASAP7_75t_L g3572 ( 
.A(n_3455),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3448),
.B(n_3389),
.Y(n_3573)
);

OAI21x1_ASAP7_75t_L g3574 ( 
.A1(n_3431),
.A2(n_3386),
.B(n_3271),
.Y(n_3574)
);

INVx2_ASAP7_75t_L g3575 ( 
.A(n_3472),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_SL g3576 ( 
.A(n_3436),
.B(n_3321),
.Y(n_3576)
);

AND2x4_ASAP7_75t_L g3577 ( 
.A(n_3428),
.B(n_3321),
.Y(n_3577)
);

OR2x6_ASAP7_75t_L g3578 ( 
.A(n_3479),
.B(n_3351),
.Y(n_3578)
);

AOI21xp5_ASAP7_75t_L g3579 ( 
.A1(n_3463),
.A2(n_3367),
.B(n_3369),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3429),
.B(n_3389),
.Y(n_3580)
);

OAI21xp5_ASAP7_75t_L g3581 ( 
.A1(n_3524),
.A2(n_3387),
.B(n_3373),
.Y(n_3581)
);

AO31x2_ASAP7_75t_L g3582 ( 
.A1(n_3507),
.A2(n_3335),
.A3(n_3288),
.B(n_3373),
.Y(n_3582)
);

OAI21x1_ASAP7_75t_L g3583 ( 
.A1(n_3507),
.A2(n_3336),
.B(n_3337),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_L g3584 ( 
.A(n_3541),
.B(n_3343),
.Y(n_3584)
);

AOI21xp5_ASAP7_75t_L g3585 ( 
.A1(n_3463),
.A2(n_3317),
.B(n_3267),
.Y(n_3585)
);

INVx6_ASAP7_75t_L g3586 ( 
.A(n_3451),
.Y(n_3586)
);

OR2x2_ASAP7_75t_L g3587 ( 
.A(n_3485),
.B(n_3321),
.Y(n_3587)
);

OAI22xp5_ASAP7_75t_L g3588 ( 
.A1(n_3441),
.A2(n_3405),
.B1(n_3317),
.B2(n_3318),
.Y(n_3588)
);

AO21x2_ASAP7_75t_L g3589 ( 
.A1(n_3527),
.A2(n_3349),
.B(n_3302),
.Y(n_3589)
);

OR2x2_ASAP7_75t_L g3590 ( 
.A(n_3513),
.B(n_3343),
.Y(n_3590)
);

AO31x2_ASAP7_75t_L g3591 ( 
.A1(n_3533),
.A2(n_3273),
.A3(n_3299),
.B(n_3293),
.Y(n_3591)
);

AOI21xp5_ASAP7_75t_L g3592 ( 
.A1(n_3479),
.A2(n_3329),
.B(n_3273),
.Y(n_3592)
);

OAI21x1_ASAP7_75t_L g3593 ( 
.A1(n_3425),
.A2(n_3293),
.B(n_3301),
.Y(n_3593)
);

OA21x2_ASAP7_75t_L g3594 ( 
.A1(n_3464),
.A2(n_3301),
.B(n_3379),
.Y(n_3594)
);

AOI21xp5_ASAP7_75t_L g3595 ( 
.A1(n_3479),
.A2(n_3379),
.B(n_3301),
.Y(n_3595)
);

OAI21x1_ASAP7_75t_SL g3596 ( 
.A1(n_3515),
.A2(n_242),
.B(n_243),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_L g3597 ( 
.A(n_3496),
.B(n_243),
.Y(n_3597)
);

CKINVDCx5p33_ASAP7_75t_R g3598 ( 
.A(n_3511),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_3499),
.B(n_245),
.Y(n_3599)
);

INVx2_ASAP7_75t_L g3600 ( 
.A(n_3498),
.Y(n_3600)
);

OA21x2_ASAP7_75t_L g3601 ( 
.A1(n_3464),
.A2(n_254),
.B(n_256),
.Y(n_3601)
);

INVx2_ASAP7_75t_L g3602 ( 
.A(n_3498),
.Y(n_3602)
);

HB1xp67_ASAP7_75t_L g3603 ( 
.A(n_3454),
.Y(n_3603)
);

INVx2_ASAP7_75t_L g3604 ( 
.A(n_3454),
.Y(n_3604)
);

OR2x2_ASAP7_75t_L g3605 ( 
.A(n_3438),
.B(n_256),
.Y(n_3605)
);

CKINVDCx8_ASAP7_75t_R g3606 ( 
.A(n_3542),
.Y(n_3606)
);

AND2x4_ASAP7_75t_L g3607 ( 
.A(n_3470),
.B(n_3438),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_3535),
.B(n_3519),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_L g3609 ( 
.A(n_3519),
.B(n_257),
.Y(n_3609)
);

AOI21x1_ASAP7_75t_L g3610 ( 
.A1(n_3462),
.A2(n_259),
.B(n_261),
.Y(n_3610)
);

AOI21xp5_ASAP7_75t_L g3611 ( 
.A1(n_3441),
.A2(n_1466),
.B(n_1463),
.Y(n_3611)
);

INVx2_ASAP7_75t_L g3612 ( 
.A(n_3490),
.Y(n_3612)
);

BUFx2_ASAP7_75t_L g3613 ( 
.A(n_3446),
.Y(n_3613)
);

INVx2_ASAP7_75t_L g3614 ( 
.A(n_3495),
.Y(n_3614)
);

HB1xp67_ASAP7_75t_L g3615 ( 
.A(n_3526),
.Y(n_3615)
);

NAND2x1p5_ASAP7_75t_L g3616 ( 
.A(n_3506),
.B(n_1428),
.Y(n_3616)
);

INVx2_ASAP7_75t_L g3617 ( 
.A(n_3518),
.Y(n_3617)
);

AO31x2_ASAP7_75t_L g3618 ( 
.A1(n_3509),
.A2(n_263),
.A3(n_266),
.B(n_279),
.Y(n_3618)
);

INVx2_ASAP7_75t_L g3619 ( 
.A(n_3462),
.Y(n_3619)
);

INVx2_ASAP7_75t_SL g3620 ( 
.A(n_3440),
.Y(n_3620)
);

AOI21xp5_ASAP7_75t_SL g3621 ( 
.A1(n_3501),
.A2(n_280),
.B(n_284),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_L g3622 ( 
.A(n_3476),
.B(n_285),
.Y(n_3622)
);

OAI21x1_ASAP7_75t_L g3623 ( 
.A1(n_3481),
.A2(n_3493),
.B(n_3489),
.Y(n_3623)
);

AND2x4_ASAP7_75t_L g3624 ( 
.A(n_3506),
.B(n_3528),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_L g3625 ( 
.A(n_3476),
.B(n_287),
.Y(n_3625)
);

INVx1_ASAP7_75t_L g3626 ( 
.A(n_3520),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_3502),
.Y(n_3627)
);

INVx2_ASAP7_75t_SL g3628 ( 
.A(n_3440),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_3534),
.Y(n_3629)
);

AND2x4_ASAP7_75t_L g3630 ( 
.A(n_3528),
.B(n_292),
.Y(n_3630)
);

OA21x2_ASAP7_75t_L g3631 ( 
.A1(n_3453),
.A2(n_294),
.B(n_295),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3445),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3445),
.Y(n_3633)
);

AND2x2_ASAP7_75t_L g3634 ( 
.A(n_3444),
.B(n_296),
.Y(n_3634)
);

OA21x2_ASAP7_75t_L g3635 ( 
.A1(n_3442),
.A2(n_297),
.B(n_298),
.Y(n_3635)
);

HB1xp67_ASAP7_75t_L g3636 ( 
.A(n_3469),
.Y(n_3636)
);

OAI21xp5_ASAP7_75t_L g3637 ( 
.A1(n_3488),
.A2(n_302),
.B(n_306),
.Y(n_3637)
);

INVx1_ASAP7_75t_L g3638 ( 
.A(n_3544),
.Y(n_3638)
);

AOI21xp5_ASAP7_75t_L g3639 ( 
.A1(n_3439),
.A2(n_1466),
.B(n_1463),
.Y(n_3639)
);

AO21x2_ASAP7_75t_L g3640 ( 
.A1(n_3492),
.A2(n_309),
.B(n_312),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3478),
.Y(n_3641)
);

NAND2x1p5_ASAP7_75t_L g3642 ( 
.A(n_3515),
.B(n_1463),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3480),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3480),
.Y(n_3644)
);

OR2x6_ASAP7_75t_L g3645 ( 
.A(n_3451),
.B(n_1466),
.Y(n_3645)
);

INVx2_ASAP7_75t_L g3646 ( 
.A(n_3466),
.Y(n_3646)
);

INVx1_ASAP7_75t_L g3647 ( 
.A(n_3466),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3494),
.Y(n_3648)
);

NOR3xp33_ASAP7_75t_L g3649 ( 
.A(n_3484),
.B(n_316),
.C(n_317),
.Y(n_3649)
);

AO21x2_ASAP7_75t_L g3650 ( 
.A1(n_3543),
.A2(n_3545),
.B(n_3477),
.Y(n_3650)
);

INVx2_ASAP7_75t_L g3651 ( 
.A(n_3461),
.Y(n_3651)
);

OR2x2_ASAP7_75t_L g3652 ( 
.A(n_3450),
.B(n_319),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_L g3653 ( 
.A(n_3615),
.B(n_3457),
.Y(n_3653)
);

AOI22xp33_ASAP7_75t_SL g3654 ( 
.A1(n_3581),
.A2(n_3439),
.B1(n_3459),
.B2(n_3525),
.Y(n_3654)
);

AOI22xp33_ASAP7_75t_L g3655 ( 
.A1(n_3584),
.A2(n_3427),
.B1(n_3443),
.B2(n_3530),
.Y(n_3655)
);

AOI22xp5_ASAP7_75t_L g3656 ( 
.A1(n_3649),
.A2(n_3497),
.B1(n_3530),
.B2(n_3486),
.Y(n_3656)
);

AOI22xp33_ASAP7_75t_L g3657 ( 
.A1(n_3584),
.A2(n_3484),
.B1(n_3468),
.B2(n_3486),
.Y(n_3657)
);

AOI22xp33_ASAP7_75t_L g3658 ( 
.A1(n_3649),
.A2(n_3468),
.B1(n_3477),
.B2(n_3494),
.Y(n_3658)
);

AND2x2_ASAP7_75t_L g3659 ( 
.A(n_3613),
.B(n_3447),
.Y(n_3659)
);

INVx2_ASAP7_75t_L g3660 ( 
.A(n_3548),
.Y(n_3660)
);

CKINVDCx6p67_ASAP7_75t_R g3661 ( 
.A(n_3557),
.Y(n_3661)
);

AOI22xp33_ASAP7_75t_SL g3662 ( 
.A1(n_3581),
.A2(n_3504),
.B1(n_3451),
.B2(n_3460),
.Y(n_3662)
);

OAI22xp33_ASAP7_75t_L g3663 ( 
.A1(n_3551),
.A2(n_3460),
.B1(n_3517),
.B2(n_3503),
.Y(n_3663)
);

AOI22xp33_ASAP7_75t_L g3664 ( 
.A1(n_3553),
.A2(n_3537),
.B1(n_3532),
.B2(n_3510),
.Y(n_3664)
);

BUFx4f_ASAP7_75t_SL g3665 ( 
.A(n_3558),
.Y(n_3665)
);

INVx2_ASAP7_75t_L g3666 ( 
.A(n_3587),
.Y(n_3666)
);

AOI22xp33_ASAP7_75t_L g3667 ( 
.A1(n_3551),
.A2(n_3537),
.B1(n_3510),
.B2(n_3521),
.Y(n_3667)
);

AO22x1_ASAP7_75t_L g3668 ( 
.A1(n_3603),
.A2(n_3430),
.B1(n_3461),
.B2(n_3514),
.Y(n_3668)
);

CKINVDCx20_ASAP7_75t_R g3669 ( 
.A(n_3561),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_L g3670 ( 
.A(n_3609),
.B(n_3474),
.Y(n_3670)
);

AOI22xp33_ASAP7_75t_SL g3671 ( 
.A1(n_3563),
.A2(n_3650),
.B1(n_3604),
.B2(n_3580),
.Y(n_3671)
);

AOI22xp33_ASAP7_75t_L g3672 ( 
.A1(n_3650),
.A2(n_3465),
.B1(n_3523),
.B2(n_3512),
.Y(n_3672)
);

OAI21xp5_ASAP7_75t_SL g3673 ( 
.A1(n_3579),
.A2(n_3580),
.B(n_3546),
.Y(n_3673)
);

AND2x2_ASAP7_75t_L g3674 ( 
.A(n_3607),
.B(n_3473),
.Y(n_3674)
);

AOI22xp33_ASAP7_75t_L g3675 ( 
.A1(n_3637),
.A2(n_3465),
.B1(n_3505),
.B2(n_3540),
.Y(n_3675)
);

AOI22xp33_ASAP7_75t_SL g3676 ( 
.A1(n_3571),
.A2(n_3531),
.B1(n_3505),
.B2(n_3482),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_L g3677 ( 
.A(n_3601),
.B(n_3491),
.Y(n_3677)
);

NAND2xp5_ASAP7_75t_L g3678 ( 
.A(n_3601),
.B(n_3529),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3552),
.Y(n_3679)
);

NAND2xp5_ASAP7_75t_L g3680 ( 
.A(n_3629),
.B(n_3565),
.Y(n_3680)
);

CKINVDCx5p33_ASAP7_75t_R g3681 ( 
.A(n_3598),
.Y(n_3681)
);

AND2x4_ASAP7_75t_L g3682 ( 
.A(n_3578),
.B(n_3487),
.Y(n_3682)
);

AOI222xp33_ASAP7_75t_L g3683 ( 
.A1(n_3549),
.A2(n_3475),
.B1(n_3508),
.B2(n_326),
.C1(n_328),
.C2(n_329),
.Y(n_3683)
);

BUFx4f_ASAP7_75t_L g3684 ( 
.A(n_3547),
.Y(n_3684)
);

OAI222xp33_ASAP7_75t_L g3685 ( 
.A1(n_3585),
.A2(n_320),
.B1(n_325),
.B2(n_332),
.C1(n_333),
.C2(n_340),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3555),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_3590),
.Y(n_3687)
);

INVx1_ASAP7_75t_L g3688 ( 
.A(n_3597),
.Y(n_3688)
);

INVx3_ASAP7_75t_L g3689 ( 
.A(n_3557),
.Y(n_3689)
);

INVx3_ASAP7_75t_L g3690 ( 
.A(n_3557),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_3597),
.Y(n_3691)
);

CKINVDCx14_ASAP7_75t_R g3692 ( 
.A(n_3547),
.Y(n_3692)
);

BUFx3_ASAP7_75t_L g3693 ( 
.A(n_3606),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_L g3694 ( 
.A(n_3554),
.B(n_349),
.Y(n_3694)
);

OAI22xp5_ASAP7_75t_L g3695 ( 
.A1(n_3586),
.A2(n_1452),
.B1(n_357),
.B2(n_365),
.Y(n_3695)
);

AND2x2_ASAP7_75t_L g3696 ( 
.A(n_3570),
.B(n_369),
.Y(n_3696)
);

AOI22xp33_ASAP7_75t_L g3697 ( 
.A1(n_3556),
.A2(n_388),
.B1(n_389),
.B2(n_390),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_3599),
.Y(n_3698)
);

OAI222xp33_ASAP7_75t_L g3699 ( 
.A1(n_3585),
.A2(n_401),
.B1(n_402),
.B2(n_406),
.C1(n_407),
.C2(n_410),
.Y(n_3699)
);

OAI22xp33_ASAP7_75t_L g3700 ( 
.A1(n_3639),
.A2(n_418),
.B1(n_420),
.B2(n_421),
.Y(n_3700)
);

CKINVDCx20_ASAP7_75t_R g3701 ( 
.A(n_3566),
.Y(n_3701)
);

INVx2_ASAP7_75t_SL g3702 ( 
.A(n_3566),
.Y(n_3702)
);

AOI22xp33_ASAP7_75t_L g3703 ( 
.A1(n_3556),
.A2(n_425),
.B1(n_427),
.B2(n_428),
.Y(n_3703)
);

OAI22xp5_ASAP7_75t_L g3704 ( 
.A1(n_3645),
.A2(n_3605),
.B1(n_3608),
.B2(n_3620),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3599),
.Y(n_3705)
);

OAI22xp5_ASAP7_75t_L g3706 ( 
.A1(n_3645),
.A2(n_3628),
.B1(n_3622),
.B2(n_3625),
.Y(n_3706)
);

AOI22xp5_ASAP7_75t_L g3707 ( 
.A1(n_3640),
.A2(n_3627),
.B1(n_3559),
.B2(n_3631),
.Y(n_3707)
);

AOI222xp33_ASAP7_75t_L g3708 ( 
.A1(n_3571),
.A2(n_3564),
.B1(n_3562),
.B2(n_3573),
.C1(n_3622),
.C2(n_3625),
.Y(n_3708)
);

AND2x2_ASAP7_75t_L g3709 ( 
.A(n_3572),
.B(n_3624),
.Y(n_3709)
);

AOI22xp33_ASAP7_75t_L g3710 ( 
.A1(n_3640),
.A2(n_3559),
.B1(n_3652),
.B2(n_3639),
.Y(n_3710)
);

NOR2xp33_ASAP7_75t_L g3711 ( 
.A(n_3638),
.B(n_3572),
.Y(n_3711)
);

BUFx3_ASAP7_75t_L g3712 ( 
.A(n_3596),
.Y(n_3712)
);

AND2x2_ASAP7_75t_L g3713 ( 
.A(n_3624),
.B(n_3577),
.Y(n_3713)
);

OAI22xp5_ASAP7_75t_L g3714 ( 
.A1(n_3611),
.A2(n_3573),
.B1(n_3568),
.B2(n_3562),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_3554),
.B(n_3568),
.Y(n_3715)
);

OAI21xp5_ASAP7_75t_SL g3716 ( 
.A1(n_3611),
.A2(n_3642),
.B(n_3588),
.Y(n_3716)
);

AOI22xp33_ASAP7_75t_SL g3717 ( 
.A1(n_3631),
.A2(n_3633),
.B1(n_3632),
.B2(n_3560),
.Y(n_3717)
);

OAI21xp5_ASAP7_75t_SL g3718 ( 
.A1(n_3642),
.A2(n_3588),
.B(n_3651),
.Y(n_3718)
);

NAND2xp5_ASAP7_75t_L g3719 ( 
.A(n_3554),
.B(n_3626),
.Y(n_3719)
);

AOI22xp5_ASAP7_75t_L g3720 ( 
.A1(n_3635),
.A2(n_3564),
.B1(n_3569),
.B2(n_3575),
.Y(n_3720)
);

OAI222xp33_ASAP7_75t_L g3721 ( 
.A1(n_3641),
.A2(n_3567),
.B1(n_3648),
.B2(n_3647),
.C1(n_3643),
.C2(n_3644),
.Y(n_3721)
);

INVx1_ASAP7_75t_SL g3722 ( 
.A(n_3630),
.Y(n_3722)
);

INVx2_ASAP7_75t_SL g3723 ( 
.A(n_3577),
.Y(n_3723)
);

AOI22xp33_ASAP7_75t_L g3724 ( 
.A1(n_3635),
.A2(n_3600),
.B1(n_3602),
.B2(n_3617),
.Y(n_3724)
);

BUFx4f_ASAP7_75t_SL g3725 ( 
.A(n_3634),
.Y(n_3725)
);

OR2x2_ASAP7_75t_L g3726 ( 
.A(n_3582),
.B(n_3619),
.Y(n_3726)
);

HB1xp67_ASAP7_75t_L g3727 ( 
.A(n_3636),
.Y(n_3727)
);

CKINVDCx5p33_ASAP7_75t_R g3728 ( 
.A(n_3621),
.Y(n_3728)
);

AOI22xp33_ASAP7_75t_L g3729 ( 
.A1(n_3612),
.A2(n_3614),
.B1(n_3646),
.B2(n_3550),
.Y(n_3729)
);

AOI22xp33_ASAP7_75t_SL g3730 ( 
.A1(n_3550),
.A2(n_3582),
.B1(n_3594),
.B2(n_3623),
.Y(n_3730)
);

AND2x2_ASAP7_75t_L g3731 ( 
.A(n_3616),
.B(n_3576),
.Y(n_3731)
);

OAI22xp33_ASAP7_75t_L g3732 ( 
.A1(n_3595),
.A2(n_3592),
.B1(n_3610),
.B2(n_3582),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_3583),
.Y(n_3733)
);

AOI22xp33_ASAP7_75t_L g3734 ( 
.A1(n_3589),
.A2(n_3592),
.B1(n_3593),
.B2(n_3594),
.Y(n_3734)
);

BUFx3_ASAP7_75t_L g3735 ( 
.A(n_3616),
.Y(n_3735)
);

INVx3_ASAP7_75t_SL g3736 ( 
.A(n_3618),
.Y(n_3736)
);

OAI222xp33_ASAP7_75t_L g3737 ( 
.A1(n_3618),
.A2(n_3574),
.B1(n_3591),
.B2(n_3615),
.C1(n_3584),
.C2(n_3548),
.Y(n_3737)
);

AOI22xp33_ASAP7_75t_L g3738 ( 
.A1(n_3618),
.A2(n_3169),
.B1(n_3584),
.B2(n_3649),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3591),
.Y(n_3739)
);

OR2x2_ASAP7_75t_L g3740 ( 
.A(n_3591),
.B(n_3549),
.Y(n_3740)
);

AOI21xp33_ASAP7_75t_L g3741 ( 
.A1(n_3615),
.A2(n_3580),
.B(n_3650),
.Y(n_3741)
);

CKINVDCx11_ASAP7_75t_R g3742 ( 
.A(n_3606),
.Y(n_3742)
);

OAI21xp5_ASAP7_75t_SL g3743 ( 
.A1(n_3551),
.A2(n_3524),
.B(n_3286),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_L g3744 ( 
.A(n_3615),
.B(n_3500),
.Y(n_3744)
);

AOI22xp33_ASAP7_75t_SL g3745 ( 
.A1(n_3615),
.A2(n_3581),
.B1(n_3603),
.B2(n_3551),
.Y(n_3745)
);

OR2x2_ASAP7_75t_L g3746 ( 
.A(n_3688),
.B(n_3691),
.Y(n_3746)
);

AND2x2_ASAP7_75t_L g3747 ( 
.A(n_3713),
.B(n_3709),
.Y(n_3747)
);

OR2x2_ASAP7_75t_L g3748 ( 
.A(n_3698),
.B(n_3705),
.Y(n_3748)
);

NAND2xp5_ASAP7_75t_L g3749 ( 
.A(n_3673),
.B(n_3667),
.Y(n_3749)
);

INVx2_ASAP7_75t_L g3750 ( 
.A(n_3736),
.Y(n_3750)
);

INVx2_ASAP7_75t_L g3751 ( 
.A(n_3736),
.Y(n_3751)
);

INVx2_ASAP7_75t_L g3752 ( 
.A(n_3739),
.Y(n_3752)
);

INVx2_ASAP7_75t_L g3753 ( 
.A(n_3726),
.Y(n_3753)
);

BUFx6f_ASAP7_75t_L g3754 ( 
.A(n_3684),
.Y(n_3754)
);

AND2x2_ASAP7_75t_L g3755 ( 
.A(n_3731),
.B(n_3659),
.Y(n_3755)
);

AND2x2_ASAP7_75t_L g3756 ( 
.A(n_3723),
.B(n_3674),
.Y(n_3756)
);

OA21x2_ASAP7_75t_L g3757 ( 
.A1(n_3741),
.A2(n_3737),
.B(n_3734),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_3679),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3686),
.Y(n_3759)
);

BUFx6f_ASAP7_75t_L g3760 ( 
.A(n_3684),
.Y(n_3760)
);

OR2x2_ASAP7_75t_L g3761 ( 
.A(n_3744),
.B(n_3680),
.Y(n_3761)
);

INVx2_ASAP7_75t_L g3762 ( 
.A(n_3666),
.Y(n_3762)
);

OAI21x1_ASAP7_75t_L g3763 ( 
.A1(n_3729),
.A2(n_3721),
.B(n_3715),
.Y(n_3763)
);

BUFx3_ASAP7_75t_L g3764 ( 
.A(n_3669),
.Y(n_3764)
);

BUFx2_ASAP7_75t_L g3765 ( 
.A(n_3701),
.Y(n_3765)
);

AND2x2_ASAP7_75t_L g3766 ( 
.A(n_3702),
.B(n_3735),
.Y(n_3766)
);

CKINVDCx5p33_ASAP7_75t_R g3767 ( 
.A(n_3742),
.Y(n_3767)
);

BUFx3_ASAP7_75t_L g3768 ( 
.A(n_3661),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_3727),
.Y(n_3769)
);

AOI22xp33_ASAP7_75t_L g3770 ( 
.A1(n_3745),
.A2(n_3654),
.B1(n_3655),
.B2(n_3738),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_3727),
.Y(n_3771)
);

HB1xp67_ASAP7_75t_L g3772 ( 
.A(n_3678),
.Y(n_3772)
);

OR2x2_ASAP7_75t_L g3773 ( 
.A(n_3719),
.B(n_3653),
.Y(n_3773)
);

INVx2_ASAP7_75t_L g3774 ( 
.A(n_3740),
.Y(n_3774)
);

AO21x2_ASAP7_75t_L g3775 ( 
.A1(n_3721),
.A2(n_3732),
.B(n_3737),
.Y(n_3775)
);

INVx2_ASAP7_75t_L g3776 ( 
.A(n_3677),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3687),
.Y(n_3777)
);

AND2x2_ASAP7_75t_L g3778 ( 
.A(n_3745),
.B(n_3711),
.Y(n_3778)
);

BUFx2_ASAP7_75t_L g3779 ( 
.A(n_3692),
.Y(n_3779)
);

INVx2_ASAP7_75t_L g3780 ( 
.A(n_3660),
.Y(n_3780)
);

HB1xp67_ASAP7_75t_L g3781 ( 
.A(n_3670),
.Y(n_3781)
);

HB1xp67_ASAP7_75t_L g3782 ( 
.A(n_3733),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3707),
.Y(n_3783)
);

AOI221xp5_ASAP7_75t_L g3784 ( 
.A1(n_3743),
.A2(n_3732),
.B1(n_3714),
.B2(n_3668),
.C(n_3657),
.Y(n_3784)
);

OA21x2_ASAP7_75t_L g3785 ( 
.A1(n_3716),
.A2(n_3710),
.B(n_3672),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_3656),
.Y(n_3786)
);

AO21x2_ASAP7_75t_L g3787 ( 
.A1(n_3663),
.A2(n_3720),
.B(n_3718),
.Y(n_3787)
);

AND2x2_ASAP7_75t_L g3788 ( 
.A(n_3689),
.B(n_3690),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3658),
.Y(n_3789)
);

AO21x2_ASAP7_75t_L g3790 ( 
.A1(n_3663),
.A2(n_3699),
.B(n_3685),
.Y(n_3790)
);

AND2x2_ASAP7_75t_L g3791 ( 
.A(n_3689),
.B(n_3690),
.Y(n_3791)
);

AND2x2_ASAP7_75t_L g3792 ( 
.A(n_3662),
.B(n_3682),
.Y(n_3792)
);

OAI21xp5_ASAP7_75t_L g3793 ( 
.A1(n_3654),
.A2(n_3662),
.B(n_3667),
.Y(n_3793)
);

INVx3_ASAP7_75t_L g3794 ( 
.A(n_3712),
.Y(n_3794)
);

AND2x2_ASAP7_75t_L g3795 ( 
.A(n_3682),
.B(n_3722),
.Y(n_3795)
);

INVx3_ASAP7_75t_L g3796 ( 
.A(n_3693),
.Y(n_3796)
);

INVx1_ASAP7_75t_L g3797 ( 
.A(n_3706),
.Y(n_3797)
);

AND2x2_ASAP7_75t_L g3798 ( 
.A(n_3671),
.B(n_3704),
.Y(n_3798)
);

INVx2_ASAP7_75t_L g3799 ( 
.A(n_3665),
.Y(n_3799)
);

AOI22xp33_ASAP7_75t_L g3800 ( 
.A1(n_3708),
.A2(n_3717),
.B1(n_3671),
.B2(n_3724),
.Y(n_3800)
);

INVx2_ASAP7_75t_L g3801 ( 
.A(n_3665),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3717),
.Y(n_3802)
);

INVx1_ASAP7_75t_L g3803 ( 
.A(n_3676),
.Y(n_3803)
);

INVx1_ASAP7_75t_L g3804 ( 
.A(n_3676),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3664),
.Y(n_3805)
);

AO21x2_ASAP7_75t_L g3806 ( 
.A1(n_3685),
.A2(n_3699),
.B(n_3700),
.Y(n_3806)
);

AND2x2_ASAP7_75t_L g3807 ( 
.A(n_3675),
.B(n_3730),
.Y(n_3807)
);

AND2x2_ASAP7_75t_L g3808 ( 
.A(n_3730),
.B(n_3696),
.Y(n_3808)
);

NAND2xp5_ASAP7_75t_L g3809 ( 
.A(n_3683),
.B(n_3725),
.Y(n_3809)
);

BUFx3_ASAP7_75t_L g3810 ( 
.A(n_3681),
.Y(n_3810)
);

INVx2_ASAP7_75t_L g3811 ( 
.A(n_3728),
.Y(n_3811)
);

AND2x4_ASAP7_75t_L g3812 ( 
.A(n_3697),
.B(n_3703),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3725),
.Y(n_3813)
);

AO21x2_ASAP7_75t_L g3814 ( 
.A1(n_3695),
.A2(n_3741),
.B(n_3721),
.Y(n_3814)
);

HB1xp67_ASAP7_75t_L g3815 ( 
.A(n_3688),
.Y(n_3815)
);

OA21x2_ASAP7_75t_L g3816 ( 
.A1(n_3673),
.A2(n_3741),
.B(n_3737),
.Y(n_3816)
);

AND2x4_ASAP7_75t_L g3817 ( 
.A(n_3709),
.B(n_3713),
.Y(n_3817)
);

INVx2_ASAP7_75t_L g3818 ( 
.A(n_3736),
.Y(n_3818)
);

AOI22xp33_ASAP7_75t_L g3819 ( 
.A1(n_3736),
.A2(n_3745),
.B1(n_3654),
.B2(n_3655),
.Y(n_3819)
);

INVx2_ASAP7_75t_L g3820 ( 
.A(n_3736),
.Y(n_3820)
);

HB1xp67_ASAP7_75t_L g3821 ( 
.A(n_3688),
.Y(n_3821)
);

INVx2_ASAP7_75t_L g3822 ( 
.A(n_3736),
.Y(n_3822)
);

HB1xp67_ASAP7_75t_L g3823 ( 
.A(n_3688),
.Y(n_3823)
);

INVx2_ASAP7_75t_L g3824 ( 
.A(n_3736),
.Y(n_3824)
);

BUFx2_ASAP7_75t_L g3825 ( 
.A(n_3701),
.Y(n_3825)
);

OR2x6_ASAP7_75t_L g3826 ( 
.A(n_3694),
.B(n_3639),
.Y(n_3826)
);

AND2x2_ASAP7_75t_L g3827 ( 
.A(n_3713),
.B(n_3709),
.Y(n_3827)
);

AO21x2_ASAP7_75t_L g3828 ( 
.A1(n_3741),
.A2(n_3721),
.B(n_3694),
.Y(n_3828)
);

HB1xp67_ASAP7_75t_L g3829 ( 
.A(n_3688),
.Y(n_3829)
);

BUFx3_ASAP7_75t_L g3830 ( 
.A(n_3684),
.Y(n_3830)
);

HB1xp67_ASAP7_75t_L g3831 ( 
.A(n_3688),
.Y(n_3831)
);

AND2x2_ASAP7_75t_L g3832 ( 
.A(n_3713),
.B(n_3709),
.Y(n_3832)
);

NOR2xp33_ASAP7_75t_L g3833 ( 
.A(n_3742),
.B(n_3661),
.Y(n_3833)
);

INVx6_ASAP7_75t_SL g3834 ( 
.A(n_3817),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3752),
.Y(n_3835)
);

AND2x2_ASAP7_75t_SL g3836 ( 
.A(n_3802),
.B(n_3803),
.Y(n_3836)
);

INVx3_ASAP7_75t_L g3837 ( 
.A(n_3775),
.Y(n_3837)
);

INVx2_ASAP7_75t_L g3838 ( 
.A(n_3775),
.Y(n_3838)
);

AND2x2_ASAP7_75t_L g3839 ( 
.A(n_3788),
.B(n_3791),
.Y(n_3839)
);

AND2x4_ASAP7_75t_L g3840 ( 
.A(n_3817),
.B(n_3779),
.Y(n_3840)
);

INVxp67_ASAP7_75t_L g3841 ( 
.A(n_3765),
.Y(n_3841)
);

OR2x2_ASAP7_75t_SL g3842 ( 
.A(n_3802),
.B(n_3803),
.Y(n_3842)
);

AOI22xp33_ASAP7_75t_SL g3843 ( 
.A1(n_3775),
.A2(n_3778),
.B1(n_3816),
.B2(n_3807),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3752),
.Y(n_3844)
);

AND2x2_ASAP7_75t_L g3845 ( 
.A(n_3788),
.B(n_3791),
.Y(n_3845)
);

AND2x2_ASAP7_75t_L g3846 ( 
.A(n_3747),
.B(n_3827),
.Y(n_3846)
);

OR2x2_ASAP7_75t_L g3847 ( 
.A(n_3804),
.B(n_3746),
.Y(n_3847)
);

AND2x2_ASAP7_75t_L g3848 ( 
.A(n_3747),
.B(n_3827),
.Y(n_3848)
);

BUFx3_ASAP7_75t_L g3849 ( 
.A(n_3764),
.Y(n_3849)
);

INVx1_ASAP7_75t_L g3850 ( 
.A(n_3769),
.Y(n_3850)
);

INVx1_ASAP7_75t_L g3851 ( 
.A(n_3769),
.Y(n_3851)
);

INVx3_ASAP7_75t_L g3852 ( 
.A(n_3830),
.Y(n_3852)
);

BUFx4f_ASAP7_75t_L g3853 ( 
.A(n_3754),
.Y(n_3853)
);

INVx2_ASAP7_75t_L g3854 ( 
.A(n_3790),
.Y(n_3854)
);

AND2x2_ASAP7_75t_L g3855 ( 
.A(n_3832),
.B(n_3755),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3771),
.Y(n_3856)
);

OR2x2_ASAP7_75t_L g3857 ( 
.A(n_3804),
.B(n_3746),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_L g3858 ( 
.A(n_3781),
.B(n_3749),
.Y(n_3858)
);

NAND2xp5_ASAP7_75t_L g3859 ( 
.A(n_3808),
.B(n_3815),
.Y(n_3859)
);

INVx3_ASAP7_75t_L g3860 ( 
.A(n_3830),
.Y(n_3860)
);

AOI221xp5_ASAP7_75t_L g3861 ( 
.A1(n_3800),
.A2(n_3770),
.B1(n_3819),
.B2(n_3784),
.C(n_3793),
.Y(n_3861)
);

AND2x2_ASAP7_75t_L g3862 ( 
.A(n_3832),
.B(n_3755),
.Y(n_3862)
);

INVx2_ASAP7_75t_L g3863 ( 
.A(n_3790),
.Y(n_3863)
);

BUFx6f_ASAP7_75t_L g3864 ( 
.A(n_3764),
.Y(n_3864)
);

AND2x4_ASAP7_75t_L g3865 ( 
.A(n_3817),
.B(n_3779),
.Y(n_3865)
);

INVx2_ASAP7_75t_L g3866 ( 
.A(n_3790),
.Y(n_3866)
);

INVx2_ASAP7_75t_L g3867 ( 
.A(n_3828),
.Y(n_3867)
);

INVx2_ASAP7_75t_L g3868 ( 
.A(n_3828),
.Y(n_3868)
);

BUFx3_ASAP7_75t_L g3869 ( 
.A(n_3767),
.Y(n_3869)
);

NAND2x1p5_ASAP7_75t_L g3870 ( 
.A(n_3812),
.B(n_3830),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_L g3871 ( 
.A(n_3808),
.B(n_3821),
.Y(n_3871)
);

INVx1_ASAP7_75t_L g3872 ( 
.A(n_3771),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_3823),
.B(n_3829),
.Y(n_3873)
);

INVx2_ASAP7_75t_L g3874 ( 
.A(n_3828),
.Y(n_3874)
);

AOI22xp33_ASAP7_75t_L g3875 ( 
.A1(n_3789),
.A2(n_3805),
.B1(n_3806),
.B2(n_3812),
.Y(n_3875)
);

OR2x2_ASAP7_75t_L g3876 ( 
.A(n_3748),
.B(n_3777),
.Y(n_3876)
);

AND2x2_ASAP7_75t_L g3877 ( 
.A(n_3817),
.B(n_3765),
.Y(n_3877)
);

AND2x2_ASAP7_75t_L g3878 ( 
.A(n_3825),
.B(n_3756),
.Y(n_3878)
);

HB1xp67_ASAP7_75t_L g3879 ( 
.A(n_3825),
.Y(n_3879)
);

OA21x2_ASAP7_75t_L g3880 ( 
.A1(n_3763),
.A2(n_3783),
.B(n_3798),
.Y(n_3880)
);

INVx2_ASAP7_75t_L g3881 ( 
.A(n_3806),
.Y(n_3881)
);

BUFx2_ASAP7_75t_L g3882 ( 
.A(n_3796),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_L g3883 ( 
.A(n_3831),
.B(n_3807),
.Y(n_3883)
);

AND2x2_ASAP7_75t_L g3884 ( 
.A(n_3756),
.B(n_3794),
.Y(n_3884)
);

AND2x4_ASAP7_75t_L g3885 ( 
.A(n_3796),
.B(n_3794),
.Y(n_3885)
);

NAND2xp5_ASAP7_75t_L g3886 ( 
.A(n_3772),
.B(n_3786),
.Y(n_3886)
);

OR2x2_ASAP7_75t_L g3887 ( 
.A(n_3748),
.B(n_3777),
.Y(n_3887)
);

INVx2_ASAP7_75t_L g3888 ( 
.A(n_3806),
.Y(n_3888)
);

HB1xp67_ASAP7_75t_L g3889 ( 
.A(n_3796),
.Y(n_3889)
);

INVx3_ASAP7_75t_L g3890 ( 
.A(n_3754),
.Y(n_3890)
);

AND2x2_ASAP7_75t_L g3891 ( 
.A(n_3794),
.B(n_3766),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_L g3892 ( 
.A(n_3786),
.B(n_3778),
.Y(n_3892)
);

AND2x2_ASAP7_75t_L g3893 ( 
.A(n_3766),
.B(n_3813),
.Y(n_3893)
);

INVx1_ASAP7_75t_L g3894 ( 
.A(n_3758),
.Y(n_3894)
);

AND2x2_ASAP7_75t_L g3895 ( 
.A(n_3813),
.B(n_3795),
.Y(n_3895)
);

AND2x2_ASAP7_75t_L g3896 ( 
.A(n_3795),
.B(n_3797),
.Y(n_3896)
);

BUFx3_ASAP7_75t_L g3897 ( 
.A(n_3767),
.Y(n_3897)
);

INVxp67_ASAP7_75t_L g3898 ( 
.A(n_3799),
.Y(n_3898)
);

INVx2_ASAP7_75t_L g3899 ( 
.A(n_3816),
.Y(n_3899)
);

AND2x2_ASAP7_75t_L g3900 ( 
.A(n_3797),
.B(n_3768),
.Y(n_3900)
);

INVx2_ASAP7_75t_L g3901 ( 
.A(n_3816),
.Y(n_3901)
);

HB1xp67_ASAP7_75t_L g3902 ( 
.A(n_3782),
.Y(n_3902)
);

AND2x2_ASAP7_75t_L g3903 ( 
.A(n_3768),
.B(n_3798),
.Y(n_3903)
);

AND2x4_ASAP7_75t_SL g3904 ( 
.A(n_3754),
.B(n_3760),
.Y(n_3904)
);

NAND2xp5_ASAP7_75t_L g3905 ( 
.A(n_3750),
.B(n_3751),
.Y(n_3905)
);

INVx2_ASAP7_75t_L g3906 ( 
.A(n_3816),
.Y(n_3906)
);

AND2x2_ASAP7_75t_L g3907 ( 
.A(n_3768),
.B(n_3792),
.Y(n_3907)
);

AND2x4_ASAP7_75t_SL g3908 ( 
.A(n_3754),
.B(n_3760),
.Y(n_3908)
);

INVx2_ASAP7_75t_L g3909 ( 
.A(n_3814),
.Y(n_3909)
);

INVx4_ASAP7_75t_L g3910 ( 
.A(n_3754),
.Y(n_3910)
);

HB1xp67_ASAP7_75t_L g3911 ( 
.A(n_3799),
.Y(n_3911)
);

INVx2_ASAP7_75t_L g3912 ( 
.A(n_3814),
.Y(n_3912)
);

OR2x2_ASAP7_75t_L g3913 ( 
.A(n_3761),
.B(n_3773),
.Y(n_3913)
);

OR2x2_ASAP7_75t_L g3914 ( 
.A(n_3761),
.B(n_3773),
.Y(n_3914)
);

BUFx3_ASAP7_75t_L g3915 ( 
.A(n_3760),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3759),
.Y(n_3916)
);

NOR2xp33_ASAP7_75t_L g3917 ( 
.A(n_3760),
.B(n_3833),
.Y(n_3917)
);

AND2x2_ASAP7_75t_L g3918 ( 
.A(n_3792),
.B(n_3809),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_3899),
.Y(n_3919)
);

NAND2xp5_ASAP7_75t_L g3920 ( 
.A(n_3843),
.B(n_3899),
.Y(n_3920)
);

INVx2_ASAP7_75t_L g3921 ( 
.A(n_3842),
.Y(n_3921)
);

INVx2_ASAP7_75t_L g3922 ( 
.A(n_3842),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3901),
.Y(n_3923)
);

INVx4_ASAP7_75t_L g3924 ( 
.A(n_3864),
.Y(n_3924)
);

AND2x4_ASAP7_75t_L g3925 ( 
.A(n_3840),
.B(n_3787),
.Y(n_3925)
);

INVx2_ASAP7_75t_L g3926 ( 
.A(n_3837),
.Y(n_3926)
);

AND2x2_ASAP7_75t_L g3927 ( 
.A(n_3877),
.B(n_3814),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3901),
.Y(n_3928)
);

INVxp67_ASAP7_75t_SL g3929 ( 
.A(n_3837),
.Y(n_3929)
);

CKINVDCx5p33_ASAP7_75t_R g3930 ( 
.A(n_3869),
.Y(n_3930)
);

INVx2_ASAP7_75t_L g3931 ( 
.A(n_3837),
.Y(n_3931)
);

INVx2_ASAP7_75t_L g3932 ( 
.A(n_3836),
.Y(n_3932)
);

BUFx2_ASAP7_75t_L g3933 ( 
.A(n_3834),
.Y(n_3933)
);

NOR2xp33_ASAP7_75t_L g3934 ( 
.A(n_3864),
.B(n_3760),
.Y(n_3934)
);

AND2x2_ASAP7_75t_L g3935 ( 
.A(n_3877),
.B(n_3787),
.Y(n_3935)
);

INVx2_ASAP7_75t_L g3936 ( 
.A(n_3836),
.Y(n_3936)
);

HB1xp67_ASAP7_75t_L g3937 ( 
.A(n_3879),
.Y(n_3937)
);

AND2x2_ASAP7_75t_L g3938 ( 
.A(n_3878),
.B(n_3787),
.Y(n_3938)
);

HB1xp67_ASAP7_75t_L g3939 ( 
.A(n_3841),
.Y(n_3939)
);

INVx3_ASAP7_75t_L g3940 ( 
.A(n_3870),
.Y(n_3940)
);

INVx2_ASAP7_75t_L g3941 ( 
.A(n_3836),
.Y(n_3941)
);

BUFx3_ASAP7_75t_L g3942 ( 
.A(n_3869),
.Y(n_3942)
);

AND2x2_ASAP7_75t_L g3943 ( 
.A(n_3878),
.B(n_3763),
.Y(n_3943)
);

OR2x2_ASAP7_75t_L g3944 ( 
.A(n_3906),
.B(n_3789),
.Y(n_3944)
);

BUFx6f_ASAP7_75t_L g3945 ( 
.A(n_3864),
.Y(n_3945)
);

AND2x2_ASAP7_75t_L g3946 ( 
.A(n_3855),
.B(n_3785),
.Y(n_3946)
);

INVx2_ASAP7_75t_L g3947 ( 
.A(n_3867),
.Y(n_3947)
);

HB1xp67_ASAP7_75t_L g3948 ( 
.A(n_3911),
.Y(n_3948)
);

OR2x2_ASAP7_75t_L g3949 ( 
.A(n_3906),
.B(n_3785),
.Y(n_3949)
);

INVx2_ASAP7_75t_L g3950 ( 
.A(n_3867),
.Y(n_3950)
);

AND2x4_ASAP7_75t_L g3951 ( 
.A(n_3840),
.B(n_3826),
.Y(n_3951)
);

AND2x2_ASAP7_75t_L g3952 ( 
.A(n_3855),
.B(n_3785),
.Y(n_3952)
);

INVx2_ASAP7_75t_L g3953 ( 
.A(n_3868),
.Y(n_3953)
);

INVx2_ASAP7_75t_L g3954 ( 
.A(n_3868),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3874),
.Y(n_3955)
);

HB1xp67_ASAP7_75t_L g3956 ( 
.A(n_3870),
.Y(n_3956)
);

INVx2_ASAP7_75t_L g3957 ( 
.A(n_3874),
.Y(n_3957)
);

INVx2_ASAP7_75t_L g3958 ( 
.A(n_3909),
.Y(n_3958)
);

INVx1_ASAP7_75t_L g3959 ( 
.A(n_3881),
.Y(n_3959)
);

INVxp67_ASAP7_75t_L g3960 ( 
.A(n_3864),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3881),
.Y(n_3961)
);

HB1xp67_ASAP7_75t_L g3962 ( 
.A(n_3870),
.Y(n_3962)
);

CKINVDCx5p33_ASAP7_75t_R g3963 ( 
.A(n_3897),
.Y(n_3963)
);

INVx2_ASAP7_75t_L g3964 ( 
.A(n_3909),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3888),
.Y(n_3965)
);

INVx1_ASAP7_75t_L g3966 ( 
.A(n_3888),
.Y(n_3966)
);

HB1xp67_ASAP7_75t_L g3967 ( 
.A(n_3898),
.Y(n_3967)
);

BUFx12f_ASAP7_75t_L g3968 ( 
.A(n_3864),
.Y(n_3968)
);

INVx2_ASAP7_75t_L g3969 ( 
.A(n_3912),
.Y(n_3969)
);

AND2x2_ASAP7_75t_L g3970 ( 
.A(n_3862),
.B(n_3785),
.Y(n_3970)
);

INVxp67_ASAP7_75t_L g3971 ( 
.A(n_3849),
.Y(n_3971)
);

HB1xp67_ASAP7_75t_L g3972 ( 
.A(n_3849),
.Y(n_3972)
);

AND2x2_ASAP7_75t_L g3973 ( 
.A(n_3972),
.B(n_3862),
.Y(n_3973)
);

INVx1_ASAP7_75t_L g3974 ( 
.A(n_3929),
.Y(n_3974)
);

INVx2_ASAP7_75t_L g3975 ( 
.A(n_3921),
.Y(n_3975)
);

NAND2xp5_ASAP7_75t_L g3976 ( 
.A(n_3938),
.B(n_3854),
.Y(n_3976)
);

INVx1_ASAP7_75t_L g3977 ( 
.A(n_3929),
.Y(n_3977)
);

NOR2xp33_ASAP7_75t_L g3978 ( 
.A(n_3942),
.B(n_3897),
.Y(n_3978)
);

INVx1_ASAP7_75t_L g3979 ( 
.A(n_3921),
.Y(n_3979)
);

INVx2_ASAP7_75t_L g3980 ( 
.A(n_3921),
.Y(n_3980)
);

AND2x4_ASAP7_75t_L g3981 ( 
.A(n_3921),
.B(n_3840),
.Y(n_3981)
);

INVx2_ASAP7_75t_L g3982 ( 
.A(n_3922),
.Y(n_3982)
);

INVx1_ASAP7_75t_L g3983 ( 
.A(n_3922),
.Y(n_3983)
);

BUFx2_ASAP7_75t_L g3984 ( 
.A(n_3938),
.Y(n_3984)
);

NOR2xp33_ASAP7_75t_L g3985 ( 
.A(n_3942),
.B(n_3801),
.Y(n_3985)
);

NAND2x1p5_ASAP7_75t_L g3986 ( 
.A(n_3924),
.B(n_3910),
.Y(n_3986)
);

NOR2xp33_ASAP7_75t_L g3987 ( 
.A(n_3942),
.B(n_3801),
.Y(n_3987)
);

NAND2xp5_ASAP7_75t_L g3988 ( 
.A(n_3938),
.B(n_3854),
.Y(n_3988)
);

HB1xp67_ASAP7_75t_L g3989 ( 
.A(n_3972),
.Y(n_3989)
);

AND2x2_ASAP7_75t_L g3990 ( 
.A(n_3943),
.B(n_3846),
.Y(n_3990)
);

NOR2xp33_ASAP7_75t_L g3991 ( 
.A(n_3942),
.B(n_3810),
.Y(n_3991)
);

INVx2_ASAP7_75t_L g3992 ( 
.A(n_3922),
.Y(n_3992)
);

INVx1_ASAP7_75t_L g3993 ( 
.A(n_3922),
.Y(n_3993)
);

INVxp67_ASAP7_75t_L g3994 ( 
.A(n_3967),
.Y(n_3994)
);

INVx2_ASAP7_75t_L g3995 ( 
.A(n_3932),
.Y(n_3995)
);

INVx1_ASAP7_75t_L g3996 ( 
.A(n_3920),
.Y(n_3996)
);

INVx1_ASAP7_75t_SL g3997 ( 
.A(n_3920),
.Y(n_3997)
);

AND2x2_ASAP7_75t_L g3998 ( 
.A(n_3943),
.B(n_3846),
.Y(n_3998)
);

HB1xp67_ASAP7_75t_L g3999 ( 
.A(n_3948),
.Y(n_3999)
);

AND2x2_ASAP7_75t_L g4000 ( 
.A(n_3943),
.B(n_3848),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_3926),
.Y(n_4001)
);

HB1xp67_ASAP7_75t_L g4002 ( 
.A(n_3948),
.Y(n_4002)
);

AND2x2_ASAP7_75t_L g4003 ( 
.A(n_3946),
.B(n_3848),
.Y(n_4003)
);

AND2x2_ASAP7_75t_L g4004 ( 
.A(n_3946),
.B(n_3865),
.Y(n_4004)
);

NAND3xp33_ASAP7_75t_L g4005 ( 
.A(n_3932),
.B(n_3912),
.C(n_3875),
.Y(n_4005)
);

AND2x4_ASAP7_75t_L g4006 ( 
.A(n_3932),
.B(n_3865),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3926),
.Y(n_4007)
);

AND2x2_ASAP7_75t_L g4008 ( 
.A(n_3946),
.B(n_3865),
.Y(n_4008)
);

AND2x2_ASAP7_75t_L g4009 ( 
.A(n_3952),
.B(n_3907),
.Y(n_4009)
);

AND2x2_ASAP7_75t_L g4010 ( 
.A(n_3952),
.B(n_3907),
.Y(n_4010)
);

NAND2xp5_ASAP7_75t_L g4011 ( 
.A(n_3935),
.B(n_3863),
.Y(n_4011)
);

INVx1_ASAP7_75t_L g4012 ( 
.A(n_3926),
.Y(n_4012)
);

INVx2_ASAP7_75t_L g4013 ( 
.A(n_3932),
.Y(n_4013)
);

OR2x2_ASAP7_75t_L g4014 ( 
.A(n_3936),
.B(n_3883),
.Y(n_4014)
);

OAI21xp33_ASAP7_75t_L g4015 ( 
.A1(n_3927),
.A2(n_3903),
.B(n_3859),
.Y(n_4015)
);

HB1xp67_ASAP7_75t_L g4016 ( 
.A(n_3945),
.Y(n_4016)
);

NOR2xp33_ASAP7_75t_SL g4017 ( 
.A(n_3936),
.B(n_3941),
.Y(n_4017)
);

AOI22xp33_ASAP7_75t_L g4018 ( 
.A1(n_3925),
.A2(n_3863),
.B1(n_3866),
.B2(n_3838),
.Y(n_4018)
);

HB1xp67_ASAP7_75t_L g4019 ( 
.A(n_3945),
.Y(n_4019)
);

NAND2xp5_ASAP7_75t_L g4020 ( 
.A(n_3935),
.B(n_3866),
.Y(n_4020)
);

AND2x2_ASAP7_75t_L g4021 ( 
.A(n_3952),
.B(n_3903),
.Y(n_4021)
);

AND2x2_ASAP7_75t_L g4022 ( 
.A(n_3970),
.B(n_3891),
.Y(n_4022)
);

BUFx2_ASAP7_75t_L g4023 ( 
.A(n_3968),
.Y(n_4023)
);

AND2x2_ASAP7_75t_L g4024 ( 
.A(n_3970),
.B(n_3891),
.Y(n_4024)
);

INVxp67_ASAP7_75t_SL g4025 ( 
.A(n_3984),
.Y(n_4025)
);

INVx1_ASAP7_75t_L g4026 ( 
.A(n_3984),
.Y(n_4026)
);

INVx1_ASAP7_75t_L g4027 ( 
.A(n_3975),
.Y(n_4027)
);

INVx1_ASAP7_75t_L g4028 ( 
.A(n_3975),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_3975),
.Y(n_4029)
);

OR2x2_ASAP7_75t_L g4030 ( 
.A(n_3997),
.B(n_3996),
.Y(n_4030)
);

AND2x2_ASAP7_75t_L g4031 ( 
.A(n_3990),
.B(n_3882),
.Y(n_4031)
);

BUFx2_ASAP7_75t_L g4032 ( 
.A(n_4004),
.Y(n_4032)
);

NOR2x1_ASAP7_75t_R g4033 ( 
.A(n_4023),
.B(n_3963),
.Y(n_4033)
);

INVx2_ASAP7_75t_L g4034 ( 
.A(n_3980),
.Y(n_4034)
);

AND2x2_ASAP7_75t_L g4035 ( 
.A(n_3990),
.B(n_3882),
.Y(n_4035)
);

AND2x2_ASAP7_75t_L g4036 ( 
.A(n_3998),
.B(n_3885),
.Y(n_4036)
);

OR2x2_ASAP7_75t_L g4037 ( 
.A(n_3997),
.B(n_3936),
.Y(n_4037)
);

HB1xp67_ASAP7_75t_L g4038 ( 
.A(n_4004),
.Y(n_4038)
);

INVx2_ASAP7_75t_L g4039 ( 
.A(n_3980),
.Y(n_4039)
);

BUFx2_ASAP7_75t_L g4040 ( 
.A(n_4008),
.Y(n_4040)
);

INVx1_ASAP7_75t_L g4041 ( 
.A(n_3980),
.Y(n_4041)
);

NAND2xp5_ASAP7_75t_L g4042 ( 
.A(n_3996),
.B(n_3936),
.Y(n_4042)
);

HB1xp67_ASAP7_75t_L g4043 ( 
.A(n_4008),
.Y(n_4043)
);

AND2x2_ASAP7_75t_L g4044 ( 
.A(n_3998),
.B(n_3885),
.Y(n_4044)
);

INVx1_ASAP7_75t_L g4045 ( 
.A(n_3982),
.Y(n_4045)
);

AND2x2_ASAP7_75t_L g4046 ( 
.A(n_4000),
.B(n_3885),
.Y(n_4046)
);

AND2x2_ASAP7_75t_L g4047 ( 
.A(n_4000),
.B(n_3884),
.Y(n_4047)
);

OR2x2_ASAP7_75t_L g4048 ( 
.A(n_4021),
.B(n_3941),
.Y(n_4048)
);

AND2x2_ASAP7_75t_L g4049 ( 
.A(n_4003),
.B(n_3884),
.Y(n_4049)
);

INVx2_ASAP7_75t_L g4050 ( 
.A(n_3982),
.Y(n_4050)
);

OR2x2_ASAP7_75t_L g4051 ( 
.A(n_4021),
.B(n_3941),
.Y(n_4051)
);

NAND2xp5_ASAP7_75t_L g4052 ( 
.A(n_4003),
.B(n_3941),
.Y(n_4052)
);

AND2x2_ASAP7_75t_L g4053 ( 
.A(n_4009),
.B(n_3900),
.Y(n_4053)
);

INVx1_ASAP7_75t_L g4054 ( 
.A(n_3982),
.Y(n_4054)
);

AND2x2_ASAP7_75t_L g4055 ( 
.A(n_4009),
.B(n_3900),
.Y(n_4055)
);

INVx1_ASAP7_75t_L g4056 ( 
.A(n_3992),
.Y(n_4056)
);

INVx1_ASAP7_75t_L g4057 ( 
.A(n_3992),
.Y(n_4057)
);

AND2x2_ASAP7_75t_L g4058 ( 
.A(n_4010),
.B(n_3889),
.Y(n_4058)
);

AND2x2_ASAP7_75t_L g4059 ( 
.A(n_4010),
.B(n_4022),
.Y(n_4059)
);

AND2x2_ASAP7_75t_L g4060 ( 
.A(n_4022),
.B(n_3852),
.Y(n_4060)
);

INVx2_ASAP7_75t_L g4061 ( 
.A(n_3992),
.Y(n_4061)
);

INVxp67_ASAP7_75t_L g4062 ( 
.A(n_4017),
.Y(n_4062)
);

AND2x4_ASAP7_75t_SL g4063 ( 
.A(n_3981),
.B(n_3852),
.Y(n_4063)
);

NAND3xp33_ASAP7_75t_L g4064 ( 
.A(n_4062),
.B(n_4005),
.C(n_4017),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_4032),
.Y(n_4065)
);

INVx2_ASAP7_75t_L g4066 ( 
.A(n_4034),
.Y(n_4066)
);

OR2x2_ASAP7_75t_L g4067 ( 
.A(n_4032),
.B(n_4024),
.Y(n_4067)
);

AND2x4_ASAP7_75t_L g4068 ( 
.A(n_4063),
.B(n_3981),
.Y(n_4068)
);

OR2x2_ASAP7_75t_L g4069 ( 
.A(n_4040),
.B(n_4024),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_4040),
.Y(n_4070)
);

AND2x2_ASAP7_75t_L g4071 ( 
.A(n_4053),
.B(n_4055),
.Y(n_4071)
);

NAND2xp5_ASAP7_75t_L g4072 ( 
.A(n_4053),
.B(n_3973),
.Y(n_4072)
);

OR2x2_ASAP7_75t_L g4073 ( 
.A(n_4038),
.B(n_3967),
.Y(n_4073)
);

AND2x2_ASAP7_75t_L g4074 ( 
.A(n_4055),
.B(n_3973),
.Y(n_4074)
);

OR2x2_ASAP7_75t_L g4075 ( 
.A(n_4043),
.B(n_3970),
.Y(n_4075)
);

AND2x2_ASAP7_75t_L g4076 ( 
.A(n_4059),
.B(n_3852),
.Y(n_4076)
);

INVx1_ASAP7_75t_L g4077 ( 
.A(n_4059),
.Y(n_4077)
);

NAND2xp5_ASAP7_75t_L g4078 ( 
.A(n_4031),
.B(n_3935),
.Y(n_4078)
);

AND2x2_ASAP7_75t_L g4079 ( 
.A(n_4049),
.B(n_3860),
.Y(n_4079)
);

NOR3xp33_ASAP7_75t_L g4080 ( 
.A(n_4062),
.B(n_4005),
.C(n_4015),
.Y(n_4080)
);

OR2x2_ASAP7_75t_L g4081 ( 
.A(n_4052),
.B(n_3971),
.Y(n_4081)
);

INVx3_ASAP7_75t_L g4082 ( 
.A(n_4063),
.Y(n_4082)
);

AND2x2_ASAP7_75t_L g4083 ( 
.A(n_4049),
.B(n_3860),
.Y(n_4083)
);

INVx1_ASAP7_75t_L g4084 ( 
.A(n_4027),
.Y(n_4084)
);

AND2x2_ASAP7_75t_L g4085 ( 
.A(n_4047),
.B(n_3860),
.Y(n_4085)
);

INVx1_ASAP7_75t_L g4086 ( 
.A(n_4027),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_4028),
.Y(n_4087)
);

INVx1_ASAP7_75t_L g4088 ( 
.A(n_4028),
.Y(n_4088)
);

INVx1_ASAP7_75t_SL g4089 ( 
.A(n_4047),
.Y(n_4089)
);

AND2x2_ASAP7_75t_L g4090 ( 
.A(n_4071),
.B(n_4031),
.Y(n_4090)
);

O2A1O1Ixp33_ASAP7_75t_L g4091 ( 
.A1(n_4080),
.A2(n_4030),
.B(n_4025),
.C(n_3994),
.Y(n_4091)
);

BUFx2_ASAP7_75t_SL g4092 ( 
.A(n_4068),
.Y(n_4092)
);

INVx1_ASAP7_75t_L g4093 ( 
.A(n_4071),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_4074),
.Y(n_4094)
);

INVx1_ASAP7_75t_L g4095 ( 
.A(n_4066),
.Y(n_4095)
);

AND2x2_ASAP7_75t_L g4096 ( 
.A(n_4076),
.B(n_4035),
.Y(n_4096)
);

AND2x2_ASAP7_75t_L g4097 ( 
.A(n_4076),
.B(n_4035),
.Y(n_4097)
);

AND2x2_ASAP7_75t_L g4098 ( 
.A(n_4089),
.B(n_4036),
.Y(n_4098)
);

AND2x2_ASAP7_75t_L g4099 ( 
.A(n_4079),
.B(n_4036),
.Y(n_4099)
);

INVx2_ASAP7_75t_L g4100 ( 
.A(n_4066),
.Y(n_4100)
);

NAND2xp5_ASAP7_75t_L g4101 ( 
.A(n_4068),
.B(n_4044),
.Y(n_4101)
);

NAND2xp5_ASAP7_75t_L g4102 ( 
.A(n_4068),
.B(n_4044),
.Y(n_4102)
);

OR2x2_ASAP7_75t_L g4103 ( 
.A(n_4067),
.B(n_3971),
.Y(n_4103)
);

HB1xp67_ASAP7_75t_L g4104 ( 
.A(n_4064),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_4069),
.Y(n_4105)
);

OR2x2_ASAP7_75t_L g4106 ( 
.A(n_4075),
.B(n_3871),
.Y(n_4106)
);

INVx2_ASAP7_75t_SL g4107 ( 
.A(n_4079),
.Y(n_4107)
);

NAND2xp5_ASAP7_75t_L g4108 ( 
.A(n_4083),
.B(n_4046),
.Y(n_4108)
);

CKINVDCx16_ASAP7_75t_R g4109 ( 
.A(n_4073),
.Y(n_4109)
);

NOR3xp33_ASAP7_75t_L g4110 ( 
.A(n_4109),
.B(n_4030),
.C(n_4080),
.Y(n_4110)
);

INVx2_ASAP7_75t_L g4111 ( 
.A(n_4090),
.Y(n_4111)
);

A2O1A1Ixp33_ASAP7_75t_L g4112 ( 
.A1(n_4091),
.A2(n_3927),
.B(n_3925),
.C(n_4015),
.Y(n_4112)
);

INVx2_ASAP7_75t_L g4113 ( 
.A(n_4090),
.Y(n_4113)
);

AND2x2_ASAP7_75t_L g4114 ( 
.A(n_4099),
.B(n_4046),
.Y(n_4114)
);

OR2x2_ASAP7_75t_L g4115 ( 
.A(n_4107),
.B(n_4072),
.Y(n_4115)
);

O2A1O1Ixp33_ASAP7_75t_L g4116 ( 
.A1(n_4104),
.A2(n_4025),
.B(n_4037),
.C(n_4042),
.Y(n_4116)
);

AND2x2_ASAP7_75t_L g4117 ( 
.A(n_4099),
.B(n_4060),
.Y(n_4117)
);

INVx1_ASAP7_75t_L g4118 ( 
.A(n_4100),
.Y(n_4118)
);

AND2x2_ASAP7_75t_L g4119 ( 
.A(n_4098),
.B(n_4060),
.Y(n_4119)
);

OR2x2_ASAP7_75t_L g4120 ( 
.A(n_4107),
.B(n_4078),
.Y(n_4120)
);

OR2x2_ASAP7_75t_L g4121 ( 
.A(n_4093),
.B(n_4077),
.Y(n_4121)
);

NAND2x1_ASAP7_75t_L g4122 ( 
.A(n_4096),
.B(n_3940),
.Y(n_4122)
);

INVx1_ASAP7_75t_L g4123 ( 
.A(n_4100),
.Y(n_4123)
);

NAND2xp5_ASAP7_75t_L g4124 ( 
.A(n_4096),
.B(n_4058),
.Y(n_4124)
);

NAND2xp5_ASAP7_75t_L g4125 ( 
.A(n_4097),
.B(n_4058),
.Y(n_4125)
);

OR2x2_ASAP7_75t_L g4126 ( 
.A(n_4092),
.B(n_4065),
.Y(n_4126)
);

NAND2xp5_ASAP7_75t_L g4127 ( 
.A(n_4114),
.B(n_3927),
.Y(n_4127)
);

OR2x2_ASAP7_75t_L g4128 ( 
.A(n_4124),
.B(n_4108),
.Y(n_4128)
);

INVx2_ASAP7_75t_L g4129 ( 
.A(n_4117),
.Y(n_4129)
);

AND2x2_ASAP7_75t_L g4130 ( 
.A(n_4119),
.B(n_4097),
.Y(n_4130)
);

HB1xp67_ASAP7_75t_L g4131 ( 
.A(n_4125),
.Y(n_4131)
);

NAND2xp5_ASAP7_75t_L g4132 ( 
.A(n_4111),
.B(n_4083),
.Y(n_4132)
);

AND2x2_ASAP7_75t_L g4133 ( 
.A(n_4113),
.B(n_4085),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_L g4134 ( 
.A(n_4110),
.B(n_4085),
.Y(n_4134)
);

AND2x2_ASAP7_75t_L g4135 ( 
.A(n_4115),
.B(n_3896),
.Y(n_4135)
);

INVx1_ASAP7_75t_L g4136 ( 
.A(n_4118),
.Y(n_4136)
);

NAND2xp5_ASAP7_75t_L g4137 ( 
.A(n_4118),
.B(n_3981),
.Y(n_4137)
);

INVx1_ASAP7_75t_L g4138 ( 
.A(n_4123),
.Y(n_4138)
);

AND2x2_ASAP7_75t_L g4139 ( 
.A(n_4130),
.B(n_3896),
.Y(n_4139)
);

INVx1_ASAP7_75t_L g4140 ( 
.A(n_4135),
.Y(n_4140)
);

INVx1_ASAP7_75t_SL g4141 ( 
.A(n_4133),
.Y(n_4141)
);

INVx1_ASAP7_75t_L g4142 ( 
.A(n_4137),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_4127),
.Y(n_4143)
);

INVx2_ASAP7_75t_L g4144 ( 
.A(n_4128),
.Y(n_4144)
);

INVx2_ASAP7_75t_L g4145 ( 
.A(n_4129),
.Y(n_4145)
);

INVxp33_ASAP7_75t_L g4146 ( 
.A(n_4131),
.Y(n_4146)
);

OAI21xp5_ASAP7_75t_L g4147 ( 
.A1(n_4146),
.A2(n_4127),
.B(n_4116),
.Y(n_4147)
);

NAND2xp5_ASAP7_75t_L g4148 ( 
.A(n_4139),
.B(n_3981),
.Y(n_4148)
);

AOI322xp5_ASAP7_75t_L g4149 ( 
.A1(n_4142),
.A2(n_3988),
.A3(n_3976),
.B1(n_4011),
.B2(n_4020),
.C1(n_3838),
.C2(n_3979),
.Y(n_4149)
);

NAND3xp33_ASAP7_75t_L g4150 ( 
.A(n_4146),
.B(n_4104),
.C(n_4134),
.Y(n_4150)
);

AOI22xp5_ASAP7_75t_L g4151 ( 
.A1(n_4141),
.A2(n_4013),
.B1(n_3995),
.B2(n_4037),
.Y(n_4151)
);

NAND2xp5_ASAP7_75t_L g4152 ( 
.A(n_4141),
.B(n_4063),
.Y(n_4152)
);

NAND2xp5_ASAP7_75t_L g4153 ( 
.A(n_4144),
.B(n_4006),
.Y(n_4153)
);

NAND4xp75_ASAP7_75t_L g4154 ( 
.A(n_4143),
.B(n_4132),
.C(n_4105),
.D(n_4095),
.Y(n_4154)
);

NAND2xp5_ASAP7_75t_L g4155 ( 
.A(n_4145),
.B(n_4006),
.Y(n_4155)
);

NOR2xp33_ASAP7_75t_L g4156 ( 
.A(n_4140),
.B(n_4048),
.Y(n_4156)
);

AND2x2_ASAP7_75t_L g4157 ( 
.A(n_4139),
.B(n_3978),
.Y(n_4157)
);

INVx1_ASAP7_75t_L g4158 ( 
.A(n_4139),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_4139),
.Y(n_4159)
);

OR2x2_ASAP7_75t_L g4160 ( 
.A(n_4148),
.B(n_4048),
.Y(n_4160)
);

AOI22xp5_ASAP7_75t_L g4161 ( 
.A1(n_4151),
.A2(n_4013),
.B1(n_3995),
.B2(n_4042),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_4153),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_L g4163 ( 
.A(n_4149),
.B(n_4006),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_4155),
.Y(n_4164)
);

INVx1_ASAP7_75t_L g4165 ( 
.A(n_4156),
.Y(n_4165)
);

OAI211xp5_ASAP7_75t_L g4166 ( 
.A1(n_4147),
.A2(n_4126),
.B(n_4138),
.C(n_4136),
.Y(n_4166)
);

NOR3xp33_ASAP7_75t_L g4167 ( 
.A(n_4150),
.B(n_4123),
.C(n_4120),
.Y(n_4167)
);

INVx1_ASAP7_75t_SL g4168 ( 
.A(n_4157),
.Y(n_4168)
);

OAI21xp5_ASAP7_75t_L g4169 ( 
.A1(n_4152),
.A2(n_4112),
.B(n_4102),
.Y(n_4169)
);

INVx2_ASAP7_75t_L g4170 ( 
.A(n_4154),
.Y(n_4170)
);

OAI21xp5_ASAP7_75t_L g4171 ( 
.A1(n_4158),
.A2(n_4101),
.B(n_4052),
.Y(n_4171)
);

OAI21xp5_ASAP7_75t_L g4172 ( 
.A1(n_4159),
.A2(n_4026),
.B(n_4070),
.Y(n_4172)
);

AND2x2_ASAP7_75t_L g4173 ( 
.A(n_4157),
.B(n_3991),
.Y(n_4173)
);

NAND2xp5_ASAP7_75t_L g4174 ( 
.A(n_4151),
.B(n_4006),
.Y(n_4174)
);

AOI221xp5_ASAP7_75t_L g4175 ( 
.A1(n_4147),
.A2(n_3979),
.B1(n_3993),
.B2(n_3983),
.C(n_3988),
.Y(n_4175)
);

NAND3xp33_ASAP7_75t_L g4176 ( 
.A(n_4150),
.B(n_3976),
.C(n_4011),
.Y(n_4176)
);

AND2x2_ASAP7_75t_L g4177 ( 
.A(n_4157),
.B(n_3893),
.Y(n_4177)
);

NAND2xp5_ASAP7_75t_SL g4178 ( 
.A(n_4151),
.B(n_3945),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_4151),
.Y(n_4179)
);

NAND2xp5_ASAP7_75t_L g4180 ( 
.A(n_4151),
.B(n_3918),
.Y(n_4180)
);

AOI21xp5_ASAP7_75t_L g4181 ( 
.A1(n_4148),
.A2(n_4122),
.B(n_4086),
.Y(n_4181)
);

OAI31xp33_ASAP7_75t_SL g4182 ( 
.A1(n_4176),
.A2(n_4026),
.A3(n_4094),
.B(n_3977),
.Y(n_4182)
);

AOI221x1_ASAP7_75t_L g4183 ( 
.A1(n_4167),
.A2(n_4084),
.B1(n_4088),
.B2(n_4087),
.C(n_3974),
.Y(n_4183)
);

AOI21xp5_ASAP7_75t_L g4184 ( 
.A1(n_4178),
.A2(n_3977),
.B(n_3974),
.Y(n_4184)
);

NAND3xp33_ASAP7_75t_L g4185 ( 
.A(n_4176),
.B(n_4171),
.C(n_4166),
.Y(n_4185)
);

OAI21xp5_ASAP7_75t_L g4186 ( 
.A1(n_4174),
.A2(n_4163),
.B(n_4180),
.Y(n_4186)
);

OAI21xp5_ASAP7_75t_L g4187 ( 
.A1(n_4160),
.A2(n_3993),
.B(n_3983),
.Y(n_4187)
);

INVxp67_ASAP7_75t_L g4188 ( 
.A(n_4173),
.Y(n_4188)
);

OAI221xp5_ASAP7_75t_L g4189 ( 
.A1(n_4161),
.A2(n_3940),
.B1(n_4051),
.B2(n_3956),
.C(n_3962),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_4177),
.Y(n_4190)
);

AOI221x1_ASAP7_75t_L g4191 ( 
.A1(n_4179),
.A2(n_4082),
.B1(n_3985),
.B2(n_3987),
.C(n_3924),
.Y(n_4191)
);

INVx1_ASAP7_75t_SL g4192 ( 
.A(n_4168),
.Y(n_4192)
);

OAI21xp33_ASAP7_75t_L g4193 ( 
.A1(n_4165),
.A2(n_3934),
.B(n_4103),
.Y(n_4193)
);

NAND2xp5_ASAP7_75t_SL g4194 ( 
.A(n_4175),
.B(n_3963),
.Y(n_4194)
);

AOI222xp33_ASAP7_75t_L g4195 ( 
.A1(n_4169),
.A2(n_4020),
.B1(n_3923),
.B2(n_3928),
.C1(n_3919),
.C2(n_3926),
.Y(n_4195)
);

AND2x2_ASAP7_75t_L g4196 ( 
.A(n_4172),
.B(n_3893),
.Y(n_4196)
);

OAI22xp33_ASAP7_75t_SL g4197 ( 
.A1(n_4170),
.A2(n_4051),
.B1(n_3949),
.B2(n_4041),
.Y(n_4197)
);

OAI22xp5_ASAP7_75t_L g4198 ( 
.A1(n_4181),
.A2(n_4014),
.B1(n_4106),
.B2(n_4081),
.Y(n_4198)
);

OAI22xp5_ASAP7_75t_L g4199 ( 
.A1(n_4162),
.A2(n_4014),
.B1(n_3940),
.B2(n_3962),
.Y(n_4199)
);

OAI322xp33_ASAP7_75t_L g4200 ( 
.A1(n_4164),
.A2(n_4121),
.A3(n_3949),
.B1(n_4054),
.B2(n_4057),
.C1(n_4056),
.C2(n_4045),
.Y(n_4200)
);

NAND4xp25_ASAP7_75t_L g4201 ( 
.A(n_4167),
.B(n_4023),
.C(n_4082),
.D(n_3934),
.Y(n_4201)
);

OAI21xp33_ASAP7_75t_L g4202 ( 
.A1(n_4168),
.A2(n_3960),
.B(n_4082),
.Y(n_4202)
);

INVx2_ASAP7_75t_L g4203 ( 
.A(n_4177),
.Y(n_4203)
);

OAI32xp33_ASAP7_75t_L g4204 ( 
.A1(n_4168),
.A2(n_3924),
.A3(n_3960),
.B1(n_3989),
.B2(n_4002),
.Y(n_4204)
);

O2A1O1Ixp33_ASAP7_75t_SL g4205 ( 
.A1(n_4178),
.A2(n_3999),
.B(n_3939),
.C(n_3937),
.Y(n_4205)
);

NAND2xp5_ASAP7_75t_L g4206 ( 
.A(n_4175),
.B(n_3918),
.Y(n_4206)
);

AOI221xp5_ASAP7_75t_L g4207 ( 
.A1(n_4175),
.A2(n_3995),
.B1(n_4013),
.B2(n_3923),
.C(n_3919),
.Y(n_4207)
);

NOR3xp33_ASAP7_75t_L g4208 ( 
.A(n_4185),
.B(n_4033),
.C(n_3930),
.Y(n_4208)
);

OAI21xp5_ASAP7_75t_L g4209 ( 
.A1(n_4186),
.A2(n_4041),
.B(n_4029),
.Y(n_4209)
);

AOI222xp33_ASAP7_75t_L g4210 ( 
.A1(n_4207),
.A2(n_4045),
.B1(n_4057),
.B2(n_4056),
.C1(n_4054),
.C2(n_4029),
.Y(n_4210)
);

NAND3xp33_ASAP7_75t_L g4211 ( 
.A(n_4182),
.B(n_4039),
.C(n_4034),
.Y(n_4211)
);

AOI21xp5_ASAP7_75t_L g4212 ( 
.A1(n_4197),
.A2(n_4007),
.B(n_4001),
.Y(n_4212)
);

AOI221xp5_ASAP7_75t_L g4213 ( 
.A1(n_4200),
.A2(n_3919),
.B1(n_3923),
.B2(n_3928),
.C(n_4001),
.Y(n_4213)
);

NAND4xp25_ASAP7_75t_L g4214 ( 
.A(n_4191),
.B(n_4018),
.C(n_3924),
.D(n_4039),
.Y(n_4214)
);

AOI21xp33_ASAP7_75t_SL g4215 ( 
.A1(n_4198),
.A2(n_3949),
.B(n_4050),
.Y(n_4215)
);

AOI21xp5_ASAP7_75t_L g4216 ( 
.A1(n_4184),
.A2(n_4206),
.B(n_4192),
.Y(n_4216)
);

OAI22xp33_ASAP7_75t_L g4217 ( 
.A1(n_4190),
.A2(n_4012),
.B1(n_4007),
.B2(n_3940),
.Y(n_4217)
);

AOI21xp33_ASAP7_75t_L g4218 ( 
.A1(n_4187),
.A2(n_4061),
.B(n_4050),
.Y(n_4218)
);

AOI221xp5_ASAP7_75t_L g4219 ( 
.A1(n_4199),
.A2(n_3928),
.B1(n_4012),
.B2(n_4039),
.C(n_4034),
.Y(n_4219)
);

NOR2xp33_ASAP7_75t_L g4220 ( 
.A(n_4189),
.B(n_4050),
.Y(n_4220)
);

AOI221xp5_ASAP7_75t_L g4221 ( 
.A1(n_4205),
.A2(n_4061),
.B1(n_3931),
.B2(n_3958),
.C(n_3969),
.Y(n_4221)
);

AOI21xp5_ASAP7_75t_L g4222 ( 
.A1(n_4183),
.A2(n_4033),
.B(n_4061),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_L g4223 ( 
.A(n_4195),
.B(n_3931),
.Y(n_4223)
);

OAI221xp5_ASAP7_75t_SL g4224 ( 
.A1(n_4202),
.A2(n_3933),
.B1(n_3940),
.B2(n_3956),
.C(n_3944),
.Y(n_4224)
);

OAI21xp5_ASAP7_75t_L g4225 ( 
.A1(n_4188),
.A2(n_4203),
.B(n_4196),
.Y(n_4225)
);

OR2x2_ASAP7_75t_L g4226 ( 
.A(n_4201),
.B(n_3937),
.Y(n_4226)
);

NOR2xp33_ASAP7_75t_L g4227 ( 
.A(n_4193),
.B(n_3968),
.Y(n_4227)
);

NOR3xp33_ASAP7_75t_L g4228 ( 
.A(n_4194),
.B(n_4204),
.C(n_3924),
.Y(n_4228)
);

NOR2xp33_ASAP7_75t_L g4229 ( 
.A(n_4197),
.B(n_3968),
.Y(n_4229)
);

NAND2xp33_ASAP7_75t_SL g4230 ( 
.A(n_4196),
.B(n_3945),
.Y(n_4230)
);

OAI311xp33_ASAP7_75t_L g4231 ( 
.A1(n_4201),
.A2(n_3955),
.A3(n_3961),
.B1(n_3959),
.C1(n_3965),
.Y(n_4231)
);

NOR2xp33_ASAP7_75t_L g4232 ( 
.A(n_4224),
.B(n_3968),
.Y(n_4232)
);

OAI21xp33_ASAP7_75t_L g4233 ( 
.A1(n_4225),
.A2(n_3945),
.B(n_3939),
.Y(n_4233)
);

AOI22xp5_ASAP7_75t_SL g4234 ( 
.A1(n_4229),
.A2(n_3917),
.B1(n_3924),
.B2(n_3940),
.Y(n_4234)
);

NAND2xp5_ASAP7_75t_L g4235 ( 
.A(n_4215),
.B(n_3931),
.Y(n_4235)
);

AOI22xp5_ASAP7_75t_L g4236 ( 
.A1(n_4211),
.A2(n_3931),
.B1(n_3933),
.B2(n_3945),
.Y(n_4236)
);

AOI21xp5_ASAP7_75t_L g4237 ( 
.A1(n_4230),
.A2(n_3858),
.B(n_3958),
.Y(n_4237)
);

AOI21xp5_ASAP7_75t_L g4238 ( 
.A1(n_4218),
.A2(n_3964),
.B(n_3958),
.Y(n_4238)
);

NAND2xp33_ASAP7_75t_L g4239 ( 
.A(n_4208),
.B(n_3945),
.Y(n_4239)
);

AOI22xp5_ASAP7_75t_L g4240 ( 
.A1(n_4213),
.A2(n_3933),
.B1(n_3945),
.B2(n_3925),
.Y(n_4240)
);

O2A1O1Ixp33_ASAP7_75t_L g4241 ( 
.A1(n_4209),
.A2(n_3925),
.B(n_3986),
.C(n_3964),
.Y(n_4241)
);

NAND4xp25_ASAP7_75t_SL g4242 ( 
.A(n_4222),
.B(n_3861),
.C(n_3895),
.D(n_3905),
.Y(n_4242)
);

AOI211xp5_ASAP7_75t_L g4243 ( 
.A1(n_4231),
.A2(n_3945),
.B(n_3925),
.C(n_4019),
.Y(n_4243)
);

AOI221xp5_ASAP7_75t_L g4244 ( 
.A1(n_4214),
.A2(n_3958),
.B1(n_3969),
.B2(n_3964),
.C(n_3925),
.Y(n_4244)
);

OAI221xp5_ASAP7_75t_L g4245 ( 
.A1(n_4221),
.A2(n_3986),
.B1(n_4016),
.B2(n_3910),
.C(n_3853),
.Y(n_4245)
);

NAND3xp33_ASAP7_75t_L g4246 ( 
.A(n_4216),
.B(n_3964),
.C(n_3969),
.Y(n_4246)
);

NOR3xp33_ASAP7_75t_L g4247 ( 
.A(n_4220),
.B(n_3910),
.C(n_3969),
.Y(n_4247)
);

AOI211xp5_ASAP7_75t_L g4248 ( 
.A1(n_4217),
.A2(n_3944),
.B(n_3961),
.C(n_3966),
.Y(n_4248)
);

AOI21xp33_ASAP7_75t_L g4249 ( 
.A1(n_4235),
.A2(n_4223),
.B(n_4226),
.Y(n_4249)
);

AOI211xp5_ASAP7_75t_L g4250 ( 
.A1(n_4233),
.A2(n_4227),
.B(n_4212),
.C(n_4228),
.Y(n_4250)
);

NAND4xp25_ASAP7_75t_L g4251 ( 
.A(n_4246),
.B(n_4210),
.C(n_4219),
.D(n_3944),
.Y(n_4251)
);

NAND4xp25_ASAP7_75t_L g4252 ( 
.A(n_4232),
.B(n_3892),
.C(n_3966),
.D(n_3965),
.Y(n_4252)
);

NOR3xp33_ASAP7_75t_L g4253 ( 
.A(n_4239),
.B(n_3961),
.C(n_3959),
.Y(n_4253)
);

NAND3xp33_ASAP7_75t_SL g4254 ( 
.A(n_4243),
.B(n_3966),
.C(n_3965),
.Y(n_4254)
);

OAI21xp33_ASAP7_75t_L g4255 ( 
.A1(n_4242),
.A2(n_3986),
.B(n_3904),
.Y(n_4255)
);

AND2x2_ASAP7_75t_SL g4256 ( 
.A(n_4247),
.B(n_3951),
.Y(n_4256)
);

NAND2xp5_ASAP7_75t_L g4257 ( 
.A(n_4237),
.B(n_3959),
.Y(n_4257)
);

AOI22xp5_ASAP7_75t_L g4258 ( 
.A1(n_4244),
.A2(n_3880),
.B1(n_3951),
.B2(n_3915),
.Y(n_4258)
);

NOR3xp33_ASAP7_75t_SL g4259 ( 
.A(n_4245),
.B(n_3955),
.C(n_3886),
.Y(n_4259)
);

NAND5xp2_ASAP7_75t_L g4260 ( 
.A(n_4241),
.B(n_3955),
.C(n_3895),
.D(n_3783),
.E(n_3805),
.Y(n_4260)
);

NOR3x1_ASAP7_75t_L g4261 ( 
.A(n_4234),
.B(n_3857),
.C(n_3847),
.Y(n_4261)
);

OR2x2_ASAP7_75t_L g4262 ( 
.A(n_4236),
.B(n_3947),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_4248),
.Y(n_4263)
);

OAI211xp5_ASAP7_75t_SL g4264 ( 
.A1(n_4249),
.A2(n_4250),
.B(n_4263),
.C(n_4240),
.Y(n_4264)
);

NOR3xp33_ASAP7_75t_L g4265 ( 
.A(n_4251),
.B(n_4238),
.C(n_3957),
.Y(n_4265)
);

NAND4xp25_ASAP7_75t_L g4266 ( 
.A(n_4260),
.B(n_3957),
.C(n_3954),
.D(n_3953),
.Y(n_4266)
);

AOI21xp5_ASAP7_75t_L g4267 ( 
.A1(n_4257),
.A2(n_3957),
.B(n_3954),
.Y(n_4267)
);

AOI21xp33_ASAP7_75t_L g4268 ( 
.A1(n_4262),
.A2(n_3957),
.B(n_3954),
.Y(n_4268)
);

AOI21xp5_ASAP7_75t_L g4269 ( 
.A1(n_4256),
.A2(n_3954),
.B(n_3953),
.Y(n_4269)
);

NAND4xp25_ASAP7_75t_L g4270 ( 
.A(n_4261),
.B(n_3953),
.C(n_3947),
.D(n_3950),
.Y(n_4270)
);

NAND5xp2_ASAP7_75t_L g4271 ( 
.A(n_4255),
.B(n_3880),
.C(n_3950),
.D(n_3947),
.E(n_3953),
.Y(n_4271)
);

AOI211xp5_ASAP7_75t_SL g4272 ( 
.A1(n_4254),
.A2(n_4258),
.B(n_4253),
.C(n_3951),
.Y(n_4272)
);

NAND4xp25_ASAP7_75t_L g4273 ( 
.A(n_4252),
.B(n_3950),
.C(n_3947),
.D(n_3915),
.Y(n_4273)
);

OR2x2_ASAP7_75t_L g4274 ( 
.A(n_4259),
.B(n_3950),
.Y(n_4274)
);

HB1xp67_ASAP7_75t_L g4275 ( 
.A(n_4262),
.Y(n_4275)
);

NOR3xp33_ASAP7_75t_L g4276 ( 
.A(n_4249),
.B(n_3810),
.C(n_3890),
.Y(n_4276)
);

NOR2x1_ASAP7_75t_L g4277 ( 
.A(n_4251),
.B(n_3890),
.Y(n_4277)
);

NAND4xp75_ASAP7_75t_L g4278 ( 
.A(n_4249),
.B(n_3880),
.C(n_3757),
.D(n_3873),
.Y(n_4278)
);

OAI22xp5_ASAP7_75t_L g4279 ( 
.A1(n_4258),
.A2(n_3890),
.B1(n_3951),
.B2(n_3857),
.Y(n_4279)
);

OAI211xp5_ASAP7_75t_SL g4280 ( 
.A1(n_4249),
.A2(n_3847),
.B(n_3872),
.C(n_3856),
.Y(n_4280)
);

NOR3xp33_ASAP7_75t_L g4281 ( 
.A(n_4249),
.B(n_3810),
.C(n_3951),
.Y(n_4281)
);

OAI211xp5_ASAP7_75t_L g4282 ( 
.A1(n_4275),
.A2(n_3880),
.B(n_3902),
.C(n_3822),
.Y(n_4282)
);

NOR2x1_ASAP7_75t_L g4283 ( 
.A(n_4264),
.B(n_4274),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_4270),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_4277),
.Y(n_4285)
);

NAND5xp2_ASAP7_75t_L g4286 ( 
.A(n_4281),
.B(n_3839),
.C(n_3845),
.D(n_3872),
.E(n_3850),
.Y(n_4286)
);

AOI221xp5_ASAP7_75t_L g4287 ( 
.A1(n_4268),
.A2(n_3951),
.B1(n_3853),
.B2(n_3904),
.C(n_3908),
.Y(n_4287)
);

NOR2x1_ASAP7_75t_L g4288 ( 
.A(n_4266),
.B(n_3750),
.Y(n_4288)
);

OA22x2_ASAP7_75t_L g4289 ( 
.A1(n_4279),
.A2(n_4271),
.B1(n_4272),
.B2(n_4276),
.Y(n_4289)
);

INVxp67_ASAP7_75t_L g4290 ( 
.A(n_4265),
.Y(n_4290)
);

AND2x2_ASAP7_75t_L g4291 ( 
.A(n_4269),
.B(n_3839),
.Y(n_4291)
);

AND2x2_ASAP7_75t_L g4292 ( 
.A(n_4278),
.B(n_3845),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_4273),
.Y(n_4293)
);

INVx1_ASAP7_75t_L g4294 ( 
.A(n_4267),
.Y(n_4294)
);

AND2x2_ASAP7_75t_L g4295 ( 
.A(n_4280),
.B(n_3908),
.Y(n_4295)
);

AND2x4_ASAP7_75t_L g4296 ( 
.A(n_4281),
.B(n_3811),
.Y(n_4296)
);

INVx1_ASAP7_75t_L g4297 ( 
.A(n_4275),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_4275),
.Y(n_4298)
);

NAND5xp2_ASAP7_75t_L g4299 ( 
.A(n_4297),
.B(n_3850),
.C(n_3851),
.D(n_3856),
.E(n_3853),
.Y(n_4299)
);

NOR2x1_ASAP7_75t_L g4300 ( 
.A(n_4298),
.B(n_3811),
.Y(n_4300)
);

NAND3xp33_ASAP7_75t_SL g4301 ( 
.A(n_4285),
.B(n_3913),
.C(n_3914),
.Y(n_4301)
);

NOR3xp33_ASAP7_75t_L g4302 ( 
.A(n_4283),
.B(n_3751),
.C(n_3818),
.Y(n_4302)
);

OR2x2_ASAP7_75t_L g4303 ( 
.A(n_4286),
.B(n_3851),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_4291),
.Y(n_4304)
);

NOR2x1_ASAP7_75t_L g4305 ( 
.A(n_4294),
.B(n_3818),
.Y(n_4305)
);

NAND3xp33_ASAP7_75t_L g4306 ( 
.A(n_4290),
.B(n_3822),
.C(n_3824),
.Y(n_4306)
);

AO211x2_ASAP7_75t_L g4307 ( 
.A1(n_4284),
.A2(n_3835),
.B(n_3844),
.C(n_3916),
.Y(n_4307)
);

OAI211xp5_ASAP7_75t_L g4308 ( 
.A1(n_4293),
.A2(n_3820),
.B(n_3824),
.C(n_3914),
.Y(n_4308)
);

NAND2xp5_ASAP7_75t_L g4309 ( 
.A(n_4292),
.B(n_3776),
.Y(n_4309)
);

NOR3xp33_ASAP7_75t_L g4310 ( 
.A(n_4304),
.B(n_4288),
.C(n_4295),
.Y(n_4310)
);

NOR3xp33_ASAP7_75t_L g4311 ( 
.A(n_4300),
.B(n_4296),
.C(n_4282),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_4309),
.Y(n_4312)
);

NOR2x1_ASAP7_75t_L g4313 ( 
.A(n_4305),
.B(n_4289),
.Y(n_4313)
);

NOR3xp33_ASAP7_75t_L g4314 ( 
.A(n_4301),
.B(n_4287),
.C(n_3820),
.Y(n_4314)
);

AOI221xp5_ASAP7_75t_L g4315 ( 
.A1(n_4302),
.A2(n_3835),
.B1(n_3844),
.B2(n_3774),
.C(n_3913),
.Y(n_4315)
);

CKINVDCx6p67_ASAP7_75t_R g4316 ( 
.A(n_4312),
.Y(n_4316)
);

INVx3_ASAP7_75t_L g4317 ( 
.A(n_4313),
.Y(n_4317)
);

INVx2_ASAP7_75t_SL g4318 ( 
.A(n_4311),
.Y(n_4318)
);

INVx1_ASAP7_75t_L g4319 ( 
.A(n_4317),
.Y(n_4319)
);

INVx1_ASAP7_75t_L g4320 ( 
.A(n_4316),
.Y(n_4320)
);

INVx2_ASAP7_75t_L g4321 ( 
.A(n_4319),
.Y(n_4321)
);

INVx1_ASAP7_75t_L g4322 ( 
.A(n_4321),
.Y(n_4322)
);

INVx1_ASAP7_75t_L g4323 ( 
.A(n_4322),
.Y(n_4323)
);

NAND3xp33_ASAP7_75t_L g4324 ( 
.A(n_4323),
.B(n_4320),
.C(n_4310),
.Y(n_4324)
);

OAI22x1_ASAP7_75t_L g4325 ( 
.A1(n_4324),
.A2(n_4318),
.B1(n_4303),
.B2(n_4306),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4325),
.Y(n_4326)
);

AOI21xp5_ASAP7_75t_L g4327 ( 
.A1(n_4326),
.A2(n_4314),
.B(n_4307),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_4327),
.Y(n_4328)
);

OAI21xp5_ASAP7_75t_L g4329 ( 
.A1(n_4328),
.A2(n_4308),
.B(n_4315),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_4329),
.Y(n_4330)
);

OR2x2_ASAP7_75t_L g4331 ( 
.A(n_4330),
.B(n_4299),
.Y(n_4331)
);

AOI221xp5_ASAP7_75t_L g4332 ( 
.A1(n_4331),
.A2(n_3776),
.B1(n_3774),
.B2(n_3753),
.C(n_3876),
.Y(n_4332)
);

AOI221xp5_ASAP7_75t_L g4333 ( 
.A1(n_4331),
.A2(n_3753),
.B1(n_3887),
.B2(n_3876),
.C(n_3916),
.Y(n_4333)
);

AOI22xp5_ASAP7_75t_L g4334 ( 
.A1(n_4333),
.A2(n_3780),
.B1(n_3834),
.B2(n_3762),
.Y(n_4334)
);

AOI211xp5_ASAP7_75t_L g4335 ( 
.A1(n_4334),
.A2(n_4332),
.B(n_3887),
.C(n_3894),
.Y(n_4335)
);


endmodule