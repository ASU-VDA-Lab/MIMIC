module fake_jpeg_24570_n_44 (n_3, n_2, n_1, n_0, n_4, n_5, n_44);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_5),
.B(n_0),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_17),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_15),
.A2(n_20),
.B1(n_8),
.B2(n_9),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_16),
.A2(n_10),
.B1(n_12),
.B2(n_20),
.Y(n_27)
);

BUFx4f_ASAP7_75t_SL g17 ( 
.A(n_11),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_2),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_18),
.B(n_21),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_6),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_6),
.B(n_1),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_27),
.B1(n_28),
.B2(n_22),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_8),
.C(n_9),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_26),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_21),
.A2(n_9),
.B(n_10),
.Y(n_26)
);

NOR3xp33_ASAP7_75t_SL g30 ( 
.A(n_26),
.B(n_17),
.C(n_18),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_24),
.A2(n_17),
.B1(n_19),
.B2(n_12),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_33),
.B1(n_34),
.B2(n_30),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_25),
.A2(n_17),
.B1(n_19),
.B2(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_36),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_33),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_22),
.C(n_28),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_35),
.A2(n_29),
.B1(n_31),
.B2(n_38),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_37),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_43),
.B(n_39),
.Y(n_44)
);


endmodule