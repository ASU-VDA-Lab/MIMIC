module fake_jpeg_31544_n_342 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_51),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_52),
.Y(n_57)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx5_ASAP7_75t_SL g67 ( 
.A(n_49),
.Y(n_67)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_22),
.B(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_30),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_22),
.B(n_1),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_54),
.B(n_23),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_55),
.B(n_63),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_58),
.B(n_62),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_44),
.B(n_27),
.Y(n_63)
);

OR2x2_ASAP7_75t_SL g65 ( 
.A(n_40),
.B(n_24),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_71),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_20),
.B1(n_24),
.B2(n_38),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_66),
.A2(n_29),
.B1(n_32),
.B2(n_31),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_20),
.B1(n_24),
.B2(n_38),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_69),
.A2(n_35),
.B1(n_2),
.B2(n_3),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_43),
.Y(n_71)
);

OR2x2_ASAP7_75t_SL g72 ( 
.A(n_53),
.B(n_28),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_75),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_28),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_78),
.Y(n_104)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_47),
.A2(n_25),
.B1(n_23),
.B2(n_37),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_27),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_77),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_25),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_41),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_17),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_81),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_41),
.Y(n_82)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_41),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_91),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_37),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_84),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_49),
.A2(n_17),
.B1(n_34),
.B2(n_33),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g113 ( 
.A1(n_85),
.A2(n_35),
.B1(n_32),
.B2(n_29),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_26),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_44),
.B(n_34),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_51),
.B(n_33),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_94),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_51),
.B(n_26),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_95),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_96),
.Y(n_142)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_61),
.A2(n_19),
.B1(n_32),
.B2(n_31),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_61),
.A2(n_35),
.B1(n_32),
.B2(n_31),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_106),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_107),
.A2(n_129),
.B1(n_131),
.B2(n_132),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_69),
.A2(n_64),
.B1(n_86),
.B2(n_92),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_110),
.A2(n_114),
.B1(n_130),
.B2(n_71),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_126),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_68),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_64),
.A2(n_35),
.B1(n_2),
.B2(n_3),
.Y(n_114)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_118),
.Y(n_167)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_67),
.Y(n_127)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_80),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_L g131 ( 
.A1(n_73),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_91),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_59),
.C(n_65),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_133),
.B(n_134),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_109),
.B(n_59),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_135),
.B(n_136),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_59),
.C(n_72),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_128),
.B(n_94),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_138),
.B(n_117),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_55),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_143),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_78),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_100),
.B(n_89),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_144),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_146),
.A2(n_153),
.B1(n_163),
.B2(n_157),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_121),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_155),
.Y(n_169)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_103),
.B(n_83),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_157),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_103),
.B(n_79),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_152),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_93),
.B1(n_80),
.B2(n_67),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_154),
.A2(n_119),
.B1(n_87),
.B2(n_68),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_120),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_98),
.B(n_82),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_97),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_159),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_124),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_115),
.B(n_60),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_101),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_112),
.A2(n_93),
.B1(n_80),
.B2(n_56),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_103),
.B(n_87),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_165),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_98),
.B(n_113),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_98),
.A2(n_70),
.B1(n_90),
.B2(n_87),
.Y(n_166)
);

NOR2x1_ASAP7_75t_R g181 ( 
.A(n_166),
.B(n_113),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_143),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_173),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_137),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_175),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_161),
.A2(n_96),
.B1(n_108),
.B2(n_99),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_176),
.A2(n_203),
.B(n_8),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_161),
.A2(n_127),
.B1(n_122),
.B2(n_70),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_177),
.A2(n_181),
.B(n_194),
.Y(n_225)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_183),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_137),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_184),
.Y(n_221)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_186),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_141),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_188),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_189),
.B(n_195),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_190),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_168),
.A2(n_113),
.B1(n_131),
.B2(n_107),
.Y(n_192)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_192),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_145),
.A2(n_142),
.B1(n_122),
.B2(n_166),
.Y(n_194)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_197),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_142),
.B(n_140),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_198),
.B(n_202),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_153),
.A2(n_123),
.B1(n_119),
.B2(n_118),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_199),
.A2(n_164),
.B1(n_168),
.B2(n_149),
.Y(n_212)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_141),
.Y(n_200)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_200),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_133),
.B(n_123),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_152),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_136),
.B(n_8),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_153),
.A2(n_111),
.B1(n_74),
.B2(n_101),
.Y(n_203)
);

AO21x2_ASAP7_75t_L g208 ( 
.A1(n_181),
.A2(n_165),
.B(n_163),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_208),
.A2(n_190),
.B1(n_191),
.B2(n_199),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_211),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_170),
.B(n_150),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_213),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_170),
.B(n_139),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_157),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_215),
.C(n_216),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_146),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_149),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_111),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_219),
.B(n_203),
.C(n_186),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_226),
.B(n_230),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_173),
.B(n_8),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_232),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_178),
.B(n_10),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_171),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_182),
.Y(n_230)
);

AND2x6_ASAP7_75t_L g231 ( 
.A(n_176),
.B(n_15),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_231),
.A2(n_189),
.B(n_202),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_179),
.B(n_10),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_204),
.Y(n_234)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_234),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_235),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_227),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_244),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_220),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_197),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_207),
.A2(n_191),
.B(n_179),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_243),
.A2(n_254),
.B(n_208),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_227),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_206),
.B(n_169),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_245),
.B(n_246),
.Y(n_261)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_233),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_247),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_172),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_248),
.B(n_250),
.Y(n_266)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_249),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_205),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_217),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_251),
.B(n_252),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_221),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_219),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_207),
.A2(n_172),
.B(n_171),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_214),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_224),
.A2(n_185),
.B1(n_180),
.B2(n_187),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_256),
.A2(n_211),
.B1(n_208),
.B2(n_222),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_209),
.B(n_174),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_215),
.C(n_216),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_250),
.B(n_210),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_260),
.B(n_262),
.Y(n_288)
);

AO22x1_ASAP7_75t_L g262 ( 
.A1(n_235),
.A2(n_208),
.B1(n_226),
.B2(n_213),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_263),
.A2(n_270),
.B1(n_274),
.B2(n_256),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_264),
.B(n_272),
.Y(n_289)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_245),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_269),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_246),
.B(n_232),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_239),
.A2(n_231),
.B1(n_225),
.B2(n_212),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_277),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_237),
.A2(n_243),
.B1(n_254),
.B2(n_249),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_238),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_293),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_279),
.A2(n_281),
.B1(n_276),
.B2(n_262),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_276),
.A2(n_225),
.B1(n_251),
.B2(n_252),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_238),
.C(n_257),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_284),
.C(n_286),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_253),
.C(n_255),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_275),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_285),
.B(n_291),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_266),
.A2(n_237),
.B1(n_248),
.B2(n_236),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_287),
.A2(n_258),
.B1(n_268),
.B2(n_241),
.Y(n_306)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_290),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_229),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_292),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_236),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_268),
.Y(n_294)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_294),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_295),
.B(n_296),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_281),
.A2(n_259),
.B(n_265),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_288),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_265),
.C(n_242),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_308),
.C(n_289),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_283),
.Y(n_299)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_299),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_242),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_303),
.B(n_304),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_280),
.B(n_234),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_306),
.A2(n_244),
.B1(n_240),
.B2(n_308),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_247),
.C(n_218),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_312),
.Y(n_325)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_307),
.Y(n_311)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_311),
.Y(n_322)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_300),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_317),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_299),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_315),
.Y(n_327)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_297),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_319),
.Y(n_321)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_298),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_295),
.C(n_305),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_324),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_303),
.C(n_301),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_301),
.C(n_284),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_326),
.B(n_318),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_331),
.Y(n_334)
);

A2O1A1Ixp33_ASAP7_75t_SL g330 ( 
.A1(n_325),
.A2(n_310),
.B(n_289),
.C(n_315),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_330),
.A2(n_327),
.B1(n_174),
.B2(n_183),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_309),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_321),
.A2(n_312),
.B(n_218),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_332),
.B(n_333),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_322),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_335),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_334),
.A2(n_328),
.B(n_330),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_338),
.Y(n_339)
);

AOI321xp33_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_336),
.A3(n_335),
.B1(n_337),
.B2(n_184),
.C(n_175),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_336),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_341),
.B(n_188),
.Y(n_342)
);


endmodule