module fake_jpeg_4677_n_113 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_113);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_113;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_111;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_100;
wire n_82;
wire n_96;

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_33),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_5),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_12),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_30),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_22),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_13),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_69),
.A2(n_64),
.B1(n_60),
.B2(n_53),
.Y(n_79)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_74),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_47),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_74),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_79),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_78),
.A2(n_67),
.B1(n_57),
.B2(n_54),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_56),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_62),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_51),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_59),
.B1(n_46),
.B2(n_49),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_86),
.B(n_25),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_92),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_88),
.A2(n_94),
.B1(n_0),
.B2(n_1),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_84),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_90),
.Y(n_98)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_51),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_55),
.Y(n_93)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_91),
.A2(n_52),
.B(n_81),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_94),
.B(n_80),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_99),
.A2(n_75),
.B1(n_2),
.B2(n_6),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_100),
.A2(n_101),
.B(n_95),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_98),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_97),
.C(n_66),
.Y(n_104)
);

NOR2x1_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_20),
.Y(n_105)
);

NOR2x1_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_23),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_106),
.A2(n_19),
.B(n_3),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_107),
.A2(n_27),
.B(n_7),
.Y(n_108)
);

AOI322xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_29),
.A3(n_9),
.B1(n_11),
.B2(n_14),
.C1(n_15),
.C2(n_16),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_36),
.B1(n_18),
.B2(n_34),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_110),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_111),
.A2(n_35),
.B1(n_43),
.B2(n_44),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_45),
.Y(n_113)
);


endmodule