module real_jpeg_13911_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_215;
wire n_221;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_225;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_202;
wire n_179;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_2),
.A2(n_63),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_2),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_2),
.A2(n_37),
.B1(n_38),
.B2(n_69),
.Y(n_88)
);

BUFx16f_ASAP7_75t_L g85 ( 
.A(n_3),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_4),
.A2(n_63),
.B1(n_70),
.B2(n_72),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_4),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_4),
.A2(n_37),
.B1(n_38),
.B2(n_72),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_5),
.A2(n_46),
.B1(n_47),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_5),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_57),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_5),
.A2(n_37),
.B1(n_38),
.B2(n_57),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_5),
.A2(n_57),
.B1(n_63),
.B2(n_70),
.Y(n_187)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_7),
.A2(n_37),
.B1(n_38),
.B2(n_41),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_7),
.A2(n_41),
.B1(n_63),
.B2(n_70),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_8),
.A2(n_63),
.B1(n_70),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_8),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_27)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_10),
.A2(n_31),
.B1(n_46),
.B2(n_47),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_10),
.A2(n_31),
.B1(n_37),
.B2(n_38),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_10),
.A2(n_31),
.B1(n_63),
.B2(n_70),
.Y(n_182)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_12),
.Y(n_76)
);

AOI21xp33_ASAP7_75t_L g103 ( 
.A1(n_12),
.A2(n_46),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_12),
.B(n_58),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_L g172 ( 
.A1(n_12),
.A2(n_37),
.B1(n_38),
.B2(n_76),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_12),
.A2(n_38),
.B(n_85),
.C(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_12),
.B(n_42),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_12),
.B(n_67),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_12),
.B(n_98),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_12),
.A2(n_28),
.B(n_32),
.C(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_13),
.A2(n_37),
.B1(n_38),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_13),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_81),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_13),
.A2(n_63),
.B1(n_70),
.B2(n_81),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_48),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_14),
.A2(n_37),
.B1(n_38),
.B2(n_48),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_14),
.A2(n_48),
.B1(n_63),
.B2(n_70),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_15),
.A2(n_63),
.B1(n_70),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_15),
.Y(n_93)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_130),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_129),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_105),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_22),
.B(n_105),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_77),
.C(n_94),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_23),
.B(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_59),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_43),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_25),
.B(n_43),
.C(n_59),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B1(n_39),
.B2(n_42),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_27),
.A2(n_36),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_29),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_28),
.A2(n_29),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_28),
.B(n_52),
.Y(n_74)
);

OAI32xp33_ASAP7_75t_L g150 ( 
.A1(n_28),
.A2(n_34),
.A3(n_37),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

OAI32xp33_ASAP7_75t_L g73 ( 
.A1(n_29),
.A2(n_46),
.A3(n_53),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_29),
.B(n_76),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_32),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_32),
.A2(n_42),
.B1(n_137),
.B2(n_139),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_35),
.B(n_38),
.Y(n_152)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_36),
.A2(n_40),
.B1(n_100),
.B2(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_36),
.A2(n_138),
.B(n_208),
.Y(n_207)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_37),
.A2(n_38),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_49),
.B1(n_55),
.B2(n_58),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_45),
.A2(n_50),
.B1(n_51),
.B2(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_46),
.A2(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_54)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_47),
.B(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_50),
.A2(n_51),
.B1(n_56),
.B2(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_73),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_60),
.A2(n_61),
.B1(n_73),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_62),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_62),
.A2(n_67),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_62),
.A2(n_67),
.B1(n_68),
.B2(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_62),
.A2(n_67),
.B1(n_143),
.B2(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_62),
.A2(n_67),
.B1(n_154),
.B2(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_62),
.A2(n_67),
.B1(n_76),
.B2(n_194),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_62),
.A2(n_67),
.B1(n_187),
.B2(n_194),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_70),
.B1(n_85),
.B2(n_86),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_63),
.B(n_196),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_66),
.A2(n_90),
.B1(n_186),
.B2(n_188),
.Y(n_185)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_L g175 ( 
.A1(n_70),
.A2(n_76),
.B(n_86),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_71),
.Y(n_91)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_73),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_77),
.B(n_94),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_89),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_89),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B1(n_87),
.B2(n_88),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_83),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_82),
.A2(n_87),
.B1(n_146),
.B2(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_83),
.A2(n_98),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_83),
.A2(n_97),
.B1(n_98),
.B2(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_83),
.A2(n_98),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_83),
.A2(n_98),
.B1(n_173),
.B2(n_180),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.C(n_102),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_95),
.A2(n_96),
.B1(n_99),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_102),
.B(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_128),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_117),
.B1(n_126),
.B2(n_127),
.Y(n_106)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_112),
.B2(n_116),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_112),
.Y(n_116)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_226),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_222),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_165),
.B(n_221),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_155),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_134),
.B(n_155),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_144),
.C(n_147),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_135),
.B(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_140),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_141),
.C(n_142),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_144),
.A2(n_147),
.B1(n_148),
.B2(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_144),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_153),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_149),
.A2(n_150),
.B1(n_153),
.B2(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_151),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_153),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_160),
.B2(n_164),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_156),
.B(n_161),
.C(n_163),
.Y(n_223)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_160),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_215),
.B(n_220),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_203),
.B(n_214),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_183),
.B(n_202),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_176),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_169),
.B(n_176),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_174),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_170),
.A2(n_171),
.B1(n_174),
.B2(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_179),
.C(n_181),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_182),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_191),
.B(n_201),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_189),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_185),
.B(n_189),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_197),
.B(n_200),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_198),
.B(n_199),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_204),
.B(n_205),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_212),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_210),
.C(n_212),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_216),
.B(n_217),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_223),
.B(n_224),
.Y(n_226)
);


endmodule