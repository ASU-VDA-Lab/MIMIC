module fake_netlist_6_248_n_3853 (n_52, n_591, n_435, n_1, n_91, n_793, n_326, n_801, n_256, n_440, n_587, n_695, n_507, n_580, n_762, n_209, n_367, n_465, n_680, n_741, n_760, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_740, n_578, n_703, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_783, n_106, n_725, n_358, n_160, n_751, n_449, n_131, n_749, n_798, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_805, n_396, n_495, n_350, n_78, n_84, n_585, n_732, n_568, n_392, n_442, n_480, n_142, n_724, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_698, n_255, n_807, n_739, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_768, n_38, n_471, n_289, n_421, n_781, n_424, n_789, n_615, n_59, n_181, n_182, n_238, n_573, n_769, n_202, n_320, n_108, n_639, n_676, n_327, n_794, n_727, n_369, n_597, n_685, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_747, n_667, n_71, n_74, n_229, n_542, n_644, n_682, n_621, n_305, n_72, n_721, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_791, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_704, n_748, n_506, n_56, n_763, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_710, n_387, n_452, n_616, n_658, n_744, n_39, n_344, n_73, n_581, n_428, n_761, n_785, n_746, n_609, n_765, n_432, n_641, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_758, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_772, n_96, n_8, n_797, n_666, n_371, n_795, n_770, n_567, n_189, n_738, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_752, n_112, n_172, n_713, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_782, n_490, n_803, n_290, n_220, n_809, n_118, n_224, n_48, n_25, n_93, n_80, n_734, n_708, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_779, n_9, n_800, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_366, n_777, n_407, n_450, n_103, n_808, n_272, n_526, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_717, n_46, n_330, n_771, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_686, n_796, n_252, n_757, n_228, n_565, n_594, n_719, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_745, n_654, n_323, n_606, n_393, n_411, n_503, n_716, n_152, n_623, n_92, n_599, n_513, n_776, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_731, n_406, n_483, n_735, n_102, n_204, n_482, n_755, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_792, n_476, n_714, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_788, n_325, n_767, n_804, n_329, n_464, n_600, n_802, n_561, n_33, n_477, n_549, n_533, n_408, n_806, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_345, n_409, n_231, n_354, n_689, n_40, n_799, n_505, n_240, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_810, n_635, n_95, n_787, n_311, n_10, n_403, n_723, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_764, n_556, n_159, n_157, n_162, n_692, n_733, n_754, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_753, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_737, n_318, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_790, n_582, n_4, n_199, n_138, n_266, n_296, n_674, n_775, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_759, n_355, n_426, n_317, n_149, n_632, n_702, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_780, n_773, n_675, n_85, n_99, n_257, n_730, n_655, n_13, n_706, n_786, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_690, n_29, n_75, n_401, n_324, n_743, n_766, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_728, n_681, n_729, n_110, n_151, n_774, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_784, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_688, n_722, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_637, n_295, n_385, n_701, n_629, n_388, n_190, n_262, n_484, n_613, n_736, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_778, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_3853);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_793;
input n_326;
input n_801;
input n_256;
input n_440;
input n_587;
input n_695;
input n_507;
input n_580;
input n_762;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_760;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_740;
input n_578;
input n_703;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_783;
input n_106;
input n_725;
input n_358;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_798;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_805;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_732;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_724;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_255;
input n_807;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_768;
input n_38;
input n_471;
input n_289;
input n_421;
input n_781;
input n_424;
input n_789;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_769;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_794;
input n_727;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_747;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_682;
input n_621;
input n_305;
input n_72;
input n_721;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_791;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_704;
input n_748;
input n_506;
input n_56;
input n_763;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_387;
input n_452;
input n_616;
input n_658;
input n_744;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_761;
input n_785;
input n_746;
input n_609;
input n_765;
input n_432;
input n_641;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_758;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_772;
input n_96;
input n_8;
input n_797;
input n_666;
input n_371;
input n_795;
input n_770;
input n_567;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_752;
input n_112;
input n_172;
input n_713;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_782;
input n_490;
input n_803;
input n_290;
input n_220;
input n_809;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_734;
input n_708;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_779;
input n_9;
input n_800;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_366;
input n_777;
input n_407;
input n_450;
input n_103;
input n_808;
input n_272;
input n_526;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_717;
input n_46;
input n_330;
input n_771;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_686;
input n_796;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_745;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_716;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_776;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_731;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_755;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_792;
input n_476;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_788;
input n_325;
input n_767;
input n_804;
input n_329;
input n_464;
input n_600;
input n_802;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_806;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_799;
input n_505;
input n_240;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_810;
input n_635;
input n_95;
input n_787;
input n_311;
input n_10;
input n_403;
input n_723;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_764;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_733;
input n_754;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_753;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_790;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_674;
input n_775;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_759;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_780;
input n_773;
input n_675;
input n_85;
input n_99;
input n_257;
input n_730;
input n_655;
input n_13;
input n_706;
input n_786;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_690;
input n_29;
input n_75;
input n_401;
input n_324;
input n_743;
input n_766;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_728;
input n_681;
input n_729;
input n_110;
input n_151;
input n_774;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_784;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_688;
input n_722;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_637;
input n_295;
input n_385;
input n_701;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_778;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_3853;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_3813;
wire n_3766;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_3254;
wire n_3684;
wire n_1199;
wire n_1674;
wire n_3392;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_1189;
wire n_3152;
wire n_3579;
wire n_1212;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3783;
wire n_3773;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_3849;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_3844;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_1357;
wire n_1853;
wire n_3741;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_1342;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_1708;
wire n_1151;
wire n_2977;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_3332;
wire n_3465;
wire n_1975;
wire n_1930;
wire n_1743;
wire n_1009;
wire n_2405;
wire n_3706;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_1724;
wire n_1032;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_1264;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_3619;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_2291;
wire n_830;
wire n_2299;
wire n_3340;
wire n_1371;
wire n_873;
wire n_1285;
wire n_2886;
wire n_2974;
wire n_1985;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3626;
wire n_3757;
wire n_1393;
wire n_1867;
wire n_1517;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_3106;
wire n_2630;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_836;
wire n_3345;
wire n_2074;
wire n_2447;
wire n_2919;
wire n_3678;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_2356;
wire n_1143;
wire n_2399;
wire n_1422;
wire n_1772;
wire n_1232;
wire n_1572;
wire n_1874;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_2480;
wire n_1300;
wire n_2739;
wire n_3023;
wire n_822;
wire n_3232;
wire n_2791;
wire n_1313;
wire n_3750;
wire n_3607;
wire n_3251;
wire n_1056;
wire n_3316;
wire n_2212;
wire n_3494;
wire n_3048;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3063;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_940;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_3028;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3624;
wire n_3077;
wire n_3737;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3452;
wire n_3655;
wire n_3107;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_3765;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_1467;
wire n_3297;
wire n_976;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3368;
wire n_917;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_907;
wire n_1446;
wire n_2591;
wire n_3507;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_913;
wire n_1658;
wire n_2593;
wire n_867;
wire n_3506;
wire n_3568;
wire n_3269;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_3850;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_1986;
wire n_2397;
wire n_824;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_2907;
wire n_3438;
wire n_2735;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_2850;
wire n_1909;
wire n_813;
wire n_2080;
wire n_1481;
wire n_3822;
wire n_1441;
wire n_818;
wire n_3373;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_1381;
wire n_2961;
wire n_3812;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_2669;
wire n_2925;
wire n_3728;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_2522;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_3798;
wire n_939;
wire n_3488;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_3732;
wire n_982;
wire n_2674;
wire n_2832;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_2831;
wire n_2998;
wire n_3446;
wire n_3317;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_3716;
wire n_1873;
wire n_905;
wire n_3630;
wire n_3518;
wire n_3824;
wire n_1866;
wire n_1680;
wire n_2692;
wire n_993;
wire n_3842;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1605;
wire n_1413;
wire n_1330;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_2355;
wire n_966;
wire n_2908;
wire n_3168;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_3403;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_3055;
wire n_3092;
wire n_3492;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_3294;
wire n_1014;
wire n_3734;
wire n_3686;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_882;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_3746;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_1265;
wire n_2711;
wire n_3490;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_3369;
wire n_3419;
wire n_1982;
wire n_2878;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3772;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_3794;
wire n_3247;
wire n_871;
wire n_3069;
wire n_922;
wire n_1760;
wire n_1335;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_1722;
wire n_1664;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_2749;
wire n_2008;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2254;
wire n_2345;
wire n_3346;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_3691;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_1801;
wire n_1214;
wire n_835;
wire n_850;
wire n_928;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3428;
wire n_3153;
wire n_3410;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_825;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_1588;
wire n_3785;
wire n_2963;
wire n_2947;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_1624;
wire n_1124;
wire n_2096;
wire n_2980;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_3434;
wire n_1515;
wire n_961;
wire n_3510;
wire n_1317;
wire n_1082;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_890;
wire n_2377;
wire n_3271;
wire n_2178;
wire n_950;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_3526;
wire n_3707;
wire n_2075;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_3545;
wire n_968;
wire n_909;
wire n_1369;
wire n_3578;
wire n_881;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_3073;
wire n_2431;
wire n_2987;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_3696;
wire n_3780;
wire n_2078;
wire n_1634;
wire n_3252;
wire n_2932;
wire n_1767;
wire n_3253;
wire n_1779;
wire n_1465;
wire n_3337;
wire n_3431;
wire n_3450;
wire n_3209;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2893;
wire n_2775;
wire n_1208;
wire n_1627;
wire n_1295;
wire n_1164;
wire n_2954;
wire n_3477;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_3421;
wire n_840;
wire n_2913;
wire n_3614;
wire n_874;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1565;
wire n_1067;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_3616;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_3436;
wire n_1932;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_3366;
wire n_3442;
wire n_2631;
wire n_1364;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_963;
wire n_2767;
wire n_3793;
wire n_894;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_1514;
wire n_1863;
wire n_826;
wire n_3385;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_872;
wire n_1714;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_2897;
wire n_847;
wire n_851;
wire n_2537;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_1513;
wire n_2747;
wire n_3171;
wire n_1913;
wire n_3608;
wire n_837;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_3491;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_3158;
wire n_1788;
wire n_3426;
wire n_1999;
wire n_2731;
wire n_2643;
wire n_2590;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_3782;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_3470;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_1492;
wire n_987;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_3104;
wire n_3435;
wire n_842;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_3611;
wire n_1432;
wire n_2208;
wire n_843;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_899;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_3580;
wire n_3775;
wire n_3537;
wire n_1004;
wire n_2134;
wire n_1176;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_3835;
wire n_1809;
wire n_3119;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_947;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1448;
wire n_1087;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_1049;
wire n_3223;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_3770;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_1849;
wire n_2848;
wire n_919;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_2231;
wire n_3609;
wire n_929;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_3693;
wire n_3788;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_1299;
wire n_2896;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_2368;
wire n_2403;
wire n_1070;
wire n_3342;
wire n_2837;
wire n_998;
wire n_3200;
wire n_1665;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_3390;
wire n_3656;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_3324;
wire n_3593;
wire n_3341;
wire n_1073;
wire n_1000;
wire n_1195;
wire n_3559;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_1507;
wire n_2482;
wire n_3810;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_2481;
wire n_3561;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_2424;
wire n_1604;
wire n_2296;
wire n_1284;
wire n_3201;
wire n_3633;
wire n_3447;
wire n_1142;
wire n_2849;
wire n_1475;
wire n_1774;
wire n_1398;
wire n_2354;
wire n_884;
wire n_1048;
wire n_2682;
wire n_1201;
wire n_3032;
wire n_3103;
wire n_3638;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_1021;
wire n_931;
wire n_3393;
wire n_811;
wire n_1207;
wire n_2442;
wire n_3627;
wire n_1791;
wire n_1368;
wire n_3451;
wire n_3480;
wire n_1418;
wire n_958;
wire n_1250;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3087;
wire n_3072;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_3577;
wire n_3540;
wire n_889;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_819;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_3641;
wire n_3591;
wire n_1837;
wire n_964;
wire n_831;
wire n_2218;
wire n_1314;
wire n_2788;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2860;
wire n_2292;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2511;
wire n_2475;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2323;
wire n_1220;
wire n_1893;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_3582;
wire n_3605;
wire n_3287;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_970;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_3481;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_3033;
wire n_3724;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_2990;
wire n_3847;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_1286;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3226;
wire n_3364;
wire n_3323;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_1153;
wire n_1618;
wire n_3407;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_3425;
wire n_2384;
wire n_1745;
wire n_914;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_3646;
wire n_2920;
wire n_3547;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_3188;
wire n_3742;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_1617;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_3816;
wire n_1470;
wire n_2550;
wire n_3093;
wire n_3175;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_848;
wire n_2732;
wire n_2928;
wire n_2249;
wire n_1096;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_3284;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_3205;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_1390;
wire n_906;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_2863;
wire n_3299;
wire n_3663;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_3360;
wire n_2135;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_2049;
wire n_858;
wire n_1331;
wire n_2627;
wire n_3234;
wire n_956;
wire n_960;
wire n_2276;
wire n_856;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_2993;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3016;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_1129;
wire n_2829;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_3751;
wire n_1869;
wire n_2911;
wire n_3625;
wire n_3804;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_1889;
wire n_2379;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_1635;
wire n_2942;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_2555;
wire n_3338;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_999;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_3722;
wire n_2984;
wire n_994;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2656;
wire n_2278;
wire n_2538;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3250;
wire n_3194;
wire n_1934;
wire n_3276;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_845;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_1510;
wire n_892;
wire n_3637;
wire n_3120;
wire n_1468;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3797;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_3548;
wire n_3767;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_1847;
wire n_2052;
wire n_3634;
wire n_2302;
wire n_1667;
wire n_1206;
wire n_3230;
wire n_1397;
wire n_1037;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_901;
wire n_1499;
wire n_3592;
wire n_2755;
wire n_3141;
wire n_923;
wire n_1409;
wire n_1841;
wire n_3839;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_1818;
wire n_1108;
wire n_2439;
wire n_3730;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_2740;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_3042;
wire n_1356;
wire n_1589;
wire n_3213;
wire n_3820;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1943;
wire n_1216;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3238;
wire n_2235;
wire n_3529;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_3424;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_3784;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_1043;
wire n_3819;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_1870;
wire n_2964;
wire n_1692;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_3485;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3475;
wire n_3501;
wire n_1840;
wire n_1152;
wire n_1705;
wire n_3262;
wire n_3544;
wire n_2904;
wire n_2244;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_3692;
wire n_3845;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_1405;
wire n_972;
wire n_2376;
wire n_3826;
wire n_1406;
wire n_3790;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_962;
wire n_1041;
wire n_2346;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_2882;
wire n_3675;
wire n_3666;
wire n_3320;
wire n_2541;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_3307;
wire n_3439;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_3588;
wire n_2871;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_3502;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_2390;
wire n_3712;
wire n_959;
wire n_879;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_2986;
wire n_1900;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2962;
wire n_2154;
wire n_2727;
wire n_3377;
wire n_2939;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_1914;
wire n_1318;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_3762;
wire n_3469;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_1029;
wire n_3779;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_1706;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_3558;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_3379;
wire n_3156;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_2668;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_1375;
wire n_1941;
wire n_3483;
wire n_3613;
wire n_2128;
wire n_1650;
wire n_1794;
wire n_1962;
wire n_1045;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_3743;
wire n_1872;
wire n_3091;
wire n_834;
wire n_2695;
wire n_3818;
wire n_3124;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_3524;
wire n_2671;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2888;
wire n_1804;
wire n_2923;
wire n_3711;
wire n_3776;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_3511;
wire n_2054;
wire n_876;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_869;
wire n_1154;
wire n_3308;
wire n_1600;
wire n_1113;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_3602;
wire n_897;
wire n_846;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_1476;
wire n_841;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_3777;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_3515;
wire n_1150;
wire n_3808;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1118;
wire n_1076;
wire n_2949;
wire n_3726;
wire n_1807;
wire n_1007;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_3758;
wire n_1879;
wire n_853;
wire n_3806;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_875;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_1953;
wire n_933;
wire n_3343;
wire n_3303;
wire n_978;
wire n_2752;
wire n_3135;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_969;
wire n_2140;
wire n_988;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_3658;
wire n_1516;
wire n_1536;
wire n_3846;
wire n_2163;
wire n_2186;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3034;
wire n_823;
wire n_1132;
wire n_1074;
wire n_1394;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_955;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_2969;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_3027;
wire n_1554;
wire n_3231;
wire n_1130;
wire n_3083;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_2380;
wire n_1120;
wire n_832;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_814;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_3541;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_1461;
wire n_3432;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_1598;
wire n_3493;
wire n_2935;
wire n_3807;
wire n_863;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_918;
wire n_1848;
wire n_1785;
wire n_1114;
wire n_1147;
wire n_3268;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_3701;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_3473;
wire n_895;
wire n_866;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_3739;
wire n_2284;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_971;
wire n_2702;
wire n_3241;
wire n_946;
wire n_2906;
wire n_1303;
wire n_2769;
wire n_3622;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_1245;
wire n_838;
wire n_3215;
wire n_3336;
wire n_844;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_3553;
wire n_1561;
wire n_2741;
wire n_3114;
wire n_930;
wire n_888;
wire n_2275;
wire n_2465;
wire n_1112;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_3811;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_2430;
wire n_3486;
wire n_1414;
wire n_3584;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_3556;
wire n_2034;
wire n_1028;
wire n_3836;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_2437;
wire n_839;
wire n_2743;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_990;
wire n_1500;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_3699;
wire n_3204;
wire n_1104;
wire n_854;
wire n_1058;
wire n_3378;
wire n_2312;
wire n_3404;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_2242;
wire n_3362;
wire n_3745;
wire n_1509;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_3256;
wire n_1276;
wire n_3802;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_3796;
wire n_2999;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3643;
wire n_3697;
wire n_1584;
wire n_2425;
wire n_924;
wire n_3408;
wire n_3461;
wire n_1582;
wire n_3680;
wire n_2318;
wire n_3286;
wire n_2408;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_3098;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_1362;
wire n_829;
wire n_1156;
wire n_3123;
wire n_2600;
wire n_984;
wire n_3380;
wire n_1829;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_868;
wire n_3038;
wire n_859;
wire n_2033;
wire n_3086;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_3285;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_3361;
wire n_981;
wire n_3596;
wire n_3478;
wire n_1349;
wire n_2071;
wire n_1144;
wire n_3669;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_3521;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_1301;
wire n_2805;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_3344;
wire n_2334;
wire n_3295;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_1133;
wire n_1194;
wire n_3374;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_2640;
wire n_3695;
wire n_1051;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_2367;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_941;
wire n_3552;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_849;
wire n_2662;
wire n_3116;
wire n_3147;
wire n_3383;
wire n_3709;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_3187;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_2065;
wire n_2879;
wire n_861;
wire n_3717;
wire n_857;
wire n_967;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_2968;
wire n_1629;
wire n_1170;
wire n_2221;
wire n_1819;
wire n_2055;
wire n_1260;
wire n_3555;
wire n_1010;
wire n_3444;
wire n_2553;
wire n_1040;
wire n_915;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_3833;
wire n_3815;
wire n_2774;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3274;
wire n_3333;
wire n_3186;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_2579;
wire n_862;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_3085;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_3387;
wire n_2027;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_3504;
wire n_1449;
wire n_827;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_1742;
wire n_1612;
wire n_1240;

INVxp67_ASAP7_75t_L g811 ( 
.A(n_222),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_620),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_291),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_464),
.Y(n_814)
);

BUFx10_ASAP7_75t_L g815 ( 
.A(n_441),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_474),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_565),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_714),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_411),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_753),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_528),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_419),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_498),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_349),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_499),
.Y(n_825)
);

BUFx5_ASAP7_75t_L g826 ( 
.A(n_249),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_660),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_160),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_97),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_488),
.Y(n_830)
);

INVxp67_ASAP7_75t_L g831 ( 
.A(n_73),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_734),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_168),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_681),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_355),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_313),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_221),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_663),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_180),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_459),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_214),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_719),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_170),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_547),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_198),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_793),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_58),
.Y(n_847)
);

CKINVDCx20_ASAP7_75t_R g848 ( 
.A(n_303),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_751),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_381),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_727),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_74),
.Y(n_852)
);

BUFx8_ASAP7_75t_SL g853 ( 
.A(n_759),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_762),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_664),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_388),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_627),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_122),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_524),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_324),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_439),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_364),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_13),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_802),
.Y(n_864)
);

CKINVDCx16_ASAP7_75t_R g865 ( 
.A(n_518),
.Y(n_865)
);

BUFx3_ASAP7_75t_L g866 ( 
.A(n_32),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_469),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_647),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_728),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_313),
.Y(n_870)
);

BUFx8_ASAP7_75t_SL g871 ( 
.A(n_158),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_466),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_461),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_670),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_785),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_678),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_578),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_527),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_615),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_672),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_804),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_605),
.Y(n_882)
);

INVx1_ASAP7_75t_SL g883 ( 
.A(n_283),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_748),
.Y(n_884)
);

CKINVDCx20_ASAP7_75t_R g885 ( 
.A(n_96),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_761),
.Y(n_886)
);

INVx1_ASAP7_75t_SL g887 ( 
.A(n_514),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_112),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_84),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_113),
.Y(n_890)
);

CKINVDCx20_ASAP7_75t_R g891 ( 
.A(n_697),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_203),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_406),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_381),
.Y(n_894)
);

INVx1_ASAP7_75t_SL g895 ( 
.A(n_364),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_589),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_221),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_711),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_757),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_480),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_731),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_428),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_790),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_483),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_547),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_613),
.Y(n_906)
);

BUFx10_ASAP7_75t_L g907 ( 
.A(n_100),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_323),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_360),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_532),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_808),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_755),
.Y(n_912)
);

BUFx5_ASAP7_75t_L g913 ( 
.A(n_803),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_752),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_772),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_800),
.Y(n_916)
);

CKINVDCx20_ASAP7_75t_R g917 ( 
.A(n_612),
.Y(n_917)
);

CKINVDCx20_ASAP7_75t_R g918 ( 
.A(n_163),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_8),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_801),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_442),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_664),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_390),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_216),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_708),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_774),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_566),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_527),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_726),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_539),
.Y(n_930)
);

BUFx10_ASAP7_75t_L g931 ( 
.A(n_350),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_94),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_607),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_743),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_787),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_143),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_807),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_330),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_273),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_590),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_725),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_742),
.Y(n_942)
);

CKINVDCx20_ASAP7_75t_R g943 ( 
.A(n_413),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_408),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_454),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_569),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_766),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_105),
.Y(n_948)
);

BUFx8_ASAP7_75t_SL g949 ( 
.A(n_744),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_566),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_443),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_723),
.Y(n_952)
);

INVxp67_ASAP7_75t_L g953 ( 
.A(n_159),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_609),
.Y(n_954)
);

BUFx10_ASAP7_75t_L g955 ( 
.A(n_351),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_559),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_777),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_206),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_754),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_350),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_90),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_20),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_223),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_799),
.Y(n_964)
);

CKINVDCx20_ASAP7_75t_R g965 ( 
.A(n_689),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_95),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_78),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_370),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_349),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_652),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_581),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_695),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_623),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_383),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_285),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_512),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_194),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_190),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_724),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_736),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_558),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_751),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_230),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_358),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_61),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_177),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_567),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_34),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_746),
.Y(n_989)
);

BUFx10_ASAP7_75t_L g990 ( 
.A(n_251),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_806),
.Y(n_991)
);

INVx1_ASAP7_75t_SL g992 ( 
.A(n_715),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_377),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_180),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_610),
.Y(n_995)
);

INVx2_ASAP7_75t_SL g996 ( 
.A(n_747),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_489),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_340),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_618),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_306),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_747),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_792),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_720),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_651),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_472),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_51),
.Y(n_1006)
);

INVx1_ASAP7_75t_SL g1007 ( 
.A(n_728),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_739),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_135),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_407),
.Y(n_1010)
);

CKINVDCx20_ASAP7_75t_R g1011 ( 
.A(n_509),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_150),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_454),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_509),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_732),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_92),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_240),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_398),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_741),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_390),
.Y(n_1020)
);

INVx2_ASAP7_75t_SL g1021 ( 
.A(n_369),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_762),
.Y(n_1022)
);

INVxp33_ASAP7_75t_L g1023 ( 
.A(n_733),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_127),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_0),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_209),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_536),
.Y(n_1027)
);

CKINVDCx14_ASAP7_75t_R g1028 ( 
.A(n_301),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_810),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_469),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_133),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_760),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_19),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_209),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_491),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_120),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_303),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_613),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_156),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_749),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_316),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_694),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_1),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_136),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_265),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_640),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_384),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_654),
.Y(n_1048)
);

INVxp67_ASAP7_75t_L g1049 ( 
.A(n_700),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_434),
.Y(n_1050)
);

CKINVDCx20_ASAP7_75t_R g1051 ( 
.A(n_618),
.Y(n_1051)
);

BUFx10_ASAP7_75t_L g1052 ( 
.A(n_691),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_552),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_351),
.Y(n_1054)
);

BUFx2_ASAP7_75t_L g1055 ( 
.A(n_703),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_773),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_9),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_649),
.Y(n_1058)
);

INVx1_ASAP7_75t_SL g1059 ( 
.A(n_302),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_249),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_182),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_85),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_736),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_705),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_343),
.Y(n_1065)
);

INVx1_ASAP7_75t_SL g1066 ( 
.A(n_577),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_745),
.Y(n_1067)
);

INVx2_ASAP7_75t_SL g1068 ( 
.A(n_451),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_247),
.Y(n_1069)
);

INVx4_ASAP7_75t_R g1070 ( 
.A(n_558),
.Y(n_1070)
);

CKINVDCx14_ASAP7_75t_R g1071 ( 
.A(n_395),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_107),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_763),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_171),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_794),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_93),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_797),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_108),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_721),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_208),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_549),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_621),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_315),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_196),
.Y(n_1084)
);

INVx4_ASAP7_75t_R g1085 ( 
.A(n_149),
.Y(n_1085)
);

INVx2_ASAP7_75t_SL g1086 ( 
.A(n_463),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_329),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_505),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_434),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_665),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_525),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_654),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_809),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_624),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_577),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_31),
.Y(n_1096)
);

CKINVDCx20_ASAP7_75t_R g1097 ( 
.A(n_46),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_118),
.Y(n_1098)
);

BUFx10_ASAP7_75t_L g1099 ( 
.A(n_410),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_494),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_183),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_780),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_498),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_717),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_193),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_635),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_95),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_658),
.Y(n_1108)
);

CKINVDCx20_ASAP7_75t_R g1109 ( 
.A(n_53),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_679),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_623),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_21),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_669),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_683),
.Y(n_1114)
);

CKINVDCx20_ASAP7_75t_R g1115 ( 
.A(n_268),
.Y(n_1115)
);

BUFx3_ASAP7_75t_L g1116 ( 
.A(n_733),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_414),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_380),
.Y(n_1118)
);

INVx2_ASAP7_75t_SL g1119 ( 
.A(n_796),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_805),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_524),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_573),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_200),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_571),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_545),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_104),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_564),
.Y(n_1127)
);

CKINVDCx20_ASAP7_75t_R g1128 ( 
.A(n_484),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_213),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_368),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_110),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_440),
.Y(n_1132)
);

CKINVDCx20_ASAP7_75t_R g1133 ( 
.A(n_489),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_232),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_752),
.Y(n_1135)
);

HB1xp67_ASAP7_75t_L g1136 ( 
.A(n_379),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_517),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_685),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_523),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_205),
.Y(n_1140)
);

CKINVDCx20_ASAP7_75t_R g1141 ( 
.A(n_129),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_370),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_245),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_745),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_101),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_534),
.Y(n_1146)
);

CKINVDCx20_ASAP7_75t_R g1147 ( 
.A(n_49),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_375),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_348),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_256),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_612),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_344),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_76),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_578),
.Y(n_1154)
);

INVx1_ASAP7_75t_SL g1155 ( 
.A(n_714),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_235),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_755),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_360),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_130),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_192),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_325),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_642),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_162),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_111),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_737),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_795),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_471),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_552),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_346),
.Y(n_1169)
);

CKINVDCx20_ASAP7_75t_R g1170 ( 
.A(n_187),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_314),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_590),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_615),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_735),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_735),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_515),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_666),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_185),
.Y(n_1178)
);

BUFx10_ASAP7_75t_L g1179 ( 
.A(n_144),
.Y(n_1179)
);

INVx2_ASAP7_75t_SL g1180 ( 
.A(n_791),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_254),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_41),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_738),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_756),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_143),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_215),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_66),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_147),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_570),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_628),
.Y(n_1190)
);

CKINVDCx14_ASAP7_75t_R g1191 ( 
.A(n_644),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_0),
.Y(n_1192)
);

BUFx3_ASAP7_75t_L g1193 ( 
.A(n_632),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_584),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_16),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_377),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_298),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_798),
.Y(n_1198)
);

CKINVDCx14_ASAP7_75t_R g1199 ( 
.A(n_237),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_412),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_706),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_557),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_242),
.Y(n_1203)
);

CKINVDCx20_ASAP7_75t_R g1204 ( 
.A(n_677),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_79),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_460),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_76),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_500),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_421),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_48),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_681),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_708),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_260),
.Y(n_1213)
);

BUFx8_ASAP7_75t_SL g1214 ( 
.A(n_15),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_482),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_723),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_45),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_263),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_151),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_111),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_241),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_499),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_662),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_179),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_572),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_170),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_621),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_690),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_151),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_101),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_694),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_301),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_148),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_41),
.Y(n_1234)
);

INVx1_ASAP7_75t_SL g1235 ( 
.A(n_281),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_255),
.Y(n_1236)
);

CKINVDCx20_ASAP7_75t_R g1237 ( 
.A(n_376),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_L g1238 ( 
.A(n_444),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_560),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_426),
.Y(n_1240)
);

CKINVDCx20_ASAP7_75t_R g1241 ( 
.A(n_775),
.Y(n_1241)
);

INVx1_ASAP7_75t_SL g1242 ( 
.A(n_490),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_451),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_589),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_81),
.Y(n_1245)
);

INVx1_ASAP7_75t_SL g1246 ( 
.A(n_256),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_20),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_572),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_356),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_759),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_580),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_695),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_296),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_483),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_548),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_27),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_424),
.Y(n_1257)
);

CKINVDCx20_ASAP7_75t_R g1258 ( 
.A(n_112),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_445),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_674),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_624),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_452),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_395),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_740),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_87),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_789),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_375),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_658),
.Y(n_1268)
);

CKINVDCx20_ASAP7_75t_R g1269 ( 
.A(n_579),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_779),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_83),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_705),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_443),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_674),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_373),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_716),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_37),
.Y(n_1277)
);

BUFx8_ASAP7_75t_SL g1278 ( 
.A(n_722),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_753),
.Y(n_1279)
);

BUFx10_ASAP7_75t_L g1280 ( 
.A(n_161),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_515),
.Y(n_1281)
);

INVx1_ASAP7_75t_SL g1282 ( 
.A(n_473),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_446),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_431),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_462),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_253),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_580),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_324),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_98),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_99),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_124),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_441),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_110),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_758),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_478),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_669),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_725),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_437),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_764),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_649),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_667),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_435),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_322),
.Y(n_1303)
);

CKINVDCx20_ASAP7_75t_R g1304 ( 
.A(n_343),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_83),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_18),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_182),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_98),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_357),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_5),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_293),
.Y(n_1311)
);

INVx1_ASAP7_75t_SL g1312 ( 
.A(n_337),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_600),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_168),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_608),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_189),
.Y(n_1316)
);

CKINVDCx16_ASAP7_75t_R g1317 ( 
.A(n_634),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_51),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_460),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_340),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_567),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_732),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_492),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_729),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_153),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_750),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_253),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_730),
.Y(n_1328)
);

BUFx5_ASAP7_75t_L g1329 ( 
.A(n_21),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_28),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_405),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_405),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_357),
.Y(n_1333)
);

BUFx2_ASAP7_75t_L g1334 ( 
.A(n_688),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_322),
.Y(n_1335)
);

CKINVDCx16_ASAP7_75t_R g1336 ( 
.A(n_93),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_503),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_6),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_299),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_616),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_191),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_183),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_703),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_607),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_367),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_640),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_207),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_60),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_26),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_11),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_297),
.Y(n_1351)
);

CKINVDCx14_ASAP7_75t_R g1352 ( 
.A(n_1028),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_826),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_826),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_826),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_826),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_853),
.Y(n_1357)
);

INVxp33_ASAP7_75t_SL g1358 ( 
.A(n_1136),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_826),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_826),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_826),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1329),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1329),
.Y(n_1363)
);

CKINVDCx16_ASAP7_75t_R g1364 ( 
.A(n_865),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1329),
.Y(n_1365)
);

CKINVDCx20_ASAP7_75t_R g1366 ( 
.A(n_1241),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1329),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_845),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1329),
.Y(n_1369)
);

CKINVDCx20_ASAP7_75t_R g1370 ( 
.A(n_1241),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1329),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1329),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1351),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1351),
.Y(n_1374)
);

INVxp67_ASAP7_75t_SL g1375 ( 
.A(n_1351),
.Y(n_1375)
);

CKINVDCx16_ASAP7_75t_R g1376 ( 
.A(n_1317),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_866),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_866),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_878),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_878),
.Y(n_1380)
);

BUFx3_ASAP7_75t_L g1381 ( 
.A(n_1270),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_899),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_899),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_948),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_948),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_973),
.Y(n_1386)
);

BUFx2_ASAP7_75t_SL g1387 ( 
.A(n_1270),
.Y(n_1387)
);

INVxp67_ASAP7_75t_L g1388 ( 
.A(n_1234),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_973),
.Y(n_1389)
);

INVxp33_ASAP7_75t_L g1390 ( 
.A(n_1346),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1010),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1010),
.Y(n_1392)
);

BUFx6f_ASAP7_75t_L g1393 ( 
.A(n_903),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1060),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_845),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_871),
.Y(n_1396)
);

CKINVDCx20_ASAP7_75t_R g1397 ( 
.A(n_1071),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1060),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1116),
.Y(n_1399)
);

BUFx3_ASAP7_75t_L g1400 ( 
.A(n_1116),
.Y(n_1400)
);

CKINVDCx20_ASAP7_75t_R g1401 ( 
.A(n_1191),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_820),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1193),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1193),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1213),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1213),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1296),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1296),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_949),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1331),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1331),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1345),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1345),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_820),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_820),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_820),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_820),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_843),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1214),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_843),
.Y(n_1420)
);

NOR2xp67_ASAP7_75t_L g1421 ( 
.A(n_811),
.B(n_1),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_843),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_996),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_843),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_843),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_893),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_893),
.Y(n_1427)
);

INVxp67_ASAP7_75t_SL g1428 ( 
.A(n_893),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_893),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_893),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_902),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_902),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_902),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_1199),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_1278),
.Y(n_1435)
);

CKINVDCx16_ASAP7_75t_R g1436 ( 
.A(n_1336),
.Y(n_1436)
);

CKINVDCx14_ASAP7_75t_R g1437 ( 
.A(n_875),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_902),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_911),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_902),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_905),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_905),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_905),
.Y(n_1443)
);

CKINVDCx20_ASAP7_75t_R g1444 ( 
.A(n_915),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_996),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_905),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_905),
.Y(n_1447)
);

INVxp67_ASAP7_75t_SL g1448 ( 
.A(n_1221),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1221),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1221),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_920),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1221),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_935),
.Y(n_1453)
);

INVxp67_ASAP7_75t_SL g1454 ( 
.A(n_1221),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1238),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1238),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1238),
.Y(n_1457)
);

INVxp67_ASAP7_75t_L g1458 ( 
.A(n_1272),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1238),
.Y(n_1459)
);

INVxp67_ASAP7_75t_SL g1460 ( 
.A(n_1238),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_903),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_937),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1259),
.Y(n_1463)
);

INVx3_ASAP7_75t_L g1464 ( 
.A(n_1259),
.Y(n_1464)
);

CKINVDCx14_ASAP7_75t_R g1465 ( 
.A(n_875),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1259),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1259),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1259),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_822),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_823),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_832),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_833),
.Y(n_1472)
);

INVxp67_ASAP7_75t_SL g1473 ( 
.A(n_824),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_836),
.Y(n_1474)
);

INVxp33_ASAP7_75t_L g1475 ( 
.A(n_976),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_840),
.Y(n_1476)
);

INVxp67_ASAP7_75t_L g1477 ( 
.A(n_1055),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_842),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_844),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_849),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_863),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_913),
.Y(n_1482)
);

CKINVDCx16_ASAP7_75t_R g1483 ( 
.A(n_815),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_868),
.Y(n_1484)
);

INVxp33_ASAP7_75t_SL g1485 ( 
.A(n_850),
.Y(n_1485)
);

INVxp67_ASAP7_75t_SL g1486 ( 
.A(n_824),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_874),
.Y(n_1487)
);

CKINVDCx20_ASAP7_75t_R g1488 ( 
.A(n_947),
.Y(n_1488)
);

INVxp33_ASAP7_75t_SL g1489 ( 
.A(n_850),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_876),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_886),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1428),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1358),
.B(n_1023),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1400),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1402),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1422),
.Y(n_1496)
);

INVx4_ASAP7_75t_L g1497 ( 
.A(n_1439),
.Y(n_1497)
);

BUFx6f_ASAP7_75t_L g1498 ( 
.A(n_1393),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_L g1499 ( 
.A(n_1393),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1403),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1447),
.Y(n_1501)
);

INVx3_ASAP7_75t_L g1502 ( 
.A(n_1464),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1428),
.Y(n_1503)
);

AND2x6_ASAP7_75t_L g1504 ( 
.A(n_1393),
.B(n_903),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1463),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1368),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1448),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_1444),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1453),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_SL g1510 ( 
.A1(n_1366),
.A2(n_848),
.B1(n_889),
.B2(n_885),
.Y(n_1510)
);

BUFx6f_ASAP7_75t_L g1511 ( 
.A(n_1393),
.Y(n_1511)
);

BUFx6f_ASAP7_75t_L g1512 ( 
.A(n_1461),
.Y(n_1512)
);

INVxp67_ASAP7_75t_L g1513 ( 
.A(n_1368),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1395),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1448),
.Y(n_1515)
);

INVx5_ASAP7_75t_L g1516 ( 
.A(n_1461),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_1461),
.Y(n_1517)
);

AND2x6_ASAP7_75t_L g1518 ( 
.A(n_1461),
.B(n_903),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_1464),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1355),
.A2(n_864),
.B(n_846),
.Y(n_1520)
);

BUFx12f_ASAP7_75t_L g1521 ( 
.A(n_1357),
.Y(n_1521)
);

CKINVDCx20_ASAP7_75t_R g1522 ( 
.A(n_1370),
.Y(n_1522)
);

INVx3_ASAP7_75t_L g1523 ( 
.A(n_1381),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1454),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1414),
.Y(n_1525)
);

BUFx8_ASAP7_75t_SL g1526 ( 
.A(n_1396),
.Y(n_1526)
);

OA21x2_ASAP7_75t_L g1527 ( 
.A1(n_1353),
.A2(n_916),
.B(n_881),
.Y(n_1527)
);

BUFx8_ASAP7_75t_SL g1528 ( 
.A(n_1409),
.Y(n_1528)
);

BUFx12f_ASAP7_75t_L g1529 ( 
.A(n_1419),
.Y(n_1529)
);

BUFx12f_ASAP7_75t_L g1530 ( 
.A(n_1435),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1395),
.Y(n_1531)
);

OA21x2_ASAP7_75t_L g1532 ( 
.A1(n_1354),
.A2(n_1002),
.B(n_926),
.Y(n_1532)
);

OA21x2_ASAP7_75t_L g1533 ( 
.A1(n_1356),
.A2(n_1075),
.B(n_1056),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1415),
.Y(n_1534)
);

NOR2x1_ASAP7_75t_L g1535 ( 
.A(n_1488),
.B(n_1266),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1416),
.Y(n_1536)
);

BUFx12f_ASAP7_75t_L g1537 ( 
.A(n_1451),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1417),
.Y(n_1538)
);

OA21x2_ASAP7_75t_L g1539 ( 
.A1(n_1359),
.A2(n_1180),
.B(n_1119),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1454),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1460),
.Y(n_1541)
);

CKINVDCx20_ASAP7_75t_R g1542 ( 
.A(n_1397),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1460),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1418),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1420),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1424),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_1462),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1425),
.Y(n_1548)
);

INVxp67_ASAP7_75t_L g1549 ( 
.A(n_1423),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1375),
.B(n_1119),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1426),
.Y(n_1551)
);

OA21x2_ASAP7_75t_L g1552 ( 
.A1(n_1360),
.A2(n_1180),
.B(n_901),
.Y(n_1552)
);

OA21x2_ASAP7_75t_L g1553 ( 
.A1(n_1361),
.A2(n_901),
.B(n_872),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1427),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1429),
.Y(n_1555)
);

INVxp33_ASAP7_75t_SL g1556 ( 
.A(n_1387),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1430),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1375),
.B(n_1334),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1421),
.B(n_815),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1431),
.Y(n_1560)
);

INVx4_ASAP7_75t_L g1561 ( 
.A(n_1362),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_1352),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1432),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1433),
.B(n_957),
.Y(n_1564)
);

INVx3_ASAP7_75t_L g1565 ( 
.A(n_1438),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1423),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1440),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1441),
.B(n_964),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1388),
.B(n_997),
.Y(n_1569)
);

BUFx6f_ASAP7_75t_L g1570 ( 
.A(n_1442),
.Y(n_1570)
);

OA21x2_ASAP7_75t_L g1571 ( 
.A1(n_1363),
.A2(n_945),
.B(n_872),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1377),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1443),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1446),
.Y(n_1574)
);

BUFx6f_ASAP7_75t_L g1575 ( 
.A(n_1449),
.Y(n_1575)
);

BUFx2_ASAP7_75t_L g1576 ( 
.A(n_1401),
.Y(n_1576)
);

OAI21x1_ASAP7_75t_L g1577 ( 
.A1(n_1372),
.A2(n_962),
.B(n_945),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1450),
.Y(n_1578)
);

BUFx3_ASAP7_75t_L g1579 ( 
.A(n_1378),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1452),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1455),
.Y(n_1581)
);

INVx3_ASAP7_75t_L g1582 ( 
.A(n_1456),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1457),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1459),
.B(n_991),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1466),
.B(n_1029),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_1352),
.Y(n_1586)
);

AND2x6_ASAP7_75t_L g1587 ( 
.A(n_1365),
.B(n_903),
.Y(n_1587)
);

AOI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1477),
.A2(n_885),
.B1(n_889),
.B2(n_848),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1437),
.B(n_815),
.Y(n_1589)
);

BUFx6f_ASAP7_75t_L g1590 ( 
.A(n_1467),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1468),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1388),
.B(n_997),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1379),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1367),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1369),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1373),
.B(n_1077),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1380),
.Y(n_1597)
);

BUFx6f_ASAP7_75t_L g1598 ( 
.A(n_1371),
.Y(n_1598)
);

BUFx6f_ASAP7_75t_L g1599 ( 
.A(n_1469),
.Y(n_1599)
);

BUFx12f_ASAP7_75t_L g1600 ( 
.A(n_1364),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1470),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1437),
.B(n_907),
.Y(n_1602)
);

INVxp67_ASAP7_75t_L g1603 ( 
.A(n_1445),
.Y(n_1603)
);

INVx6_ASAP7_75t_L g1604 ( 
.A(n_1483),
.Y(n_1604)
);

INVx4_ASAP7_75t_L g1605 ( 
.A(n_1482),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1471),
.Y(n_1606)
);

BUFx2_ASAP7_75t_L g1607 ( 
.A(n_1434),
.Y(n_1607)
);

INVx4_ASAP7_75t_L g1608 ( 
.A(n_1376),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1465),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1472),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1374),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1473),
.B(n_1093),
.Y(n_1612)
);

BUFx6f_ASAP7_75t_L g1613 ( 
.A(n_1474),
.Y(n_1613)
);

BUFx6f_ASAP7_75t_L g1614 ( 
.A(n_1476),
.Y(n_1614)
);

BUFx3_ASAP7_75t_L g1615 ( 
.A(n_1382),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1458),
.B(n_1021),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1513),
.B(n_1465),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1598),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1598),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1598),
.Y(n_1620)
);

BUFx6f_ASAP7_75t_L g1621 ( 
.A(n_1498),
.Y(n_1621)
);

INVx3_ASAP7_75t_L g1622 ( 
.A(n_1498),
.Y(n_1622)
);

BUFx2_ASAP7_75t_L g1623 ( 
.A(n_1494),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1519),
.Y(n_1624)
);

BUFx6f_ASAP7_75t_L g1625 ( 
.A(n_1498),
.Y(n_1625)
);

INVxp67_ASAP7_75t_L g1626 ( 
.A(n_1493),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1519),
.Y(n_1627)
);

BUFx6f_ASAP7_75t_L g1628 ( 
.A(n_1499),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1513),
.B(n_1475),
.Y(n_1629)
);

INVxp67_ASAP7_75t_L g1630 ( 
.A(n_1493),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1519),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1549),
.B(n_1475),
.Y(n_1632)
);

OAI21x1_ASAP7_75t_L g1633 ( 
.A1(n_1577),
.A2(n_1384),
.B(n_1383),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1615),
.Y(n_1634)
);

BUFx6f_ASAP7_75t_L g1635 ( 
.A(n_1499),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1549),
.B(n_1436),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1594),
.B(n_1595),
.Y(n_1637)
);

AND3x1_ASAP7_75t_L g1638 ( 
.A(n_1588),
.B(n_1445),
.C(n_1068),
.Y(n_1638)
);

BUFx6f_ASAP7_75t_L g1639 ( 
.A(n_1499),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1615),
.Y(n_1640)
);

BUFx6f_ASAP7_75t_L g1641 ( 
.A(n_1511),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1603),
.B(n_1390),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_SL g1643 ( 
.A(n_1556),
.B(n_1485),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1553),
.Y(n_1644)
);

INVxp67_ASAP7_75t_L g1645 ( 
.A(n_1506),
.Y(n_1645)
);

INVx1_ASAP7_75t_SL g1646 ( 
.A(n_1506),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1570),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_SL g1648 ( 
.A(n_1556),
.B(n_1489),
.Y(n_1648)
);

BUFx6f_ASAP7_75t_L g1649 ( 
.A(n_1511),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1514),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1553),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1571),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1571),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_SL g1654 ( 
.A(n_1609),
.B(n_1477),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1494),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1603),
.B(n_1390),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1492),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1503),
.Y(n_1658)
);

INVx3_ASAP7_75t_L g1659 ( 
.A(n_1511),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1507),
.Y(n_1660)
);

BUFx3_ASAP7_75t_L g1661 ( 
.A(n_1523),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1570),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1515),
.B(n_1458),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1570),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1500),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1575),
.Y(n_1666)
);

INVx1_ASAP7_75t_SL g1667 ( 
.A(n_1514),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1524),
.Y(n_1668)
);

AND2x6_ASAP7_75t_L g1669 ( 
.A(n_1589),
.B(n_962),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1540),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1531),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1575),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1541),
.B(n_1385),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1575),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1590),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1531),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1590),
.Y(n_1677)
);

AOI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1558),
.A2(n_896),
.B1(n_917),
.B2(n_891),
.Y(n_1678)
);

BUFx6f_ASAP7_75t_L g1679 ( 
.A(n_1512),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1590),
.Y(n_1680)
);

INVx3_ASAP7_75t_L g1681 ( 
.A(n_1512),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1500),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1495),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_SL g1684 ( 
.A(n_1609),
.B(n_1602),
.Y(n_1684)
);

INVx3_ASAP7_75t_L g1685 ( 
.A(n_1512),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1496),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1501),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_1547),
.Y(n_1688)
);

BUFx6f_ASAP7_75t_L g1689 ( 
.A(n_1517),
.Y(n_1689)
);

INVx3_ASAP7_75t_L g1690 ( 
.A(n_1517),
.Y(n_1690)
);

INVx3_ASAP7_75t_L g1691 ( 
.A(n_1517),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1543),
.Y(n_1692)
);

BUFx6f_ASAP7_75t_L g1693 ( 
.A(n_1520),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1572),
.Y(n_1694)
);

AOI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1558),
.A2(n_896),
.B1(n_917),
.B2(n_891),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1505),
.Y(n_1696)
);

HB1xp67_ASAP7_75t_L g1697 ( 
.A(n_1566),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1566),
.B(n_1386),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1561),
.B(n_1473),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1561),
.B(n_1486),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1579),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1525),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1593),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1605),
.B(n_1486),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1534),
.Y(n_1705)
);

AND2x6_ASAP7_75t_L g1706 ( 
.A(n_1535),
.B(n_966),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1597),
.Y(n_1707)
);

INVx1_ASAP7_75t_SL g1708 ( 
.A(n_1542),
.Y(n_1708)
);

BUFx6f_ASAP7_75t_L g1709 ( 
.A(n_1599),
.Y(n_1709)
);

AND2x4_ASAP7_75t_L g1710 ( 
.A(n_1523),
.B(n_1389),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1536),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1502),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1538),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1502),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1605),
.B(n_913),
.Y(n_1715)
);

INVx1_ASAP7_75t_SL g1716 ( 
.A(n_1542),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1552),
.B(n_913),
.Y(n_1717)
);

INVxp67_ASAP7_75t_L g1718 ( 
.A(n_1612),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1509),
.B(n_1391),
.Y(n_1719)
);

BUFx6f_ASAP7_75t_L g1720 ( 
.A(n_1599),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1611),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1599),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1613),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1562),
.B(n_1102),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1613),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1612),
.B(n_1392),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1613),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1614),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1614),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1544),
.Y(n_1730)
);

BUFx3_ASAP7_75t_L g1731 ( 
.A(n_1537),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1545),
.Y(n_1732)
);

INVxp67_ASAP7_75t_L g1733 ( 
.A(n_1596),
.Y(n_1733)
);

INVx1_ASAP7_75t_SL g1734 ( 
.A(n_1522),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1614),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1546),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1548),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1554),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1551),
.Y(n_1739)
);

BUFx6f_ASAP7_75t_L g1740 ( 
.A(n_1552),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1555),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1569),
.B(n_1394),
.Y(n_1742)
);

INVx3_ASAP7_75t_L g1743 ( 
.A(n_1516),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1560),
.Y(n_1744)
);

INVx1_ASAP7_75t_SL g1745 ( 
.A(n_1522),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1557),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1563),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1569),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1567),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1578),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1721),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1683),
.Y(n_1752)
);

AND2x6_ASAP7_75t_L g1753 ( 
.A(n_1644),
.B(n_1651),
.Y(n_1753)
);

INVx3_ASAP7_75t_L g1754 ( 
.A(n_1661),
.Y(n_1754)
);

BUFx2_ASAP7_75t_L g1755 ( 
.A(n_1650),
.Y(n_1755)
);

INVx4_ASAP7_75t_L g1756 ( 
.A(n_1709),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1657),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1718),
.B(n_1550),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1658),
.Y(n_1759)
);

INVx2_ASAP7_75t_SL g1760 ( 
.A(n_1623),
.Y(n_1760)
);

AO21x2_ASAP7_75t_L g1761 ( 
.A1(n_1652),
.A2(n_1550),
.B(n_1564),
.Y(n_1761)
);

INVx4_ASAP7_75t_L g1762 ( 
.A(n_1709),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_SL g1763 ( 
.A(n_1718),
.B(n_1733),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1686),
.Y(n_1764)
);

INVx3_ASAP7_75t_L g1765 ( 
.A(n_1633),
.Y(n_1765)
);

OAI21xp33_ASAP7_75t_SL g1766 ( 
.A1(n_1653),
.A2(n_1559),
.B(n_1596),
.Y(n_1766)
);

OR2x6_ASAP7_75t_L g1767 ( 
.A(n_1731),
.B(n_1600),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1687),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1646),
.B(n_1592),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_L g1770 ( 
.A(n_1646),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1660),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1668),
.Y(n_1772)
);

INVx2_ASAP7_75t_SL g1773 ( 
.A(n_1719),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1667),
.B(n_1592),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1670),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1692),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1696),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1712),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1714),
.Y(n_1779)
);

INVx3_ASAP7_75t_L g1780 ( 
.A(n_1719),
.Y(n_1780)
);

BUFx10_ASAP7_75t_L g1781 ( 
.A(n_1688),
.Y(n_1781)
);

AOI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1733),
.A2(n_1547),
.B1(n_1497),
.B2(n_1564),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1702),
.Y(n_1783)
);

INVx2_ASAP7_75t_SL g1784 ( 
.A(n_1655),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1710),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1726),
.B(n_1568),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1699),
.B(n_1568),
.Y(n_1787)
);

AND2x6_ASAP7_75t_L g1788 ( 
.A(n_1740),
.B(n_1616),
.Y(n_1788)
);

INVx3_ASAP7_75t_L g1789 ( 
.A(n_1710),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1699),
.B(n_1584),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1634),
.B(n_1640),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1626),
.A2(n_1497),
.B1(n_1584),
.B2(n_1585),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1700),
.B(n_1585),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1705),
.Y(n_1794)
);

BUFx3_ASAP7_75t_L g1795 ( 
.A(n_1694),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1667),
.B(n_1608),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1736),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1711),
.Y(n_1798)
);

NAND2xp33_ASAP7_75t_L g1799 ( 
.A(n_1669),
.B(n_1504),
.Y(n_1799)
);

INVx5_ASAP7_75t_L g1800 ( 
.A(n_1669),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_SL g1801 ( 
.A(n_1626),
.B(n_1562),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1738),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1746),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1630),
.B(n_1586),
.Y(n_1804)
);

AND2x6_ASAP7_75t_L g1805 ( 
.A(n_1740),
.B(n_1616),
.Y(n_1805)
);

OR2x6_ASAP7_75t_L g1806 ( 
.A(n_1650),
.B(n_1604),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1642),
.B(n_1656),
.Y(n_1807)
);

NOR2xp33_ASAP7_75t_L g1808 ( 
.A(n_1630),
.B(n_1608),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1645),
.B(n_1604),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_1734),
.Y(n_1810)
);

INVx4_ASAP7_75t_L g1811 ( 
.A(n_1709),
.Y(n_1811)
);

NAND2x1p5_ASAP7_75t_L g1812 ( 
.A(n_1720),
.B(n_1601),
.Y(n_1812)
);

INVx4_ASAP7_75t_L g1813 ( 
.A(n_1720),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_1734),
.Y(n_1814)
);

INVx1_ASAP7_75t_SL g1815 ( 
.A(n_1629),
.Y(n_1815)
);

BUFx3_ASAP7_75t_L g1816 ( 
.A(n_1701),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_SL g1817 ( 
.A(n_1636),
.B(n_1521),
.Y(n_1817)
);

NAND2x1p5_ASAP7_75t_L g1818 ( 
.A(n_1720),
.B(n_1606),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1713),
.Y(n_1819)
);

HB1xp67_ASAP7_75t_L g1820 ( 
.A(n_1671),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1632),
.B(n_1559),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1617),
.B(n_1586),
.Y(n_1822)
);

AND3x2_ASAP7_75t_L g1823 ( 
.A(n_1748),
.B(n_1607),
.C(n_1576),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1747),
.Y(n_1824)
);

XNOR2x2_ASAP7_75t_SL g1825 ( 
.A(n_1678),
.B(n_1588),
.Y(n_1825)
);

NOR2xp33_ASAP7_75t_SL g1826 ( 
.A(n_1671),
.B(n_1529),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1749),
.Y(n_1827)
);

AND2x6_ASAP7_75t_L g1828 ( 
.A(n_1740),
.B(n_966),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_SL g1829 ( 
.A(n_1748),
.B(n_1508),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1750),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1700),
.B(n_1539),
.Y(n_1831)
);

BUFx2_ASAP7_75t_L g1832 ( 
.A(n_1676),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1730),
.Y(n_1833)
);

BUFx4f_ASAP7_75t_L g1834 ( 
.A(n_1706),
.Y(n_1834)
);

BUFx2_ASAP7_75t_L g1835 ( 
.A(n_1676),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1732),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1737),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1697),
.B(n_1508),
.Y(n_1838)
);

INVx1_ASAP7_75t_SL g1839 ( 
.A(n_1745),
.Y(n_1839)
);

INVx4_ASAP7_75t_SL g1840 ( 
.A(n_1706),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1704),
.B(n_1539),
.Y(n_1841)
);

AND2x4_ASAP7_75t_L g1842 ( 
.A(n_1703),
.B(n_1610),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1739),
.Y(n_1843)
);

INVx4_ASAP7_75t_L g1844 ( 
.A(n_1621),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1704),
.B(n_1527),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1637),
.B(n_1618),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1741),
.Y(n_1847)
);

INVx2_ASAP7_75t_SL g1848 ( 
.A(n_1665),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1697),
.B(n_1510),
.Y(n_1849)
);

OR2x6_ASAP7_75t_L g1850 ( 
.A(n_1645),
.B(n_1604),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_SL g1851 ( 
.A(n_1663),
.B(n_1120),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1744),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1637),
.Y(n_1853)
);

AOI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1669),
.A2(n_1198),
.B1(n_1299),
.B2(n_1166),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1619),
.B(n_1527),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1622),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_SL g1857 ( 
.A(n_1707),
.B(n_1583),
.Y(n_1857)
);

INVx3_ASAP7_75t_L g1858 ( 
.A(n_1622),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_SL g1859 ( 
.A(n_1643),
.B(n_1580),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1659),
.Y(n_1860)
);

INVx3_ASAP7_75t_L g1861 ( 
.A(n_1659),
.Y(n_1861)
);

HB1xp67_ASAP7_75t_L g1862 ( 
.A(n_1682),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1620),
.B(n_1532),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1715),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_L g1865 ( 
.A(n_1648),
.B(n_1530),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_SL g1866 ( 
.A(n_1745),
.B(n_1526),
.Y(n_1866)
);

AND2x4_ASAP7_75t_L g1867 ( 
.A(n_1722),
.B(n_1478),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1715),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1681),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1669),
.B(n_1532),
.Y(n_1870)
);

INVx4_ASAP7_75t_L g1871 ( 
.A(n_1621),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1624),
.Y(n_1872)
);

BUFx3_ASAP7_75t_L g1873 ( 
.A(n_1723),
.Y(n_1873)
);

AOI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1706),
.A2(n_1533),
.B1(n_1581),
.B2(n_1587),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_L g1875 ( 
.A(n_1654),
.B(n_883),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1673),
.B(n_1533),
.Y(n_1876)
);

INVx3_ASAP7_75t_L g1877 ( 
.A(n_1681),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1706),
.B(n_1573),
.Y(n_1878)
);

NAND3x1_ASAP7_75t_L g1879 ( 
.A(n_1678),
.B(n_959),
.C(n_938),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1627),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1631),
.Y(n_1881)
);

INVx3_ASAP7_75t_L g1882 ( 
.A(n_1647),
.Y(n_1882)
);

NAND2xp33_ASAP7_75t_L g1883 ( 
.A(n_1693),
.B(n_1504),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1685),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1662),
.B(n_1574),
.Y(n_1885)
);

BUFx4f_ASAP7_75t_L g1886 ( 
.A(n_1698),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1742),
.B(n_1398),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1695),
.B(n_1399),
.Y(n_1888)
);

INVx3_ASAP7_75t_L g1889 ( 
.A(n_1664),
.Y(n_1889)
);

INVx3_ASAP7_75t_R g1890 ( 
.A(n_1708),
.Y(n_1890)
);

INVx6_ASAP7_75t_L g1891 ( 
.A(n_1621),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1685),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1725),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1727),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_SL g1895 ( 
.A(n_1728),
.B(n_913),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1666),
.B(n_1591),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1729),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1672),
.B(n_1565),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1735),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1674),
.B(n_1565),
.Y(n_1900)
);

CKINVDCx5p33_ASAP7_75t_R g1901 ( 
.A(n_1708),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1690),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_SL g1903 ( 
.A(n_1684),
.B(n_913),
.Y(n_1903)
);

AND2x4_ASAP7_75t_L g1904 ( 
.A(n_1675),
.B(n_1479),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1677),
.B(n_1582),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1690),
.Y(n_1906)
);

INVx4_ASAP7_75t_L g1907 ( 
.A(n_1625),
.Y(n_1907)
);

AND2x6_ASAP7_75t_L g1908 ( 
.A(n_1717),
.B(n_1043),
.Y(n_1908)
);

BUFx6f_ASAP7_75t_L g1909 ( 
.A(n_1625),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1904),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1904),
.Y(n_1911)
);

NOR3xp33_ASAP7_75t_L g1912 ( 
.A(n_1801),
.B(n_1510),
.C(n_1716),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1752),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1764),
.Y(n_1914)
);

BUFx6f_ASAP7_75t_SL g1915 ( 
.A(n_1781),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1769),
.B(n_1695),
.Y(n_1916)
);

INVxp67_ASAP7_75t_L g1917 ( 
.A(n_1770),
.Y(n_1917)
);

AO221x1_ASAP7_75t_L g1918 ( 
.A1(n_1825),
.A2(n_1049),
.B1(n_953),
.B2(n_831),
.C(n_1638),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_L g1919 ( 
.A(n_1763),
.B(n_1716),
.Y(n_1919)
);

INVxp67_ASAP7_75t_L g1920 ( 
.A(n_1774),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1787),
.B(n_1717),
.Y(n_1921)
);

AOI22xp33_ASAP7_75t_SL g1922 ( 
.A1(n_1875),
.A2(n_918),
.B1(n_965),
.B2(n_943),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1758),
.B(n_1815),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1757),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1790),
.B(n_1680),
.Y(n_1925)
);

INVx2_ASAP7_75t_SL g1926 ( 
.A(n_1755),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1759),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1793),
.B(n_1691),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1886),
.B(n_1638),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_SL g1930 ( 
.A(n_1782),
.B(n_1792),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1786),
.B(n_1691),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1771),
.Y(n_1932)
);

NOR2xp67_ASAP7_75t_L g1933 ( 
.A(n_1865),
.B(n_1796),
.Y(n_1933)
);

AOI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1908),
.A2(n_1693),
.B1(n_913),
.B2(n_1587),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1768),
.Y(n_1935)
);

INVxp67_ASAP7_75t_L g1936 ( 
.A(n_1820),
.Y(n_1936)
);

NOR2xp33_ASAP7_75t_L g1937 ( 
.A(n_1808),
.B(n_1724),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1839),
.B(n_1526),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1853),
.B(n_1864),
.Y(n_1939)
);

INVx2_ASAP7_75t_SL g1940 ( 
.A(n_1755),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1777),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1868),
.B(n_1625),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_L g1943 ( 
.A(n_1838),
.B(n_1528),
.Y(n_1943)
);

INVxp67_ASAP7_75t_L g1944 ( 
.A(n_1832),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1788),
.B(n_1628),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_SL g1946 ( 
.A(n_1821),
.B(n_1628),
.Y(n_1946)
);

BUFx2_ASAP7_75t_L g1947 ( 
.A(n_1810),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1788),
.B(n_1628),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1772),
.Y(n_1949)
);

INVx2_ASAP7_75t_SL g1950 ( 
.A(n_1832),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1783),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1807),
.B(n_1404),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_SL g1953 ( 
.A(n_1834),
.B(n_1635),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1775),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1776),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1794),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1867),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1788),
.B(n_1805),
.Y(n_1958)
);

BUFx5_ASAP7_75t_L g1959 ( 
.A(n_1753),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1798),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1805),
.B(n_1635),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1805),
.B(n_1635),
.Y(n_1962)
);

AOI22xp33_ASAP7_75t_L g1963 ( 
.A1(n_1908),
.A2(n_1693),
.B1(n_913),
.B2(n_1587),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1887),
.B(n_1405),
.Y(n_1964)
);

NAND2x1_ASAP7_75t_L g1965 ( 
.A(n_1756),
.B(n_1639),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1835),
.B(n_1406),
.Y(n_1966)
);

BUFx3_ASAP7_75t_L g1967 ( 
.A(n_1835),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1846),
.B(n_1639),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1761),
.B(n_1639),
.Y(n_1969)
);

NAND2x1p5_ASAP7_75t_L g1970 ( 
.A(n_1800),
.B(n_1641),
.Y(n_1970)
);

NOR2xp67_ASAP7_75t_L g1971 ( 
.A(n_1760),
.B(n_1407),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1819),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1833),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1753),
.B(n_1582),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_SL g1975 ( 
.A(n_1800),
.B(n_1641),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_1862),
.B(n_1528),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1908),
.B(n_1641),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_SL g1978 ( 
.A(n_1800),
.B(n_1649),
.Y(n_1978)
);

NOR2xp33_ASAP7_75t_L g1979 ( 
.A(n_1784),
.B(n_918),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_SL g1980 ( 
.A(n_1789),
.B(n_1649),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1751),
.B(n_1649),
.Y(n_1981)
);

INVx3_ASAP7_75t_L g1982 ( 
.A(n_1858),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1797),
.B(n_1679),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_SL g1984 ( 
.A(n_1848),
.B(n_1679),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1837),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1867),
.Y(n_1986)
);

AND2x4_ASAP7_75t_L g1987 ( 
.A(n_1754),
.B(n_1480),
.Y(n_1987)
);

AOI22xp33_ASAP7_75t_L g1988 ( 
.A1(n_1828),
.A2(n_1587),
.B1(n_965),
.B2(n_1011),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1802),
.B(n_1679),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1753),
.B(n_1689),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1803),
.Y(n_1991)
);

INVx2_ASAP7_75t_SL g1992 ( 
.A(n_1806),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1824),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1827),
.B(n_1689),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_SL g1995 ( 
.A(n_1780),
.B(n_1689),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1830),
.B(n_1587),
.Y(n_1996)
);

AND2x6_ASAP7_75t_SL g1997 ( 
.A(n_1806),
.B(n_909),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1831),
.B(n_1021),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_SL g1999 ( 
.A(n_1791),
.B(n_1516),
.Y(n_1999)
);

AOI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1766),
.A2(n_1791),
.B1(n_1903),
.B2(n_1828),
.Y(n_2000)
);

AOI22xp33_ASAP7_75t_L g2001 ( 
.A1(n_1828),
.A2(n_1011),
.B1(n_1051),
.B2(n_943),
.Y(n_2001)
);

INVx4_ASAP7_75t_SL g2002 ( 
.A(n_1891),
.Y(n_2002)
);

INVx2_ASAP7_75t_SL g2003 ( 
.A(n_1814),
.Y(n_2003)
);

INVx2_ASAP7_75t_SL g2004 ( 
.A(n_1901),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1845),
.B(n_1068),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1841),
.B(n_1086),
.Y(n_2006)
);

BUFx3_ASAP7_75t_L g2007 ( 
.A(n_1781),
.Y(n_2007)
);

AO221x1_ASAP7_75t_L g2008 ( 
.A1(n_1858),
.A2(n_923),
.B1(n_934),
.B2(n_933),
.C(n_910),
.Y(n_2008)
);

INVx3_ASAP7_75t_L g2009 ( 
.A(n_1861),
.Y(n_2009)
);

INVx1_ASAP7_75t_SL g2010 ( 
.A(n_1849),
.Y(n_2010)
);

AOI22xp33_ASAP7_75t_L g2011 ( 
.A1(n_1888),
.A2(n_1051),
.B1(n_1097),
.B2(n_1079),
.Y(n_2011)
);

O2A1O1Ixp5_ASAP7_75t_L g2012 ( 
.A1(n_1876),
.A2(n_1087),
.B(n_1118),
.C(n_1043),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_SL g2013 ( 
.A(n_1773),
.B(n_1516),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1855),
.B(n_1086),
.Y(n_2014)
);

BUFx6f_ASAP7_75t_L g2015 ( 
.A(n_1909),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1809),
.B(n_1408),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1836),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1778),
.B(n_1110),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1779),
.B(n_1110),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1850),
.B(n_1410),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1843),
.B(n_1178),
.Y(n_2021)
);

NOR2xp33_ASAP7_75t_L g2022 ( 
.A(n_1804),
.B(n_1079),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1847),
.B(n_1178),
.Y(n_2023)
);

NOR2xp33_ASAP7_75t_L g2024 ( 
.A(n_1851),
.B(n_1097),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_SL g2025 ( 
.A(n_1842),
.B(n_1516),
.Y(n_2025)
);

AOI22xp33_ASAP7_75t_L g2026 ( 
.A1(n_1863),
.A2(n_1104),
.B1(n_1109),
.B2(n_1105),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1852),
.B(n_1310),
.Y(n_2027)
);

OR2x2_ASAP7_75t_L g2028 ( 
.A(n_1829),
.B(n_1411),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_SL g2029 ( 
.A(n_1842),
.B(n_1104),
.Y(n_2029)
);

INVxp67_ASAP7_75t_L g2030 ( 
.A(n_1859),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1861),
.B(n_1310),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_SL g2032 ( 
.A(n_1756),
.B(n_1105),
.Y(n_2032)
);

HB1xp67_ASAP7_75t_L g2033 ( 
.A(n_1890),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_SL g2034 ( 
.A(n_1762),
.B(n_1109),
.Y(n_2034)
);

NOR2xp33_ASAP7_75t_L g2035 ( 
.A(n_1822),
.B(n_1115),
.Y(n_2035)
);

NOR2xp33_ASAP7_75t_L g2036 ( 
.A(n_1795),
.B(n_1115),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1877),
.B(n_812),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1877),
.B(n_813),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1785),
.B(n_814),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1856),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_1870),
.B(n_887),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1893),
.B(n_816),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1860),
.Y(n_2043)
);

BUFx6f_ASAP7_75t_SL g2044 ( 
.A(n_1767),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1869),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1894),
.B(n_817),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1885),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1897),
.B(n_818),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1884),
.Y(n_2049)
);

OAI22xp33_ASAP7_75t_L g2050 ( 
.A1(n_1817),
.A2(n_1133),
.B1(n_1141),
.B2(n_1128),
.Y(n_2050)
);

BUFx3_ASAP7_75t_L g2051 ( 
.A(n_1816),
.Y(n_2051)
);

NOR2x1p5_ASAP7_75t_L g2052 ( 
.A(n_1873),
.B(n_1412),
.Y(n_2052)
);

INVx3_ASAP7_75t_L g2053 ( 
.A(n_1909),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_SL g2054 ( 
.A(n_1762),
.B(n_1128),
.Y(n_2054)
);

INVxp67_ASAP7_75t_SL g2055 ( 
.A(n_1909),
.Y(n_2055)
);

AOI22xp33_ASAP7_75t_L g2056 ( 
.A1(n_1878),
.A2(n_1141),
.B1(n_1147),
.B2(n_1133),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1899),
.B(n_819),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_SL g2058 ( 
.A(n_1811),
.B(n_1147),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_SL g2059 ( 
.A(n_1811),
.B(n_1170),
.Y(n_2059)
);

BUFx6f_ASAP7_75t_SL g2060 ( 
.A(n_1767),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_SL g2061 ( 
.A(n_1813),
.B(n_1170),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_1850),
.B(n_1413),
.Y(n_2062)
);

NOR2xp33_ASAP7_75t_L g2063 ( 
.A(n_1872),
.B(n_1187),
.Y(n_2063)
);

OAI221xp5_ASAP7_75t_L g2064 ( 
.A1(n_1857),
.A2(n_1007),
.B1(n_1015),
.B2(n_992),
.C(n_895),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_SL g2065 ( 
.A(n_1813),
.B(n_1187),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1880),
.B(n_821),
.Y(n_2066)
);

INVx2_ASAP7_75t_SL g2067 ( 
.A(n_1881),
.Y(n_2067)
);

AOI22xp33_ASAP7_75t_L g2068 ( 
.A1(n_1895),
.A2(n_1237),
.B1(n_1258),
.B2(n_1204),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1892),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1874),
.B(n_1059),
.Y(n_2070)
);

NAND2xp33_ASAP7_75t_SL g2071 ( 
.A(n_1844),
.B(n_1204),
.Y(n_2071)
);

NOR2xp33_ASAP7_75t_L g2072 ( 
.A(n_1826),
.B(n_1237),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_1840),
.B(n_1066),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_SL g2074 ( 
.A(n_1840),
.B(n_1258),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1902),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1906),
.B(n_825),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1896),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_1866),
.B(n_907),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1898),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1882),
.B(n_827),
.Y(n_2080)
);

AOI22xp5_ASAP7_75t_L g2081 ( 
.A1(n_1937),
.A2(n_1854),
.B1(n_1879),
.B2(n_1889),
.Y(n_2081)
);

INVx1_ASAP7_75t_SL g2082 ( 
.A(n_1967),
.Y(n_2082)
);

NAND2x1p5_ASAP7_75t_L g2083 ( 
.A(n_2051),
.B(n_1844),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_1923),
.B(n_1823),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1921),
.B(n_1900),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1924),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_1916),
.B(n_1812),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1927),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_SL g2089 ( 
.A(n_1933),
.B(n_1871),
.Y(n_2089)
);

CKINVDCx5p33_ASAP7_75t_R g2090 ( 
.A(n_1915),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_1921),
.B(n_1905),
.Y(n_2091)
);

AOI22xp33_ASAP7_75t_L g2092 ( 
.A1(n_1930),
.A2(n_1799),
.B1(n_1818),
.B2(n_1871),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_1993),
.Y(n_2093)
);

INVx5_ASAP7_75t_L g2094 ( 
.A(n_2015),
.Y(n_2094)
);

NOR2xp33_ASAP7_75t_L g2095 ( 
.A(n_2010),
.B(n_1907),
.Y(n_2095)
);

O2A1O1Ixp33_ASAP7_75t_SL g2096 ( 
.A1(n_1939),
.A2(n_1765),
.B(n_1235),
.C(n_1236),
.Y(n_2096)
);

AOI22xp33_ASAP7_75t_L g2097 ( 
.A1(n_2024),
.A2(n_1907),
.B1(n_1891),
.B2(n_1883),
.Y(n_2097)
);

NOR2xp33_ASAP7_75t_L g2098 ( 
.A(n_2010),
.B(n_1269),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1932),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1949),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1925),
.B(n_1155),
.Y(n_2101)
);

NAND2x1_ASAP7_75t_L g2102 ( 
.A(n_1982),
.B(n_1765),
.Y(n_2102)
);

BUFx5_ASAP7_75t_L g2103 ( 
.A(n_2079),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2041),
.B(n_1242),
.Y(n_2104)
);

INVxp67_ASAP7_75t_L g2105 ( 
.A(n_1926),
.Y(n_2105)
);

CKINVDCx8_ASAP7_75t_R g2106 ( 
.A(n_1997),
.Y(n_2106)
);

A2O1A1Ixp33_ASAP7_75t_L g2107 ( 
.A1(n_2022),
.A2(n_942),
.B(n_951),
.C(n_939),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1954),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1955),
.Y(n_2109)
);

INVx3_ASAP7_75t_L g2110 ( 
.A(n_2007),
.Y(n_2110)
);

BUFx4f_ASAP7_75t_L g2111 ( 
.A(n_1940),
.Y(n_2111)
);

NAND2xp33_ASAP7_75t_SL g2112 ( 
.A(n_1915),
.B(n_2073),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1913),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1991),
.Y(n_2114)
);

AOI21xp5_ASAP7_75t_L g2115 ( 
.A1(n_1928),
.A2(n_1743),
.B(n_1518),
.Y(n_2115)
);

NOR2xp67_ASAP7_75t_L g2116 ( 
.A(n_2003),
.B(n_765),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2017),
.Y(n_2117)
);

CKINVDCx5p33_ASAP7_75t_R g2118 ( 
.A(n_1947),
.Y(n_2118)
);

NOR2xp33_ASAP7_75t_L g2119 ( 
.A(n_1944),
.B(n_1269),
.Y(n_2119)
);

OAI22xp5_ASAP7_75t_L g2120 ( 
.A1(n_2000),
.A2(n_1304),
.B1(n_1293),
.B2(n_1282),
.Y(n_2120)
);

OAI22xp5_ASAP7_75t_SL g2121 ( 
.A1(n_1922),
.A2(n_1304),
.B1(n_1293),
.B2(n_862),
.Y(n_2121)
);

BUFx6f_ASAP7_75t_L g2122 ( 
.A(n_2015),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_SL g2123 ( 
.A(n_1920),
.B(n_1481),
.Y(n_2123)
);

BUFx2_ASAP7_75t_L g2124 ( 
.A(n_2033),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1914),
.Y(n_2125)
);

BUFx6f_ASAP7_75t_L g2126 ( 
.A(n_2015),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_1935),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_2041),
.B(n_1246),
.Y(n_2128)
);

CKINVDCx5p33_ASAP7_75t_R g2129 ( 
.A(n_2044),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1941),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1951),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_1952),
.B(n_2016),
.Y(n_2132)
);

AND2x6_ASAP7_75t_SL g2133 ( 
.A(n_1938),
.B(n_956),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1956),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1931),
.B(n_1312),
.Y(n_2135)
);

BUFx3_ASAP7_75t_L g2136 ( 
.A(n_1950),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_1960),
.Y(n_2137)
);

INVx3_ASAP7_75t_L g2138 ( 
.A(n_1987),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1972),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1973),
.Y(n_2140)
);

OAI22xp5_ASAP7_75t_L g2141 ( 
.A1(n_2070),
.A2(n_1349),
.B1(n_829),
.B2(n_830),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_1985),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2021),
.Y(n_2143)
);

INVx5_ASAP7_75t_L g2144 ( 
.A(n_1997),
.Y(n_2144)
);

INVx3_ASAP7_75t_L g2145 ( 
.A(n_1987),
.Y(n_2145)
);

BUFx8_ASAP7_75t_L g2146 ( 
.A(n_2044),
.Y(n_2146)
);

BUFx3_ASAP7_75t_L g2147 ( 
.A(n_1992),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2047),
.B(n_828),
.Y(n_2148)
);

AND2x4_ASAP7_75t_L g2149 ( 
.A(n_1957),
.B(n_1484),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2023),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_1982),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2027),
.Y(n_2152)
);

AND2x4_ASAP7_75t_L g2153 ( 
.A(n_1986),
.B(n_1487),
.Y(n_2153)
);

NAND2x1p5_ASAP7_75t_L g2154 ( 
.A(n_2053),
.B(n_1490),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_SL g2155 ( 
.A(n_2004),
.B(n_1491),
.Y(n_2155)
);

AND2x6_ASAP7_75t_L g2156 ( 
.A(n_1958),
.B(n_1087),
.Y(n_2156)
);

INVxp67_ASAP7_75t_L g2157 ( 
.A(n_1919),
.Y(n_2157)
);

INVx2_ASAP7_75t_SL g2158 ( 
.A(n_2020),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1981),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_2077),
.B(n_1964),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1968),
.B(n_834),
.Y(n_2161)
);

NOR3xp33_ASAP7_75t_SL g2162 ( 
.A(n_2050),
.B(n_852),
.C(n_851),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1983),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1989),
.Y(n_2164)
);

OAI21x1_ASAP7_75t_L g2165 ( 
.A1(n_2012),
.A2(n_1743),
.B(n_1181),
.Y(n_2165)
);

AOI22xp33_ASAP7_75t_L g2166 ( 
.A1(n_1918),
.A2(n_1181),
.B1(n_1183),
.B2(n_1118),
.Y(n_2166)
);

CKINVDCx5p33_ASAP7_75t_R g2167 ( 
.A(n_2060),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2070),
.B(n_835),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_2030),
.B(n_837),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_1966),
.B(n_838),
.Y(n_2170)
);

AOI22xp5_ASAP7_75t_L g2171 ( 
.A1(n_1912),
.A2(n_841),
.B1(n_847),
.B2(n_839),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2009),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_1942),
.B(n_884),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_2009),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_2006),
.B(n_888),
.Y(n_2175)
);

INVxp33_ASAP7_75t_SL g2176 ( 
.A(n_1943),
.Y(n_2176)
);

OR2x4_ASAP7_75t_L g2177 ( 
.A(n_2072),
.B(n_960),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2006),
.B(n_890),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_SL g2179 ( 
.A(n_1988),
.B(n_892),
.Y(n_2179)
);

NAND2x1p5_ASAP7_75t_L g2180 ( 
.A(n_2053),
.B(n_961),
.Y(n_2180)
);

NOR2xp33_ASAP7_75t_L g2181 ( 
.A(n_1917),
.B(n_894),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1994),
.Y(n_2182)
);

INVx2_ASAP7_75t_SL g2183 ( 
.A(n_2062),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2005),
.B(n_897),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2031),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_2040),
.Y(n_2186)
);

BUFx6f_ASAP7_75t_L g2187 ( 
.A(n_1984),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1910),
.Y(n_2188)
);

HB1xp67_ASAP7_75t_L g2189 ( 
.A(n_1936),
.Y(n_2189)
);

O2A1O1Ixp33_ASAP7_75t_L g2190 ( 
.A1(n_2064),
.A2(n_971),
.B(n_982),
.C(n_967),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1911),
.Y(n_2191)
);

AOI22xp5_ASAP7_75t_L g2192 ( 
.A1(n_2035),
.A2(n_900),
.B1(n_904),
.B2(n_898),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_SL g2193 ( 
.A(n_2036),
.B(n_906),
.Y(n_2193)
);

CKINVDCx5p33_ASAP7_75t_R g2194 ( 
.A(n_2060),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2018),
.Y(n_2195)
);

NOR2x1_ASAP7_75t_R g2196 ( 
.A(n_2074),
.B(n_851),
.Y(n_2196)
);

AOI22xp5_ASAP7_75t_L g2197 ( 
.A1(n_2032),
.A2(n_912),
.B1(n_914),
.B2(n_908),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_2005),
.B(n_919),
.Y(n_2198)
);

AND2x4_ASAP7_75t_L g2199 ( 
.A(n_2052),
.B(n_985),
.Y(n_2199)
);

AO21x1_ASAP7_75t_L g2200 ( 
.A1(n_1969),
.A2(n_1000),
.B(n_994),
.Y(n_2200)
);

BUFx3_ASAP7_75t_L g2201 ( 
.A(n_1976),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2019),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2043),
.Y(n_2203)
);

O2A1O1Ixp33_ASAP7_75t_L g2204 ( 
.A1(n_1929),
.A2(n_1009),
.B(n_1012),
.C(n_1004),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_1946),
.B(n_2014),
.Y(n_2205)
);

AOI22xp33_ASAP7_75t_L g2206 ( 
.A1(n_2008),
.A2(n_1184),
.B1(n_1217),
.B2(n_1183),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_1979),
.B(n_2063),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2045),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_SL g2209 ( 
.A(n_2067),
.B(n_921),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_SL g2210 ( 
.A(n_2073),
.B(n_922),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2049),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2069),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_2075),
.Y(n_2213)
);

CKINVDCx11_ASAP7_75t_R g2214 ( 
.A(n_2002),
.Y(n_2214)
);

INVxp67_ASAP7_75t_L g2215 ( 
.A(n_2028),
.Y(n_2215)
);

AOI22xp33_ASAP7_75t_L g2216 ( 
.A1(n_2071),
.A2(n_1217),
.B1(n_1228),
.B2(n_1184),
.Y(n_2216)
);

AOI22xp5_ASAP7_75t_L g2217 ( 
.A1(n_2034),
.A2(n_925),
.B1(n_927),
.B2(n_924),
.Y(n_2217)
);

AND2x4_ASAP7_75t_L g2218 ( 
.A(n_2002),
.B(n_1013),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2014),
.Y(n_2219)
);

BUFx3_ASAP7_75t_L g2220 ( 
.A(n_2078),
.Y(n_2220)
);

AND2x4_ASAP7_75t_L g2221 ( 
.A(n_2002),
.B(n_1014),
.Y(n_2221)
);

HB1xp67_ASAP7_75t_L g2222 ( 
.A(n_1971),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_1998),
.B(n_928),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_1970),
.Y(n_2224)
);

INVx2_ASAP7_75t_SL g2225 ( 
.A(n_2076),
.Y(n_2225)
);

NOR2xp33_ASAP7_75t_L g2226 ( 
.A(n_2054),
.B(n_929),
.Y(n_2226)
);

INVx5_ASAP7_75t_L g2227 ( 
.A(n_1959),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2039),
.Y(n_2228)
);

INVxp67_ASAP7_75t_L g2229 ( 
.A(n_2029),
.Y(n_2229)
);

AOI22xp5_ASAP7_75t_L g2230 ( 
.A1(n_2058),
.A2(n_932),
.B1(n_936),
.B2(n_930),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1980),
.Y(n_2231)
);

INVx2_ASAP7_75t_SL g2232 ( 
.A(n_2080),
.Y(n_2232)
);

INVxp67_ASAP7_75t_L g2233 ( 
.A(n_2042),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1995),
.Y(n_2234)
);

NAND2xp33_ASAP7_75t_SL g2235 ( 
.A(n_2132),
.B(n_2059),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_SL g2236 ( 
.A(n_2207),
.B(n_2001),
.Y(n_2236)
);

NAND2xp33_ASAP7_75t_SL g2237 ( 
.A(n_2160),
.B(n_2061),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_2104),
.B(n_2026),
.Y(n_2238)
);

NAND2xp33_ASAP7_75t_SL g2239 ( 
.A(n_2162),
.B(n_2065),
.Y(n_2239)
);

NAND2xp33_ASAP7_75t_SL g2240 ( 
.A(n_2087),
.B(n_1953),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_SL g2241 ( 
.A(n_2157),
.B(n_2056),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_SL g2242 ( 
.A(n_2233),
.B(n_2011),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_SL g2243 ( 
.A(n_2111),
.B(n_2068),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_SL g2244 ( 
.A(n_2118),
.B(n_2037),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_SL g2245 ( 
.A(n_2095),
.B(n_2038),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_SL g2246 ( 
.A(n_2098),
.B(n_2046),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_SL g2247 ( 
.A(n_2215),
.B(n_2048),
.Y(n_2247)
);

NAND2xp33_ASAP7_75t_SL g2248 ( 
.A(n_2187),
.B(n_1990),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_2128),
.B(n_2057),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_SL g2250 ( 
.A(n_2220),
.B(n_2066),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_SL g2251 ( 
.A(n_2176),
.B(n_1959),
.Y(n_2251)
);

AND2x4_ASAP7_75t_L g2252 ( 
.A(n_2138),
.B(n_2145),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2101),
.B(n_2055),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_SL g2254 ( 
.A(n_2084),
.B(n_1959),
.Y(n_2254)
);

NAND2xp33_ASAP7_75t_SL g2255 ( 
.A(n_2187),
.B(n_1990),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_SL g2256 ( 
.A(n_2158),
.B(n_1959),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_SL g2257 ( 
.A(n_2183),
.B(n_1959),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_SL g2258 ( 
.A(n_2228),
.B(n_1977),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2219),
.B(n_1999),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_SL g2260 ( 
.A(n_2136),
.B(n_1945),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_SL g2261 ( 
.A(n_2229),
.B(n_1948),
.Y(n_2261)
);

NAND2xp33_ASAP7_75t_SL g2262 ( 
.A(n_2122),
.B(n_1961),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2135),
.B(n_2025),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_SL g2264 ( 
.A(n_2144),
.B(n_1962),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_SL g2265 ( 
.A(n_2144),
.B(n_1970),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_SL g2266 ( 
.A(n_2144),
.B(n_1974),
.Y(n_2266)
);

NAND2xp33_ASAP7_75t_SL g2267 ( 
.A(n_2122),
.B(n_1975),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_SL g2268 ( 
.A(n_2225),
.B(n_1974),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_SL g2269 ( 
.A(n_2105),
.B(n_1996),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_SL g2270 ( 
.A(n_2082),
.B(n_2013),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_SL g2271 ( 
.A(n_2232),
.B(n_1934),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_SL g2272 ( 
.A(n_2120),
.B(n_1963),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_SL g2273 ( 
.A(n_2119),
.B(n_1978),
.Y(n_2273)
);

NAND2xp33_ASAP7_75t_SL g2274 ( 
.A(n_2122),
.B(n_1965),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_SL g2275 ( 
.A(n_2189),
.B(n_852),
.Y(n_2275)
);

NAND2xp33_ASAP7_75t_SL g2276 ( 
.A(n_2126),
.B(n_854),
.Y(n_2276)
);

NAND2xp33_ASAP7_75t_SL g2277 ( 
.A(n_2126),
.B(n_854),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_SL g2278 ( 
.A(n_2103),
.B(n_855),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_2085),
.B(n_1016),
.Y(n_2279)
);

AND2x2_ASAP7_75t_SL g2280 ( 
.A(n_2226),
.B(n_2166),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_SL g2281 ( 
.A(n_2103),
.B(n_855),
.Y(n_2281)
);

NOR2xp33_ASAP7_75t_L g2282 ( 
.A(n_2121),
.B(n_940),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_SL g2283 ( 
.A(n_2103),
.B(n_856),
.Y(n_2283)
);

NAND2xp33_ASAP7_75t_SL g2284 ( 
.A(n_2126),
.B(n_856),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_SL g2285 ( 
.A(n_2103),
.B(n_857),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_SL g2286 ( 
.A(n_2201),
.B(n_857),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_SL g2287 ( 
.A(n_2081),
.B(n_858),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_SL g2288 ( 
.A(n_2195),
.B(n_858),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_SL g2289 ( 
.A(n_2202),
.B(n_859),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_SL g2290 ( 
.A(n_2222),
.B(n_859),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_SL g2291 ( 
.A(n_2093),
.B(n_2159),
.Y(n_2291)
);

NAND2xp33_ASAP7_75t_SL g2292 ( 
.A(n_2110),
.B(n_860),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_SL g2293 ( 
.A(n_2163),
.B(n_860),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_SL g2294 ( 
.A(n_2164),
.B(n_861),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_2170),
.B(n_907),
.Y(n_2295)
);

AND2x4_ASAP7_75t_L g2296 ( 
.A(n_2147),
.B(n_1019),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_SL g2297 ( 
.A(n_2182),
.B(n_861),
.Y(n_2297)
);

NAND2xp33_ASAP7_75t_SL g2298 ( 
.A(n_2086),
.B(n_862),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_SL g2299 ( 
.A(n_2143),
.B(n_2150),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_SL g2300 ( 
.A(n_2152),
.B(n_867),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_SL g2301 ( 
.A(n_2094),
.B(n_867),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_SL g2302 ( 
.A(n_2094),
.B(n_869),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_SL g2303 ( 
.A(n_2094),
.B(n_869),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_SL g2304 ( 
.A(n_2148),
.B(n_870),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_SL g2305 ( 
.A(n_2168),
.B(n_870),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_SL g2306 ( 
.A(n_2185),
.B(n_873),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_SL g2307 ( 
.A(n_2169),
.B(n_873),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2091),
.B(n_2175),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_2178),
.B(n_1020),
.Y(n_2309)
);

NAND2xp33_ASAP7_75t_SL g2310 ( 
.A(n_2088),
.B(n_877),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_SL g2311 ( 
.A(n_2181),
.B(n_2191),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_SL g2312 ( 
.A(n_2099),
.B(n_877),
.Y(n_2312)
);

NAND2xp33_ASAP7_75t_SL g2313 ( 
.A(n_2100),
.B(n_879),
.Y(n_2313)
);

NAND2xp33_ASAP7_75t_SL g2314 ( 
.A(n_2108),
.B(n_879),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_SL g2315 ( 
.A(n_2109),
.B(n_880),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_SL g2316 ( 
.A(n_2114),
.B(n_880),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_SL g2317 ( 
.A(n_2188),
.B(n_882),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2184),
.B(n_1030),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_SL g2319 ( 
.A(n_2117),
.B(n_882),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_SL g2320 ( 
.A(n_2149),
.B(n_1081),
.Y(n_2320)
);

OR2x2_ASAP7_75t_L g2321 ( 
.A(n_2198),
.B(n_1081),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_SL g2322 ( 
.A(n_2149),
.B(n_1301),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_SL g2323 ( 
.A(n_2153),
.B(n_1301),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_SL g2324 ( 
.A(n_2153),
.B(n_1302),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_SL g2325 ( 
.A(n_2173),
.B(n_1302),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_SL g2326 ( 
.A(n_2113),
.B(n_1303),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_SL g2327 ( 
.A(n_2125),
.B(n_1303),
.Y(n_2327)
);

AND2x4_ASAP7_75t_L g2328 ( 
.A(n_2186),
.B(n_1033),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_2161),
.B(n_1035),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_SL g2330 ( 
.A(n_2127),
.B(n_1306),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_SL g2331 ( 
.A(n_2137),
.B(n_1306),
.Y(n_2331)
);

NAND2xp33_ASAP7_75t_SL g2332 ( 
.A(n_2097),
.B(n_1309),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_SL g2333 ( 
.A(n_2139),
.B(n_1309),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_SL g2334 ( 
.A(n_2142),
.B(n_1315),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_SL g2335 ( 
.A(n_2124),
.B(n_2155),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_SL g2336 ( 
.A(n_2083),
.B(n_1315),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_SL g2337 ( 
.A(n_2223),
.B(n_2180),
.Y(n_2337)
);

AND2x4_ASAP7_75t_L g2338 ( 
.A(n_2211),
.B(n_1036),
.Y(n_2338)
);

NAND2xp33_ASAP7_75t_SL g2339 ( 
.A(n_2090),
.B(n_1316),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_SL g2340 ( 
.A(n_2212),
.B(n_1316),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_SL g2341 ( 
.A(n_2213),
.B(n_1319),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_SL g2342 ( 
.A(n_2171),
.B(n_1319),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_SL g2343 ( 
.A(n_2130),
.B(n_1320),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_SL g2344 ( 
.A(n_2131),
.B(n_1320),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_SL g2345 ( 
.A(n_2134),
.B(n_1347),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_SL g2346 ( 
.A(n_2140),
.B(n_1347),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_SL g2347 ( 
.A(n_2116),
.B(n_1348),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_SL g2348 ( 
.A(n_2203),
.B(n_1348),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_SL g2349 ( 
.A(n_2208),
.B(n_931),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_SL g2350 ( 
.A(n_2154),
.B(n_931),
.Y(n_2350)
);

AND2x2_ASAP7_75t_L g2351 ( 
.A(n_2199),
.B(n_931),
.Y(n_2351)
);

NAND2xp33_ASAP7_75t_SL g2352 ( 
.A(n_2129),
.B(n_1228),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_SL g2353 ( 
.A(n_2151),
.B(n_955),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2205),
.B(n_1038),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_SL g2355 ( 
.A(n_2172),
.B(n_955),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_SL g2356 ( 
.A(n_2174),
.B(n_2193),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_SL g2357 ( 
.A(n_2197),
.B(n_2217),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_SL g2358 ( 
.A(n_2230),
.B(n_955),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_SL g2359 ( 
.A(n_2209),
.B(n_990),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_SL g2360 ( 
.A(n_2192),
.B(n_990),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_SL g2361 ( 
.A(n_2190),
.B(n_990),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_SL g2362 ( 
.A(n_2199),
.B(n_1052),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_2210),
.B(n_1050),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_SL g2364 ( 
.A(n_2227),
.B(n_1052),
.Y(n_2364)
);

NOR2xp33_ASAP7_75t_L g2365 ( 
.A(n_2196),
.B(n_941),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_SL g2366 ( 
.A(n_2227),
.B(n_2231),
.Y(n_2366)
);

NAND2xp33_ASAP7_75t_SL g2367 ( 
.A(n_2167),
.B(n_1260),
.Y(n_2367)
);

NAND2xp33_ASAP7_75t_SL g2368 ( 
.A(n_2194),
.B(n_1260),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2141),
.B(n_1053),
.Y(n_2369)
);

NAND2xp33_ASAP7_75t_SL g2370 ( 
.A(n_2224),
.B(n_1263),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_SL g2371 ( 
.A(n_2227),
.B(n_1052),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_SL g2372 ( 
.A(n_2234),
.B(n_1099),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_SL g2373 ( 
.A(n_2218),
.B(n_1099),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_2107),
.B(n_1058),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_SL g2375 ( 
.A(n_2218),
.B(n_1099),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_2179),
.B(n_1179),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_SL g2377 ( 
.A(n_2221),
.B(n_1179),
.Y(n_2377)
);

NAND2xp33_ASAP7_75t_SL g2378 ( 
.A(n_2089),
.B(n_1263),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_SL g2379 ( 
.A(n_2221),
.B(n_1179),
.Y(n_2379)
);

NAND2xp33_ASAP7_75t_SL g2380 ( 
.A(n_2092),
.B(n_1283),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_SL g2381 ( 
.A(n_2106),
.B(n_1280),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2123),
.B(n_1061),
.Y(n_2382)
);

AND2x4_ASAP7_75t_L g2383 ( 
.A(n_2156),
.B(n_1064),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2216),
.B(n_1065),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_2096),
.B(n_1067),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2200),
.B(n_2156),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_SL g2387 ( 
.A(n_2112),
.B(n_1280),
.Y(n_2387)
);

NAND2xp33_ASAP7_75t_SL g2388 ( 
.A(n_2214),
.B(n_1283),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2308),
.B(n_2177),
.Y(n_2389)
);

OAI22xp5_ASAP7_75t_L g2390 ( 
.A1(n_2280),
.A2(n_2206),
.B1(n_2204),
.B2(n_2102),
.Y(n_2390)
);

HB1xp67_ASAP7_75t_L g2391 ( 
.A(n_2335),
.Y(n_2391)
);

AND2x2_ASAP7_75t_L g2392 ( 
.A(n_2295),
.B(n_2156),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_2249),
.B(n_2238),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_2253),
.B(n_2133),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2236),
.B(n_944),
.Y(n_2395)
);

INVx2_ASAP7_75t_SL g2396 ( 
.A(n_2296),
.Y(n_2396)
);

BUFx12f_ASAP7_75t_L g2397 ( 
.A(n_2296),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2291),
.Y(n_2398)
);

OR2x6_ASAP7_75t_L g2399 ( 
.A(n_2251),
.B(n_2165),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_SL g2400 ( 
.A(n_2235),
.B(n_2146),
.Y(n_2400)
);

CKINVDCx8_ASAP7_75t_R g2401 ( 
.A(n_2252),
.Y(n_2401)
);

AND2x2_ASAP7_75t_SL g2402 ( 
.A(n_2282),
.B(n_2146),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2299),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_2241),
.B(n_946),
.Y(n_2404)
);

CKINVDCx8_ASAP7_75t_R g2405 ( 
.A(n_2252),
.Y(n_2405)
);

HB1xp67_ASAP7_75t_L g2406 ( 
.A(n_2261),
.Y(n_2406)
);

CKINVDCx5p33_ASAP7_75t_R g2407 ( 
.A(n_2244),
.Y(n_2407)
);

INVx1_ASAP7_75t_SL g2408 ( 
.A(n_2351),
.Y(n_2408)
);

HB1xp67_ASAP7_75t_L g2409 ( 
.A(n_2264),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_SL g2410 ( 
.A(n_2237),
.B(n_2115),
.Y(n_2410)
);

AND2x4_ASAP7_75t_L g2411 ( 
.A(n_2265),
.B(n_767),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2242),
.B(n_950),
.Y(n_2412)
);

AND3x1_ASAP7_75t_SL g2413 ( 
.A(n_2243),
.B(n_1083),
.C(n_1078),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_SL g2414 ( 
.A(n_2246),
.B(n_1280),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_2279),
.B(n_952),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_2328),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2328),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_2338),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2338),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2354),
.B(n_954),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2263),
.B(n_958),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2309),
.B(n_963),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2259),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2318),
.B(n_968),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2329),
.B(n_2245),
.Y(n_2425)
);

NOR2xp67_ASAP7_75t_L g2426 ( 
.A(n_2258),
.B(n_768),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2321),
.B(n_969),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_2268),
.Y(n_2428)
);

BUFx2_ASAP7_75t_L g2429 ( 
.A(n_2276),
.Y(n_2429)
);

BUFx2_ASAP7_75t_L g2430 ( 
.A(n_2277),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2311),
.B(n_970),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2374),
.Y(n_2432)
);

INVx3_ASAP7_75t_L g2433 ( 
.A(n_2383),
.Y(n_2433)
);

OAI22xp5_ASAP7_75t_L g2434 ( 
.A1(n_2357),
.A2(n_2287),
.B1(n_2273),
.B2(n_2250),
.Y(n_2434)
);

A2O1A1Ixp33_ASAP7_75t_L g2435 ( 
.A1(n_2239),
.A2(n_1305),
.B(n_1307),
.C(n_1289),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_SL g2436 ( 
.A(n_2240),
.B(n_1339),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2247),
.B(n_972),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2356),
.Y(n_2438)
);

BUFx4f_ASAP7_75t_SL g2439 ( 
.A(n_2270),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2337),
.B(n_974),
.Y(n_2440)
);

AND2x2_ASAP7_75t_SL g2441 ( 
.A(n_2386),
.B(n_1289),
.Y(n_2441)
);

NOR2xp33_ASAP7_75t_L g2442 ( 
.A(n_2304),
.B(n_975),
.Y(n_2442)
);

OAI21xp5_ASAP7_75t_L g2443 ( 
.A1(n_2369),
.A2(n_1090),
.B(n_1084),
.Y(n_2443)
);

INVx3_ASAP7_75t_L g2444 ( 
.A(n_2383),
.Y(n_2444)
);

NAND3xp33_ASAP7_75t_L g2445 ( 
.A(n_2358),
.B(n_978),
.C(n_977),
.Y(n_2445)
);

AND3x1_ASAP7_75t_SL g2446 ( 
.A(n_2388),
.B(n_1100),
.C(n_1095),
.Y(n_2446)
);

AOI22xp5_ASAP7_75t_L g2447 ( 
.A1(n_2272),
.A2(n_2332),
.B1(n_2360),
.B2(n_2342),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2305),
.B(n_979),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2366),
.Y(n_2449)
);

OAI221xp5_ASAP7_75t_L g2450 ( 
.A1(n_2365),
.A2(n_1114),
.B1(n_1123),
.B2(n_1108),
.C(n_1101),
.Y(n_2450)
);

AND2x2_ASAP7_75t_L g2451 ( 
.A(n_2376),
.B(n_1126),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2385),
.Y(n_2452)
);

BUFx12f_ASAP7_75t_L g2453 ( 
.A(n_2284),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2293),
.B(n_1129),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_2269),
.Y(n_2455)
);

AND2x2_ASAP7_75t_L g2456 ( 
.A(n_2294),
.B(n_1130),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2260),
.Y(n_2457)
);

BUFx8_ASAP7_75t_SL g2458 ( 
.A(n_2363),
.Y(n_2458)
);

AND3x1_ASAP7_75t_SL g2459 ( 
.A(n_2352),
.B(n_1146),
.C(n_1142),
.Y(n_2459)
);

NAND2xp33_ASAP7_75t_L g2460 ( 
.A(n_2248),
.B(n_980),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_2297),
.B(n_2288),
.Y(n_2461)
);

OAI22xp5_ASAP7_75t_L g2462 ( 
.A1(n_2325),
.A2(n_983),
.B1(n_984),
.B2(n_981),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2266),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2256),
.Y(n_2464)
);

AOI211xp5_ASAP7_75t_L g2465 ( 
.A1(n_2361),
.A2(n_1149),
.B(n_1161),
.C(n_1148),
.Y(n_2465)
);

AOI21xp33_ASAP7_75t_L g2466 ( 
.A1(n_2359),
.A2(n_1169),
.B(n_1168),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_2257),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_2271),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2289),
.B(n_986),
.Y(n_2469)
);

HB1xp67_ASAP7_75t_L g2470 ( 
.A(n_2254),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2384),
.Y(n_2471)
);

OR2x6_ASAP7_75t_L g2472 ( 
.A(n_2278),
.B(n_1305),
.Y(n_2472)
);

INVx2_ASAP7_75t_L g2473 ( 
.A(n_2382),
.Y(n_2473)
);

NOR2xp33_ASAP7_75t_R g2474 ( 
.A(n_2255),
.B(n_769),
.Y(n_2474)
);

AND2x2_ASAP7_75t_L g2475 ( 
.A(n_2300),
.B(n_1172),
.Y(n_2475)
);

AOI22xp5_ASAP7_75t_L g2476 ( 
.A1(n_2298),
.A2(n_988),
.B1(n_989),
.B2(n_987),
.Y(n_2476)
);

AND2x4_ASAP7_75t_L g2477 ( 
.A(n_2336),
.B(n_770),
.Y(n_2477)
);

INVx3_ASAP7_75t_L g2478 ( 
.A(n_2262),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2306),
.B(n_993),
.Y(n_2479)
);

INVx5_ASAP7_75t_L g2480 ( 
.A(n_2267),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_2281),
.Y(n_2481)
);

AND2x2_ASAP7_75t_L g2482 ( 
.A(n_2312),
.B(n_2315),
.Y(n_2482)
);

AND2x2_ASAP7_75t_L g2483 ( 
.A(n_2316),
.B(n_1173),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2380),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2378),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_2307),
.B(n_995),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2343),
.Y(n_2487)
);

CKINVDCx5p33_ASAP7_75t_R g2488 ( 
.A(n_2339),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2344),
.Y(n_2489)
);

INVx2_ASAP7_75t_L g2490 ( 
.A(n_2283),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2320),
.B(n_998),
.Y(n_2491)
);

OAI22xp5_ASAP7_75t_SL g2492 ( 
.A1(n_2381),
.A2(n_1205),
.B1(n_1207),
.B2(n_1202),
.Y(n_2492)
);

OR2x6_ASAP7_75t_SL g2493 ( 
.A(n_2362),
.B(n_999),
.Y(n_2493)
);

AND2x2_ASAP7_75t_L g2494 ( 
.A(n_2319),
.B(n_1208),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2285),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2326),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2322),
.B(n_1001),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_SL g2498 ( 
.A(n_2364),
.B(n_1340),
.Y(n_2498)
);

AND2x2_ASAP7_75t_L g2499 ( 
.A(n_2323),
.B(n_1209),
.Y(n_2499)
);

AND3x1_ASAP7_75t_SL g2500 ( 
.A(n_2367),
.B(n_1211),
.C(n_1210),
.Y(n_2500)
);

AND2x2_ASAP7_75t_L g2501 ( 
.A(n_2324),
.B(n_1215),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_2286),
.B(n_1003),
.Y(n_2502)
);

NAND3xp33_ASAP7_75t_SL g2503 ( 
.A(n_2350),
.B(n_1008),
.C(n_1006),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2275),
.B(n_1005),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2317),
.B(n_1017),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2345),
.Y(n_2506)
);

INVx2_ASAP7_75t_SL g2507 ( 
.A(n_2290),
.Y(n_2507)
);

AND2x2_ASAP7_75t_L g2508 ( 
.A(n_2327),
.B(n_1220),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_2371),
.B(n_1018),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_L g2510 ( 
.A(n_2346),
.B(n_1022),
.Y(n_2510)
);

AOI22x1_ASAP7_75t_L g2511 ( 
.A1(n_2370),
.A2(n_1311),
.B1(n_1335),
.B2(n_1307),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2348),
.Y(n_2512)
);

OAI21xp5_ASAP7_75t_L g2513 ( 
.A1(n_2372),
.A2(n_1224),
.B(n_1223),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2330),
.Y(n_2514)
);

CKINVDCx5p33_ASAP7_75t_R g2515 ( 
.A(n_2368),
.Y(n_2515)
);

AND2x2_ASAP7_75t_L g2516 ( 
.A(n_2331),
.B(n_1226),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_SL g2517 ( 
.A(n_2349),
.B(n_1343),
.Y(n_2517)
);

AND2x4_ASAP7_75t_L g2518 ( 
.A(n_2333),
.B(n_2340),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_SL g2519 ( 
.A(n_2347),
.B(n_1344),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_2334),
.Y(n_2520)
);

AND2x2_ASAP7_75t_L g2521 ( 
.A(n_2341),
.B(n_2301),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2274),
.Y(n_2522)
);

OAI21xp5_ASAP7_75t_L g2523 ( 
.A1(n_2353),
.A2(n_1232),
.B(n_1229),
.Y(n_2523)
);

NAND2xp33_ASAP7_75t_SL g2524 ( 
.A(n_2373),
.B(n_1350),
.Y(n_2524)
);

AND2x2_ASAP7_75t_L g2525 ( 
.A(n_2302),
.B(n_1233),
.Y(n_2525)
);

CKINVDCx5p33_ASAP7_75t_R g2526 ( 
.A(n_2292),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2355),
.Y(n_2527)
);

OAI22xp5_ASAP7_75t_SL g2528 ( 
.A1(n_2310),
.A2(n_1245),
.B1(n_1254),
.B2(n_1243),
.Y(n_2528)
);

NOR2xp33_ASAP7_75t_SL g2529 ( 
.A(n_2375),
.B(n_1025),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2377),
.B(n_1024),
.Y(n_2530)
);

AOI22x1_ASAP7_75t_L g2531 ( 
.A1(n_2452),
.A2(n_1335),
.B1(n_1341),
.B2(n_1311),
.Y(n_2531)
);

NAND2x1p5_ASAP7_75t_L g2532 ( 
.A(n_2480),
.B(n_2387),
.Y(n_2532)
);

INVx2_ASAP7_75t_SL g2533 ( 
.A(n_2397),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2468),
.Y(n_2534)
);

NAND2x1p5_ASAP7_75t_L g2535 ( 
.A(n_2480),
.B(n_2379),
.Y(n_2535)
);

OAI21x1_ASAP7_75t_L g2536 ( 
.A1(n_2410),
.A2(n_2303),
.B(n_1341),
.Y(n_2536)
);

INVx1_ASAP7_75t_SL g2537 ( 
.A(n_2408),
.Y(n_2537)
);

NAND2x1p5_ASAP7_75t_L g2538 ( 
.A(n_2480),
.B(n_1332),
.Y(n_2538)
);

HB1xp67_ASAP7_75t_L g2539 ( 
.A(n_2391),
.Y(n_2539)
);

OAI21xp5_ASAP7_75t_L g2540 ( 
.A1(n_2447),
.A2(n_2314),
.B(n_2313),
.Y(n_2540)
);

HB1xp67_ASAP7_75t_L g2541 ( 
.A(n_2406),
.Y(n_2541)
);

CKINVDCx5p33_ASAP7_75t_R g2542 ( 
.A(n_2458),
.Y(n_2542)
);

BUFx12f_ASAP7_75t_L g2543 ( 
.A(n_2453),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2403),
.Y(n_2544)
);

OAI21xp5_ASAP7_75t_L g2545 ( 
.A1(n_2447),
.A2(n_1314),
.B(n_1265),
.Y(n_2545)
);

AO21x2_ASAP7_75t_L g2546 ( 
.A1(n_2400),
.A2(n_1267),
.B(n_1262),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2398),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_2441),
.B(n_1271),
.Y(n_2548)
);

INVx6_ASAP7_75t_L g2549 ( 
.A(n_2402),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2428),
.Y(n_2550)
);

BUFx6f_ASAP7_75t_L g2551 ( 
.A(n_2401),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2393),
.B(n_1026),
.Y(n_2552)
);

OAI21x1_ASAP7_75t_L g2553 ( 
.A1(n_2464),
.A2(n_1286),
.B(n_1273),
.Y(n_2553)
);

AOI21xp5_ASAP7_75t_L g2554 ( 
.A1(n_2425),
.A2(n_1291),
.B(n_1287),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2455),
.Y(n_2555)
);

INVx2_ASAP7_75t_SL g2556 ( 
.A(n_2396),
.Y(n_2556)
);

INVx4_ASAP7_75t_L g2557 ( 
.A(n_2478),
.Y(n_2557)
);

OAI21x1_ASAP7_75t_L g2558 ( 
.A1(n_2467),
.A2(n_1297),
.B(n_1295),
.Y(n_2558)
);

INVx6_ASAP7_75t_L g2559 ( 
.A(n_2518),
.Y(n_2559)
);

AO21x1_ASAP7_75t_L g2560 ( 
.A1(n_2434),
.A2(n_1308),
.B(n_1300),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2470),
.Y(n_2561)
);

OAI21x1_ASAP7_75t_L g2562 ( 
.A1(n_2484),
.A2(n_1318),
.B(n_1313),
.Y(n_2562)
);

INVx1_ASAP7_75t_SL g2563 ( 
.A(n_2407),
.Y(n_2563)
);

INVx4_ASAP7_75t_L g2564 ( 
.A(n_2478),
.Y(n_2564)
);

INVx3_ASAP7_75t_L g2565 ( 
.A(n_2433),
.Y(n_2565)
);

BUFx6f_ASAP7_75t_SL g2566 ( 
.A(n_2518),
.Y(n_2566)
);

NOR2xp33_ASAP7_75t_L g2567 ( 
.A(n_2394),
.B(n_1027),
.Y(n_2567)
);

BUFx6f_ASAP7_75t_L g2568 ( 
.A(n_2405),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2423),
.Y(n_2569)
);

OAI21xp5_ASAP7_75t_L g2570 ( 
.A1(n_2445),
.A2(n_1324),
.B(n_1322),
.Y(n_2570)
);

BUFx3_ASAP7_75t_L g2571 ( 
.A(n_2439),
.Y(n_2571)
);

INVx6_ASAP7_75t_L g2572 ( 
.A(n_2411),
.Y(n_2572)
);

INVx1_ASAP7_75t_SL g2573 ( 
.A(n_2389),
.Y(n_2573)
);

AND2x4_ASAP7_75t_L g2574 ( 
.A(n_2449),
.B(n_771),
.Y(n_2574)
);

OAI21x1_ASAP7_75t_L g2575 ( 
.A1(n_2390),
.A2(n_1326),
.B(n_1325),
.Y(n_2575)
);

OAI21x1_ASAP7_75t_L g2576 ( 
.A1(n_2522),
.A2(n_1338),
.B(n_1333),
.Y(n_2576)
);

AO21x2_ASAP7_75t_L g2577 ( 
.A1(n_2436),
.A2(n_1342),
.B(n_1085),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2399),
.Y(n_2578)
);

BUFx3_ASAP7_75t_L g2579 ( 
.A(n_2507),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2399),
.Y(n_2580)
);

INVx2_ASAP7_75t_L g2581 ( 
.A(n_2438),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_2457),
.Y(n_2582)
);

AO21x2_ASAP7_75t_L g2583 ( 
.A1(n_2426),
.A2(n_1070),
.B(n_2),
.Y(n_2583)
);

BUFx2_ASAP7_75t_R g2584 ( 
.A(n_2488),
.Y(n_2584)
);

BUFx3_ASAP7_75t_L g2585 ( 
.A(n_2526),
.Y(n_2585)
);

OAI21xp5_ASAP7_75t_L g2586 ( 
.A1(n_2445),
.A2(n_1032),
.B(n_1031),
.Y(n_2586)
);

HB1xp67_ASAP7_75t_L g2587 ( 
.A(n_2409),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2473),
.Y(n_2588)
);

INVx2_ASAP7_75t_SL g2589 ( 
.A(n_2433),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_2416),
.Y(n_2590)
);

BUFx4_ASAP7_75t_SL g2591 ( 
.A(n_2429),
.Y(n_2591)
);

OAI22x1_ASAP7_75t_L g2592 ( 
.A1(n_2414),
.A2(n_1037),
.B1(n_1039),
.B2(n_1034),
.Y(n_2592)
);

BUFx6f_ASAP7_75t_SL g2593 ( 
.A(n_2477),
.Y(n_2593)
);

BUFx6f_ASAP7_75t_L g2594 ( 
.A(n_2444),
.Y(n_2594)
);

BUFx3_ASAP7_75t_L g2595 ( 
.A(n_2444),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2432),
.B(n_1298),
.Y(n_2596)
);

CKINVDCx8_ASAP7_75t_R g2597 ( 
.A(n_2515),
.Y(n_2597)
);

INVx5_ASAP7_75t_L g2598 ( 
.A(n_2472),
.Y(n_2598)
);

AO21x2_ASAP7_75t_L g2599 ( 
.A1(n_2426),
.A2(n_1041),
.B(n_1040),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2399),
.Y(n_2600)
);

BUFx3_ASAP7_75t_L g2601 ( 
.A(n_2430),
.Y(n_2601)
);

INVx3_ASAP7_75t_L g2602 ( 
.A(n_2418),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2463),
.Y(n_2603)
);

AND2x2_ASAP7_75t_L g2604 ( 
.A(n_2417),
.B(n_776),
.Y(n_2604)
);

OAI21xp5_ASAP7_75t_L g2605 ( 
.A1(n_2443),
.A2(n_1044),
.B(n_1042),
.Y(n_2605)
);

INVxp67_ASAP7_75t_SL g2606 ( 
.A(n_2471),
.Y(n_2606)
);

INVx6_ASAP7_75t_L g2607 ( 
.A(n_2411),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2419),
.Y(n_2608)
);

INVx3_ASAP7_75t_L g2609 ( 
.A(n_2481),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_2490),
.B(n_1337),
.Y(n_2610)
);

NAND2x1p5_ASAP7_75t_L g2611 ( 
.A(n_2392),
.B(n_778),
.Y(n_2611)
);

OA21x2_ASAP7_75t_L g2612 ( 
.A1(n_2435),
.A2(n_1046),
.B(n_1045),
.Y(n_2612)
);

AO21x2_ASAP7_75t_L g2613 ( 
.A1(n_2485),
.A2(n_2),
.B(n_3),
.Y(n_2613)
);

OR2x6_ASAP7_75t_L g2614 ( 
.A(n_2477),
.B(n_781),
.Y(n_2614)
);

AND2x2_ASAP7_75t_L g2615 ( 
.A(n_2451),
.B(n_2487),
.Y(n_2615)
);

INVx2_ASAP7_75t_SL g2616 ( 
.A(n_2496),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2495),
.Y(n_2617)
);

BUFx2_ASAP7_75t_R g2618 ( 
.A(n_2493),
.Y(n_2618)
);

BUFx2_ASAP7_75t_R g2619 ( 
.A(n_2498),
.Y(n_2619)
);

OAI21x1_ASAP7_75t_L g2620 ( 
.A1(n_2511),
.A2(n_783),
.B(n_782),
.Y(n_2620)
);

HB1xp67_ASAP7_75t_L g2621 ( 
.A(n_2514),
.Y(n_2621)
);

INVx3_ASAP7_75t_L g2622 ( 
.A(n_2520),
.Y(n_2622)
);

OAI21xp5_ASAP7_75t_L g2623 ( 
.A1(n_2442),
.A2(n_1048),
.B(n_1047),
.Y(n_2623)
);

INVxp67_ASAP7_75t_SL g2624 ( 
.A(n_2489),
.Y(n_2624)
);

CKINVDCx20_ASAP7_75t_R g2625 ( 
.A(n_2524),
.Y(n_2625)
);

BUFx3_ASAP7_75t_L g2626 ( 
.A(n_2521),
.Y(n_2626)
);

INVx1_ASAP7_75t_SL g2627 ( 
.A(n_2461),
.Y(n_2627)
);

INVx3_ASAP7_75t_L g2628 ( 
.A(n_2506),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2512),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_L g2630 ( 
.A(n_2421),
.B(n_1292),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2395),
.Y(n_2631)
);

INVxp67_ASAP7_75t_SL g2632 ( 
.A(n_2460),
.Y(n_2632)
);

AO21x2_ASAP7_75t_L g2633 ( 
.A1(n_2474),
.A2(n_3),
.B(n_4),
.Y(n_2633)
);

OAI21x1_ASAP7_75t_L g2634 ( 
.A1(n_2527),
.A2(n_786),
.B(n_784),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2544),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2544),
.Y(n_2636)
);

OAI22xp5_ASAP7_75t_L g2637 ( 
.A1(n_2614),
.A2(n_2465),
.B1(n_2492),
.B2(n_2476),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2547),
.Y(n_2638)
);

BUFx6f_ASAP7_75t_L g2639 ( 
.A(n_2551),
.Y(n_2639)
);

AND2x2_ASAP7_75t_L g2640 ( 
.A(n_2626),
.B(n_2482),
.Y(n_2640)
);

BUFx12f_ASAP7_75t_L g2641 ( 
.A(n_2543),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2547),
.Y(n_2642)
);

OAI22xp33_ASAP7_75t_L g2643 ( 
.A1(n_2614),
.A2(n_2529),
.B1(n_2472),
.B2(n_2412),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2603),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2603),
.Y(n_2645)
);

INVx3_ASAP7_75t_L g2646 ( 
.A(n_2628),
.Y(n_2646)
);

AOI22xp33_ASAP7_75t_SL g2647 ( 
.A1(n_2593),
.A2(n_2529),
.B1(n_2492),
.B2(n_2528),
.Y(n_2647)
);

NAND2x1p5_ASAP7_75t_L g2648 ( 
.A(n_2557),
.B(n_2517),
.Y(n_2648)
);

AND2x2_ASAP7_75t_L g2649 ( 
.A(n_2627),
.B(n_2525),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2561),
.Y(n_2650)
);

OAI22xp5_ASAP7_75t_L g2651 ( 
.A1(n_2593),
.A2(n_2465),
.B1(n_2476),
.B2(n_2404),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2561),
.Y(n_2652)
);

INVx2_ASAP7_75t_SL g2653 ( 
.A(n_2579),
.Y(n_2653)
);

CKINVDCx5p33_ASAP7_75t_R g2654 ( 
.A(n_2542),
.Y(n_2654)
);

BUFx2_ASAP7_75t_SL g2655 ( 
.A(n_2566),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2569),
.Y(n_2656)
);

AOI22xp33_ASAP7_75t_L g2657 ( 
.A1(n_2540),
.A2(n_2560),
.B1(n_2633),
.B2(n_2545),
.Y(n_2657)
);

CKINVDCx11_ASAP7_75t_R g2658 ( 
.A(n_2597),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2581),
.Y(n_2659)
);

AOI22xp33_ASAP7_75t_L g2660 ( 
.A1(n_2633),
.A2(n_2528),
.B1(n_2503),
.B2(n_2466),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2569),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2621),
.Y(n_2662)
);

BUFx3_ASAP7_75t_L g2663 ( 
.A(n_2571),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2624),
.Y(n_2664)
);

AOI22xp33_ASAP7_75t_SL g2665 ( 
.A1(n_2566),
.A2(n_2513),
.B1(n_2472),
.B2(n_2450),
.Y(n_2665)
);

OAI22xp5_ASAP7_75t_L g2666 ( 
.A1(n_2598),
.A2(n_2440),
.B1(n_2431),
.B2(n_2509),
.Y(n_2666)
);

BUFx12f_ASAP7_75t_L g2667 ( 
.A(n_2551),
.Y(n_2667)
);

AOI22xp33_ASAP7_75t_SL g2668 ( 
.A1(n_2632),
.A2(n_2523),
.B1(n_2501),
.B2(n_2499),
.Y(n_2668)
);

INVx2_ASAP7_75t_L g2669 ( 
.A(n_2582),
.Y(n_2669)
);

INVx2_ASAP7_75t_SL g2670 ( 
.A(n_2591),
.Y(n_2670)
);

CKINVDCx20_ASAP7_75t_R g2671 ( 
.A(n_2625),
.Y(n_2671)
);

CKINVDCx6p67_ASAP7_75t_R g2672 ( 
.A(n_2585),
.Y(n_2672)
);

OAI22xp5_ASAP7_75t_L g2673 ( 
.A1(n_2598),
.A2(n_2437),
.B1(n_2530),
.B2(n_2519),
.Y(n_2673)
);

CKINVDCx11_ASAP7_75t_R g2674 ( 
.A(n_2551),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2629),
.Y(n_2675)
);

INVx1_ASAP7_75t_SL g2676 ( 
.A(n_2563),
.Y(n_2676)
);

AOI22xp33_ASAP7_75t_L g2677 ( 
.A1(n_2572),
.A2(n_2456),
.B1(n_2475),
.B2(n_2454),
.Y(n_2677)
);

BUFx10_ASAP7_75t_L g2678 ( 
.A(n_2549),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2608),
.Y(n_2679)
);

BUFx8_ASAP7_75t_SL g2680 ( 
.A(n_2568),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2534),
.Y(n_2681)
);

INVxp67_ASAP7_75t_SL g2682 ( 
.A(n_2541),
.Y(n_2682)
);

AOI21xp33_ASAP7_75t_L g2683 ( 
.A1(n_2631),
.A2(n_2420),
.B(n_2415),
.Y(n_2683)
);

INVx2_ASAP7_75t_L g2684 ( 
.A(n_2628),
.Y(n_2684)
);

CKINVDCx11_ASAP7_75t_R g2685 ( 
.A(n_2568),
.Y(n_2685)
);

BUFx12f_ASAP7_75t_L g2686 ( 
.A(n_2568),
.Y(n_2686)
);

CKINVDCx20_ASAP7_75t_R g2687 ( 
.A(n_2549),
.Y(n_2687)
);

OAI22xp5_ASAP7_75t_L g2688 ( 
.A1(n_2598),
.A2(n_2422),
.B1(n_2424),
.B2(n_2469),
.Y(n_2688)
);

BUFx10_ASAP7_75t_L g2689 ( 
.A(n_2533),
.Y(n_2689)
);

AOI22xp33_ASAP7_75t_L g2690 ( 
.A1(n_2572),
.A2(n_2494),
.B1(n_2483),
.B2(n_2508),
.Y(n_2690)
);

AOI22xp5_ASAP7_75t_L g2691 ( 
.A1(n_2607),
.A2(n_2631),
.B1(n_2559),
.B2(n_2546),
.Y(n_2691)
);

CKINVDCx5p33_ASAP7_75t_R g2692 ( 
.A(n_2584),
.Y(n_2692)
);

OAI22xp33_ASAP7_75t_L g2693 ( 
.A1(n_2573),
.A2(n_2448),
.B1(n_2486),
.B2(n_2427),
.Y(n_2693)
);

BUFx6f_ASAP7_75t_L g2694 ( 
.A(n_2594),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2534),
.Y(n_2695)
);

BUFx4f_ASAP7_75t_SL g2696 ( 
.A(n_2601),
.Y(n_2696)
);

OR2x2_ASAP7_75t_L g2697 ( 
.A(n_2539),
.B(n_2516),
.Y(n_2697)
);

CKINVDCx8_ASAP7_75t_R g2698 ( 
.A(n_2594),
.Y(n_2698)
);

AOI22xp33_ASAP7_75t_L g2699 ( 
.A1(n_2607),
.A2(n_2479),
.B1(n_2497),
.B2(n_2491),
.Y(n_2699)
);

BUFx4f_ASAP7_75t_L g2700 ( 
.A(n_2535),
.Y(n_2700)
);

AOI22xp33_ASAP7_75t_SL g2701 ( 
.A1(n_2559),
.A2(n_2413),
.B1(n_2462),
.B2(n_2502),
.Y(n_2701)
);

AOI22xp33_ASAP7_75t_SL g2702 ( 
.A1(n_2583),
.A2(n_2505),
.B1(n_2510),
.B2(n_2504),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2587),
.Y(n_2703)
);

INVx2_ASAP7_75t_L g2704 ( 
.A(n_2617),
.Y(n_2704)
);

AOI22xp33_ASAP7_75t_SL g2705 ( 
.A1(n_2583),
.A2(n_2500),
.B1(n_2459),
.B2(n_1057),
.Y(n_2705)
);

AOI22xp5_ASAP7_75t_L g2706 ( 
.A1(n_2546),
.A2(n_2446),
.B1(n_1062),
.B2(n_1069),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2617),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2606),
.B(n_1054),
.Y(n_2708)
);

INVx4_ASAP7_75t_SL g2709 ( 
.A(n_2615),
.Y(n_2709)
);

AOI22xp33_ASAP7_75t_SL g2710 ( 
.A1(n_2548),
.A2(n_1072),
.B1(n_1073),
.B2(n_1063),
.Y(n_2710)
);

AOI22xp33_ASAP7_75t_L g2711 ( 
.A1(n_2623),
.A2(n_2567),
.B1(n_2577),
.B2(n_2605),
.Y(n_2711)
);

OAI22xp33_ASAP7_75t_L g2712 ( 
.A1(n_2538),
.A2(n_1323),
.B1(n_1279),
.B2(n_1098),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2550),
.Y(n_2713)
);

CKINVDCx16_ASAP7_75t_R g2714 ( 
.A(n_2595),
.Y(n_2714)
);

INVx6_ASAP7_75t_L g2715 ( 
.A(n_2594),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2588),
.Y(n_2716)
);

HB1xp67_ASAP7_75t_L g2717 ( 
.A(n_2662),
.Y(n_2717)
);

AND2x2_ASAP7_75t_L g2718 ( 
.A(n_2682),
.B(n_2578),
.Y(n_2718)
);

OAI21x1_ASAP7_75t_L g2719 ( 
.A1(n_2691),
.A2(n_2575),
.B(n_2536),
.Y(n_2719)
);

INVx2_ASAP7_75t_SL g2720 ( 
.A(n_2696),
.Y(n_2720)
);

INVxp67_ASAP7_75t_SL g2721 ( 
.A(n_2664),
.Y(n_2721)
);

AOI22xp33_ASAP7_75t_L g2722 ( 
.A1(n_2637),
.A2(n_2612),
.B1(n_2599),
.B2(n_2577),
.Y(n_2722)
);

AOI221xp5_ASAP7_75t_L g2723 ( 
.A1(n_2683),
.A2(n_2570),
.B1(n_2554),
.B2(n_2586),
.C(n_2592),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2703),
.B(n_2622),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2659),
.B(n_2622),
.Y(n_2725)
);

AND2x4_ASAP7_75t_L g2726 ( 
.A(n_2709),
.B(n_2578),
.Y(n_2726)
);

OAI21x1_ASAP7_75t_L g2727 ( 
.A1(n_2657),
.A2(n_2620),
.B(n_2634),
.Y(n_2727)
);

AOI21xp5_ASAP7_75t_L g2728 ( 
.A1(n_2711),
.A2(n_2532),
.B(n_2612),
.Y(n_2728)
);

OAI22xp33_ASAP7_75t_SL g2729 ( 
.A1(n_2651),
.A2(n_2609),
.B1(n_2616),
.B2(n_2555),
.Y(n_2729)
);

HB1xp67_ASAP7_75t_L g2730 ( 
.A(n_2646),
.Y(n_2730)
);

BUFx3_ASAP7_75t_L g2731 ( 
.A(n_2680),
.Y(n_2731)
);

OAI21x1_ASAP7_75t_L g2732 ( 
.A1(n_2666),
.A2(n_2600),
.B(n_2580),
.Y(n_2732)
);

OR2x2_ASAP7_75t_L g2733 ( 
.A(n_2650),
.B(n_2652),
.Y(n_2733)
);

OA21x2_ASAP7_75t_L g2734 ( 
.A1(n_2635),
.A2(n_2600),
.B(n_2580),
.Y(n_2734)
);

OAI21xp5_ASAP7_75t_L g2735 ( 
.A1(n_2702),
.A2(n_2576),
.B(n_2552),
.Y(n_2735)
);

O2A1O1Ixp33_ASAP7_75t_L g2736 ( 
.A1(n_2643),
.A2(n_2630),
.B(n_2613),
.C(n_2596),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2669),
.B(n_2609),
.Y(n_2737)
);

OR2x2_ASAP7_75t_L g2738 ( 
.A(n_2697),
.B(n_2636),
.Y(n_2738)
);

OAI221xp5_ASAP7_75t_L g2739 ( 
.A1(n_2701),
.A2(n_2610),
.B1(n_2611),
.B2(n_2537),
.C(n_2556),
.Y(n_2739)
);

HB1xp67_ASAP7_75t_L g2740 ( 
.A(n_2646),
.Y(n_2740)
);

AO21x2_ASAP7_75t_L g2741 ( 
.A1(n_2688),
.A2(n_2613),
.B(n_2562),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2638),
.Y(n_2742)
);

AO21x2_ASAP7_75t_L g2743 ( 
.A1(n_2642),
.A2(n_2645),
.B(n_2644),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2656),
.Y(n_2744)
);

OR2x6_ASAP7_75t_L g2745 ( 
.A(n_2655),
.B(n_2557),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2661),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2681),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_2675),
.Y(n_2748)
);

OAI22xp33_ASAP7_75t_L g2749 ( 
.A1(n_2706),
.A2(n_2564),
.B1(n_2589),
.B2(n_2531),
.Y(n_2749)
);

AO21x2_ASAP7_75t_L g2750 ( 
.A1(n_2708),
.A2(n_2558),
.B(n_2553),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2695),
.Y(n_2751)
);

AOI21x1_ASAP7_75t_L g2752 ( 
.A1(n_2673),
.A2(n_2590),
.B(n_2574),
.Y(n_2752)
);

AND2x4_ASAP7_75t_L g2753 ( 
.A(n_2709),
.B(n_2565),
.Y(n_2753)
);

AO31x2_ASAP7_75t_L g2754 ( 
.A1(n_2707),
.A2(n_2564),
.A3(n_2531),
.B(n_2565),
.Y(n_2754)
);

O2A1O1Ixp33_ASAP7_75t_L g2755 ( 
.A1(n_2660),
.A2(n_2574),
.B(n_2602),
.C(n_2604),
.Y(n_2755)
);

INVx1_ASAP7_75t_SL g2756 ( 
.A(n_2676),
.Y(n_2756)
);

HB1xp67_ASAP7_75t_L g2757 ( 
.A(n_2684),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2713),
.B(n_2602),
.Y(n_2758)
);

OA21x2_ASAP7_75t_L g2759 ( 
.A1(n_2704),
.A2(n_1076),
.B(n_1074),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2679),
.Y(n_2760)
);

AOI21xp5_ASAP7_75t_L g2761 ( 
.A1(n_2693),
.A2(n_2619),
.B(n_2618),
.Y(n_2761)
);

A2O1A1Ixp33_ASAP7_75t_L g2762 ( 
.A1(n_2665),
.A2(n_1290),
.B(n_1294),
.C(n_1288),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2716),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_2649),
.B(n_1080),
.Y(n_2764)
);

AOI21xp5_ASAP7_75t_L g2765 ( 
.A1(n_2700),
.A2(n_1088),
.B(n_1082),
.Y(n_2765)
);

OAI211xp5_ASAP7_75t_L g2766 ( 
.A1(n_2647),
.A2(n_1091),
.B(n_1092),
.C(n_1089),
.Y(n_2766)
);

INVx2_ASAP7_75t_SL g2767 ( 
.A(n_2678),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2640),
.Y(n_2768)
);

HB1xp67_ASAP7_75t_L g2769 ( 
.A(n_2694),
.Y(n_2769)
);

OR2x6_ASAP7_75t_L g2770 ( 
.A(n_2670),
.B(n_788),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2694),
.Y(n_2771)
);

OR2x2_ASAP7_75t_L g2772 ( 
.A(n_2714),
.B(n_2653),
.Y(n_2772)
);

AOI22xp33_ASAP7_75t_L g2773 ( 
.A1(n_2668),
.A2(n_1096),
.B1(n_1103),
.B2(n_1094),
.Y(n_2773)
);

AO31x2_ASAP7_75t_L g2774 ( 
.A1(n_2705),
.A2(n_6),
.A3(n_4),
.B(n_5),
.Y(n_2774)
);

AND2x2_ASAP7_75t_L g2775 ( 
.A(n_2639),
.B(n_7),
.Y(n_2775)
);

AND2x2_ASAP7_75t_L g2776 ( 
.A(n_2639),
.B(n_7),
.Y(n_2776)
);

AOI22xp33_ASAP7_75t_L g2777 ( 
.A1(n_2710),
.A2(n_1107),
.B1(n_1111),
.B2(n_1106),
.Y(n_2777)
);

OAI22x1_ASAP7_75t_L g2778 ( 
.A1(n_2692),
.A2(n_1113),
.B1(n_1117),
.B2(n_1112),
.Y(n_2778)
);

OR2x2_ASAP7_75t_L g2779 ( 
.A(n_2639),
.B(n_8),
.Y(n_2779)
);

AOI221xp5_ASAP7_75t_L g2780 ( 
.A1(n_2712),
.A2(n_1124),
.B1(n_1125),
.B2(n_1122),
.C(n_1121),
.Y(n_2780)
);

BUFx2_ASAP7_75t_L g2781 ( 
.A(n_2687),
.Y(n_2781)
);

AND2x2_ASAP7_75t_L g2782 ( 
.A(n_2678),
.B(n_9),
.Y(n_2782)
);

OA21x2_ASAP7_75t_L g2783 ( 
.A1(n_2690),
.A2(n_1131),
.B(n_1127),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2694),
.Y(n_2784)
);

AOI22xp33_ASAP7_75t_L g2785 ( 
.A1(n_2677),
.A2(n_1134),
.B1(n_1135),
.B2(n_1132),
.Y(n_2785)
);

CKINVDCx5p33_ASAP7_75t_R g2786 ( 
.A(n_2658),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_L g2787 ( 
.A(n_2699),
.B(n_1137),
.Y(n_2787)
);

BUFx3_ASAP7_75t_L g2788 ( 
.A(n_2663),
.Y(n_2788)
);

AOI21xp5_ASAP7_75t_L g2789 ( 
.A1(n_2648),
.A2(n_1139),
.B(n_1138),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2715),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2715),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2733),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2744),
.Y(n_2793)
);

INVx5_ASAP7_75t_L g2794 ( 
.A(n_2770),
.Y(n_2794)
);

AOI22xp5_ASAP7_75t_L g2795 ( 
.A1(n_2739),
.A2(n_2667),
.B1(n_2686),
.B2(n_2672),
.Y(n_2795)
);

OAI22xp5_ASAP7_75t_L g2796 ( 
.A1(n_2761),
.A2(n_2698),
.B1(n_2671),
.B2(n_2641),
.Y(n_2796)
);

AOI221xp5_ASAP7_75t_L g2797 ( 
.A1(n_2736),
.A2(n_1144),
.B1(n_1145),
.B2(n_1143),
.C(n_1140),
.Y(n_2797)
);

OAI22xp33_ASAP7_75t_L g2798 ( 
.A1(n_2783),
.A2(n_2654),
.B1(n_2685),
.B2(n_2674),
.Y(n_2798)
);

INVx2_ASAP7_75t_L g2799 ( 
.A(n_2738),
.Y(n_2799)
);

INVx1_ASAP7_75t_SL g2800 ( 
.A(n_2756),
.Y(n_2800)
);

AOI221xp5_ASAP7_75t_L g2801 ( 
.A1(n_2787),
.A2(n_1152),
.B1(n_1153),
.B2(n_1151),
.C(n_1150),
.Y(n_2801)
);

INVx3_ASAP7_75t_L g2802 ( 
.A(n_2726),
.Y(n_2802)
);

AND2x2_ASAP7_75t_L g2803 ( 
.A(n_2768),
.B(n_2689),
.Y(n_2803)
);

BUFx6f_ASAP7_75t_L g2804 ( 
.A(n_2731),
.Y(n_2804)
);

AOI22xp5_ASAP7_75t_L g2805 ( 
.A1(n_2723),
.A2(n_2689),
.B1(n_1157),
.B2(n_1158),
.Y(n_2805)
);

AOI221xp5_ASAP7_75t_L g2806 ( 
.A1(n_2735),
.A2(n_1159),
.B1(n_1160),
.B2(n_1156),
.C(n_1154),
.Y(n_2806)
);

OAI21xp33_ASAP7_75t_L g2807 ( 
.A1(n_2722),
.A2(n_1163),
.B(n_1162),
.Y(n_2807)
);

AOI22xp33_ASAP7_75t_L g2808 ( 
.A1(n_2783),
.A2(n_1330),
.B1(n_1328),
.B2(n_1165),
.Y(n_2808)
);

AOI22xp33_ASAP7_75t_L g2809 ( 
.A1(n_2728),
.A2(n_1167),
.B1(n_1171),
.B2(n_1164),
.Y(n_2809)
);

OAI21x1_ASAP7_75t_L g2810 ( 
.A1(n_2732),
.A2(n_10),
.B(n_11),
.Y(n_2810)
);

AOI22xp33_ASAP7_75t_L g2811 ( 
.A1(n_2741),
.A2(n_2749),
.B1(n_2729),
.B2(n_2773),
.Y(n_2811)
);

AOI22xp33_ASAP7_75t_L g2812 ( 
.A1(n_2759),
.A2(n_2750),
.B1(n_2778),
.B2(n_2785),
.Y(n_2812)
);

OAI211xp5_ASAP7_75t_L g2813 ( 
.A1(n_2766),
.A2(n_1192),
.B(n_1206),
.C(n_1176),
.Y(n_2813)
);

OAI221xp5_ASAP7_75t_L g2814 ( 
.A1(n_2762),
.A2(n_1177),
.B1(n_1182),
.B2(n_1175),
.C(n_1174),
.Y(n_2814)
);

AOI22xp33_ASAP7_75t_L g2815 ( 
.A1(n_2759),
.A2(n_1285),
.B1(n_1321),
.B2(n_1284),
.Y(n_2815)
);

OAI211xp5_ASAP7_75t_L g2816 ( 
.A1(n_2780),
.A2(n_1201),
.B(n_1227),
.C(n_1188),
.Y(n_2816)
);

AOI22xp33_ASAP7_75t_L g2817 ( 
.A1(n_2770),
.A2(n_1186),
.B1(n_1189),
.B2(n_1185),
.Y(n_2817)
);

AOI22xp33_ASAP7_75t_L g2818 ( 
.A1(n_2767),
.A2(n_1257),
.B1(n_1261),
.B2(n_1256),
.Y(n_2818)
);

OAI22xp5_ASAP7_75t_L g2819 ( 
.A1(n_2755),
.A2(n_1194),
.B1(n_1195),
.B2(n_1190),
.Y(n_2819)
);

NOR2xp33_ASAP7_75t_SL g2820 ( 
.A(n_2786),
.B(n_1275),
.Y(n_2820)
);

NAND2xp5_ASAP7_75t_L g2821 ( 
.A(n_2724),
.B(n_1196),
.Y(n_2821)
);

AOI22xp33_ASAP7_75t_L g2822 ( 
.A1(n_2781),
.A2(n_1281),
.B1(n_1327),
.B2(n_1277),
.Y(n_2822)
);

AND2x2_ASAP7_75t_L g2823 ( 
.A(n_2717),
.B(n_2730),
.Y(n_2823)
);

INVx5_ASAP7_75t_SL g2824 ( 
.A(n_2745),
.Y(n_2824)
);

AOI22xp33_ASAP7_75t_SL g2825 ( 
.A1(n_2727),
.A2(n_1200),
.B1(n_1203),
.B2(n_1197),
.Y(n_2825)
);

OAI21x1_ASAP7_75t_L g2826 ( 
.A1(n_2719),
.A2(n_10),
.B(n_12),
.Y(n_2826)
);

NOR2xp33_ASAP7_75t_L g2827 ( 
.A(n_2772),
.B(n_1212),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2740),
.Y(n_2828)
);

AOI22xp5_ASAP7_75t_L g2829 ( 
.A1(n_2745),
.A2(n_1218),
.B1(n_1219),
.B2(n_1216),
.Y(n_2829)
);

INVx3_ASAP7_75t_L g2830 ( 
.A(n_2726),
.Y(n_2830)
);

NOR2x1_ASAP7_75t_L g2831 ( 
.A(n_2743),
.B(n_12),
.Y(n_2831)
);

AND2x4_ASAP7_75t_L g2832 ( 
.A(n_2718),
.B(n_2753),
.Y(n_2832)
);

OAI21xp5_ASAP7_75t_L g2833 ( 
.A1(n_2789),
.A2(n_1225),
.B(n_1222),
.Y(n_2833)
);

INVx2_ASAP7_75t_L g2834 ( 
.A(n_2744),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_2721),
.B(n_1230),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2793),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_L g2837 ( 
.A(n_2823),
.B(n_2757),
.Y(n_2837)
);

INVx2_ASAP7_75t_L g2838 ( 
.A(n_2834),
.Y(n_2838)
);

CKINVDCx6p67_ASAP7_75t_R g2839 ( 
.A(n_2794),
.Y(n_2839)
);

INVx2_ASAP7_75t_L g2840 ( 
.A(n_2828),
.Y(n_2840)
);

OR2x2_ASAP7_75t_L g2841 ( 
.A(n_2799),
.B(n_2760),
.Y(n_2841)
);

AND2x4_ASAP7_75t_L g2842 ( 
.A(n_2802),
.B(n_2753),
.Y(n_2842)
);

AND2x2_ASAP7_75t_L g2843 ( 
.A(n_2832),
.B(n_2769),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2792),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2831),
.Y(n_2845)
);

BUFx2_ASAP7_75t_L g2846 ( 
.A(n_2802),
.Y(n_2846)
);

AND2x2_ASAP7_75t_L g2847 ( 
.A(n_2830),
.B(n_2734),
.Y(n_2847)
);

AOI221xp5_ASAP7_75t_L g2848 ( 
.A1(n_2797),
.A2(n_1240),
.B1(n_1244),
.B2(n_1239),
.C(n_1231),
.Y(n_2848)
);

AOI22xp33_ASAP7_75t_L g2849 ( 
.A1(n_2806),
.A2(n_2764),
.B1(n_2777),
.B2(n_2776),
.Y(n_2849)
);

OR2x2_ASAP7_75t_L g2850 ( 
.A(n_2800),
.B(n_2763),
.Y(n_2850)
);

AND2x4_ASAP7_75t_L g2851 ( 
.A(n_2830),
.B(n_2791),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_2831),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_2810),
.Y(n_2853)
);

OAI21xp5_ASAP7_75t_L g2854 ( 
.A1(n_2809),
.A2(n_2752),
.B(n_2782),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_L g2855 ( 
.A(n_2803),
.B(n_2748),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2832),
.Y(n_2856)
);

BUFx2_ASAP7_75t_L g2857 ( 
.A(n_2794),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2826),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2835),
.Y(n_2859)
);

OR2x2_ASAP7_75t_L g2860 ( 
.A(n_2824),
.B(n_2725),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2821),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2824),
.Y(n_2862)
);

AND2x4_ASAP7_75t_L g2863 ( 
.A(n_2794),
.B(n_2791),
.Y(n_2863)
);

HB1xp67_ASAP7_75t_L g2864 ( 
.A(n_2795),
.Y(n_2864)
);

AND2x2_ASAP7_75t_L g2865 ( 
.A(n_2811),
.B(n_2734),
.Y(n_2865)
);

BUFx2_ASAP7_75t_L g2866 ( 
.A(n_2804),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_L g2867 ( 
.A(n_2812),
.B(n_2742),
.Y(n_2867)
);

AND2x2_ASAP7_75t_L g2868 ( 
.A(n_2827),
.B(n_2790),
.Y(n_2868)
);

BUFx2_ASAP7_75t_L g2869 ( 
.A(n_2804),
.Y(n_2869)
);

AND2x2_ASAP7_75t_L g2870 ( 
.A(n_2804),
.B(n_2771),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2805),
.Y(n_2871)
);

AO22x1_ASAP7_75t_L g2872 ( 
.A1(n_2796),
.A2(n_2788),
.B1(n_2720),
.B2(n_2775),
.Y(n_2872)
);

OAI22xp33_ASAP7_75t_L g2873 ( 
.A1(n_2839),
.A2(n_2798),
.B1(n_2819),
.B2(n_2829),
.Y(n_2873)
);

A2O1A1Ixp33_ASAP7_75t_L g2874 ( 
.A1(n_2865),
.A2(n_2815),
.B(n_2808),
.C(n_2807),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2836),
.Y(n_2875)
);

INVx4_ASAP7_75t_SL g2876 ( 
.A(n_2862),
.Y(n_2876)
);

AND2x4_ASAP7_75t_L g2877 ( 
.A(n_2857),
.B(n_2784),
.Y(n_2877)
);

AND2x4_ASAP7_75t_L g2878 ( 
.A(n_2842),
.B(n_2746),
.Y(n_2878)
);

BUFx4f_ASAP7_75t_L g2879 ( 
.A(n_2839),
.Y(n_2879)
);

AOI22xp5_ASAP7_75t_L g2880 ( 
.A1(n_2864),
.A2(n_2825),
.B1(n_2816),
.B2(n_2801),
.Y(n_2880)
);

AO31x2_ASAP7_75t_L g2881 ( 
.A1(n_2852),
.A2(n_2746),
.A3(n_2751),
.B(n_2747),
.Y(n_2881)
);

AO21x2_ASAP7_75t_L g2882 ( 
.A1(n_2852),
.A2(n_2833),
.B(n_2751),
.Y(n_2882)
);

AOI21xp5_ASAP7_75t_L g2883 ( 
.A1(n_2854),
.A2(n_2814),
.B(n_2817),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2851),
.Y(n_2884)
);

INVx2_ASAP7_75t_L g2885 ( 
.A(n_2851),
.Y(n_2885)
);

AO31x2_ASAP7_75t_L g2886 ( 
.A1(n_2845),
.A2(n_2747),
.A3(n_2737),
.B(n_2758),
.Y(n_2886)
);

BUFx2_ASAP7_75t_L g2887 ( 
.A(n_2863),
.Y(n_2887)
);

INVx2_ASAP7_75t_L g2888 ( 
.A(n_2851),
.Y(n_2888)
);

HB1xp67_ASAP7_75t_L g2889 ( 
.A(n_2853),
.Y(n_2889)
);

A2O1A1Ixp33_ASAP7_75t_L g2890 ( 
.A1(n_2865),
.A2(n_2820),
.B(n_2765),
.C(n_2813),
.Y(n_2890)
);

OAI21x1_ASAP7_75t_L g2891 ( 
.A1(n_2847),
.A2(n_2779),
.B(n_2818),
.Y(n_2891)
);

INVx2_ASAP7_75t_SL g2892 ( 
.A(n_2863),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2838),
.Y(n_2893)
);

BUFx2_ASAP7_75t_L g2894 ( 
.A(n_2863),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2838),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2841),
.Y(n_2896)
);

INVx2_ASAP7_75t_SL g2897 ( 
.A(n_2866),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2844),
.Y(n_2898)
);

OAI22xp5_ASAP7_75t_L g2899 ( 
.A1(n_2864),
.A2(n_2822),
.B1(n_2774),
.B2(n_1248),
.Y(n_2899)
);

INVx2_ASAP7_75t_L g2900 ( 
.A(n_2860),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2846),
.Y(n_2901)
);

AOI21xp5_ASAP7_75t_L g2902 ( 
.A1(n_2867),
.A2(n_1249),
.B(n_1247),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_L g2903 ( 
.A(n_2859),
.B(n_2774),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2850),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2840),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2843),
.Y(n_2906)
);

OR2x2_ASAP7_75t_L g2907 ( 
.A(n_2837),
.B(n_2754),
.Y(n_2907)
);

AO21x2_ASAP7_75t_L g2908 ( 
.A1(n_2847),
.A2(n_2754),
.B(n_2774),
.Y(n_2908)
);

OAI21x1_ASAP7_75t_L g2909 ( 
.A1(n_2853),
.A2(n_2754),
.B(n_13),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2840),
.Y(n_2910)
);

INVx2_ASAP7_75t_L g2911 ( 
.A(n_2869),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2875),
.Y(n_2912)
);

AND2x2_ASAP7_75t_L g2913 ( 
.A(n_2887),
.B(n_2842),
.Y(n_2913)
);

AND2x2_ASAP7_75t_L g2914 ( 
.A(n_2876),
.B(n_2842),
.Y(n_2914)
);

INVx2_ASAP7_75t_L g2915 ( 
.A(n_2881),
.Y(n_2915)
);

NOR2xp67_ASAP7_75t_SL g2916 ( 
.A(n_2883),
.B(n_2871),
.Y(n_2916)
);

HB1xp67_ASAP7_75t_L g2917 ( 
.A(n_2894),
.Y(n_2917)
);

AND2x2_ASAP7_75t_L g2918 ( 
.A(n_2892),
.B(n_2856),
.Y(n_2918)
);

BUFx2_ASAP7_75t_L g2919 ( 
.A(n_2879),
.Y(n_2919)
);

AND2x2_ASAP7_75t_L g2920 ( 
.A(n_2884),
.B(n_2870),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2875),
.Y(n_2921)
);

OR2x2_ASAP7_75t_L g2922 ( 
.A(n_2904),
.B(n_2861),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2898),
.Y(n_2923)
);

AND2x4_ASAP7_75t_L g2924 ( 
.A(n_2876),
.B(n_2858),
.Y(n_2924)
);

AND2x2_ASAP7_75t_L g2925 ( 
.A(n_2885),
.B(n_2870),
.Y(n_2925)
);

AND2x2_ASAP7_75t_L g2926 ( 
.A(n_2888),
.B(n_2872),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2902),
.B(n_2868),
.Y(n_2927)
);

INVx1_ASAP7_75t_SL g2928 ( 
.A(n_2897),
.Y(n_2928)
);

AND2x4_ASAP7_75t_L g2929 ( 
.A(n_2901),
.B(n_2868),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_L g2930 ( 
.A(n_2911),
.B(n_2855),
.Y(n_2930)
);

AND2x4_ASAP7_75t_L g2931 ( 
.A(n_2900),
.B(n_2849),
.Y(n_2931)
);

AOI211xp5_ASAP7_75t_L g2932 ( 
.A1(n_2873),
.A2(n_2848),
.B(n_1251),
.C(n_1252),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_2881),
.Y(n_2933)
);

INVx2_ASAP7_75t_L g2934 ( 
.A(n_2881),
.Y(n_2934)
);

BUFx6f_ASAP7_75t_L g2935 ( 
.A(n_2879),
.Y(n_2935)
);

AND2x2_ASAP7_75t_L g2936 ( 
.A(n_2906),
.B(n_2849),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2905),
.Y(n_2937)
);

AND2x2_ASAP7_75t_L g2938 ( 
.A(n_2878),
.B(n_14),
.Y(n_2938)
);

AOI22xp33_ASAP7_75t_SL g2939 ( 
.A1(n_2899),
.A2(n_1253),
.B1(n_1255),
.B2(n_1250),
.Y(n_2939)
);

AND2x2_ASAP7_75t_L g2940 ( 
.A(n_2878),
.B(n_14),
.Y(n_2940)
);

AND2x2_ASAP7_75t_L g2941 ( 
.A(n_2877),
.B(n_15),
.Y(n_2941)
);

AND2x2_ASAP7_75t_L g2942 ( 
.A(n_2877),
.B(n_2896),
.Y(n_2942)
);

AOI22xp33_ASAP7_75t_SL g2943 ( 
.A1(n_2882),
.A2(n_2891),
.B1(n_2903),
.B2(n_2889),
.Y(n_2943)
);

INVx3_ASAP7_75t_L g2944 ( 
.A(n_2886),
.Y(n_2944)
);

OAI221xp5_ASAP7_75t_L g2945 ( 
.A1(n_2890),
.A2(n_1274),
.B1(n_1276),
.B2(n_1268),
.C(n_1264),
.Y(n_2945)
);

OAI31xp33_ASAP7_75t_L g2946 ( 
.A1(n_2874),
.A2(n_18),
.A3(n_16),
.B(n_17),
.Y(n_2946)
);

INVx4_ASAP7_75t_L g2947 ( 
.A(n_2882),
.Y(n_2947)
);

HB1xp67_ASAP7_75t_L g2948 ( 
.A(n_2917),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2944),
.Y(n_2949)
);

AND2x2_ASAP7_75t_L g2950 ( 
.A(n_2914),
.B(n_2896),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2912),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2921),
.Y(n_2952)
);

AND2x2_ASAP7_75t_L g2953 ( 
.A(n_2913),
.B(n_2905),
.Y(n_2953)
);

AND2x2_ASAP7_75t_L g2954 ( 
.A(n_2913),
.B(n_2910),
.Y(n_2954)
);

AND2x2_ASAP7_75t_L g2955 ( 
.A(n_2926),
.B(n_2910),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2931),
.B(n_2880),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_SL g2957 ( 
.A(n_2946),
.B(n_2907),
.Y(n_2957)
);

NAND2x1p5_ASAP7_75t_L g2958 ( 
.A(n_2924),
.B(n_2909),
.Y(n_2958)
);

NAND2x1p5_ASAP7_75t_L g2959 ( 
.A(n_2924),
.B(n_2893),
.Y(n_2959)
);

INVx2_ASAP7_75t_L g2960 ( 
.A(n_2944),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2937),
.Y(n_2961)
);

INVx3_ASAP7_75t_L g2962 ( 
.A(n_2924),
.Y(n_2962)
);

AND2x2_ASAP7_75t_L g2963 ( 
.A(n_2926),
.B(n_2895),
.Y(n_2963)
);

AND2x2_ASAP7_75t_L g2964 ( 
.A(n_2928),
.B(n_2895),
.Y(n_2964)
);

INVx2_ASAP7_75t_L g2965 ( 
.A(n_2944),
.Y(n_2965)
);

NAND2x1_ASAP7_75t_L g2966 ( 
.A(n_2947),
.B(n_2886),
.Y(n_2966)
);

INVx2_ASAP7_75t_L g2967 ( 
.A(n_2947),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2922),
.Y(n_2968)
);

INVx1_ASAP7_75t_SL g2969 ( 
.A(n_2919),
.Y(n_2969)
);

NOR2xp67_ASAP7_75t_L g2970 ( 
.A(n_2935),
.B(n_2947),
.Y(n_2970)
);

INVx3_ASAP7_75t_L g2971 ( 
.A(n_2935),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2931),
.B(n_2886),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2923),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2931),
.B(n_2908),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2915),
.Y(n_2975)
);

AND2x2_ASAP7_75t_L g2976 ( 
.A(n_2920),
.B(n_2908),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_L g2977 ( 
.A(n_2936),
.B(n_17),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_L g2978 ( 
.A(n_2941),
.B(n_19),
.Y(n_2978)
);

NAND2xp33_ASAP7_75t_SL g2979 ( 
.A(n_2916),
.B(n_22),
.Y(n_2979)
);

AND2x2_ASAP7_75t_L g2980 ( 
.A(n_2920),
.B(n_22),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2941),
.B(n_23),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2915),
.Y(n_2982)
);

AND2x2_ASAP7_75t_L g2983 ( 
.A(n_2925),
.B(n_23),
.Y(n_2983)
);

INVx2_ASAP7_75t_L g2984 ( 
.A(n_2933),
.Y(n_2984)
);

AND2x2_ASAP7_75t_L g2985 ( 
.A(n_2925),
.B(n_24),
.Y(n_2985)
);

AND2x2_ASAP7_75t_L g2986 ( 
.A(n_2942),
.B(n_24),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2938),
.Y(n_2987)
);

NOR2x1p5_ASAP7_75t_L g2988 ( 
.A(n_2935),
.B(n_25),
.Y(n_2988)
);

AND2x2_ASAP7_75t_L g2989 ( 
.A(n_2942),
.B(n_25),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2938),
.Y(n_2990)
);

AND2x2_ASAP7_75t_L g2991 ( 
.A(n_2929),
.B(n_26),
.Y(n_2991)
);

AND2x2_ASAP7_75t_L g2992 ( 
.A(n_2929),
.B(n_27),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_2933),
.Y(n_2993)
);

AND2x2_ASAP7_75t_L g2994 ( 
.A(n_2929),
.B(n_28),
.Y(n_2994)
);

NOR3xp33_ASAP7_75t_SL g2995 ( 
.A(n_2956),
.B(n_2945),
.C(n_2927),
.Y(n_2995)
);

NAND2xp5_ASAP7_75t_L g2996 ( 
.A(n_2969),
.B(n_2940),
.Y(n_2996)
);

HB1xp67_ASAP7_75t_L g2997 ( 
.A(n_2948),
.Y(n_2997)
);

NAND4xp75_ASAP7_75t_SL g2998 ( 
.A(n_2970),
.B(n_2918),
.C(n_2940),
.D(n_2943),
.Y(n_2998)
);

NAND4xp75_ASAP7_75t_SL g2999 ( 
.A(n_2950),
.B(n_2918),
.C(n_2935),
.D(n_2932),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2975),
.Y(n_3000)
);

NAND2xp5_ASAP7_75t_L g3001 ( 
.A(n_2986),
.B(n_2930),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2975),
.Y(n_3002)
);

NAND4xp25_ASAP7_75t_L g3003 ( 
.A(n_2971),
.B(n_2939),
.C(n_2934),
.D(n_31),
.Y(n_3003)
);

XOR2x2_ASAP7_75t_L g3004 ( 
.A(n_2957),
.B(n_29),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_2986),
.B(n_2934),
.Y(n_3005)
);

NAND4xp75_ASAP7_75t_L g3006 ( 
.A(n_2957),
.B(n_2974),
.C(n_2972),
.D(n_2976),
.Y(n_3006)
);

NOR2x1_ASAP7_75t_L g3007 ( 
.A(n_2962),
.B(n_29),
.Y(n_3007)
);

OR2x2_ASAP7_75t_L g3008 ( 
.A(n_2987),
.B(n_30),
.Y(n_3008)
);

AND2x2_ASAP7_75t_L g3009 ( 
.A(n_2950),
.B(n_30),
.Y(n_3009)
);

AND2x2_ASAP7_75t_L g3010 ( 
.A(n_2990),
.B(n_32),
.Y(n_3010)
);

BUFx2_ASAP7_75t_L g3011 ( 
.A(n_2962),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2982),
.Y(n_3012)
);

INVx2_ASAP7_75t_L g3013 ( 
.A(n_2962),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2982),
.Y(n_3014)
);

INVx6_ASAP7_75t_L g3015 ( 
.A(n_2988),
.Y(n_3015)
);

OR2x2_ASAP7_75t_L g3016 ( 
.A(n_2977),
.B(n_2968),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2984),
.Y(n_3017)
);

NAND4xp75_ASAP7_75t_L g3018 ( 
.A(n_2976),
.B(n_35),
.C(n_33),
.D(n_34),
.Y(n_3018)
);

AND2x2_ASAP7_75t_L g3019 ( 
.A(n_2971),
.B(n_33),
.Y(n_3019)
);

BUFx3_ASAP7_75t_L g3020 ( 
.A(n_2971),
.Y(n_3020)
);

NOR2x1_ASAP7_75t_L g3021 ( 
.A(n_2989),
.B(n_35),
.Y(n_3021)
);

AND2x4_ASAP7_75t_L g3022 ( 
.A(n_2964),
.B(n_36),
.Y(n_3022)
);

NOR2xp33_ASAP7_75t_L g3023 ( 
.A(n_2978),
.B(n_36),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_L g3024 ( 
.A(n_2989),
.B(n_37),
.Y(n_3024)
);

INVx2_ASAP7_75t_L g3025 ( 
.A(n_2959),
.Y(n_3025)
);

AND2x2_ASAP7_75t_SL g3026 ( 
.A(n_2983),
.B(n_38),
.Y(n_3026)
);

BUFx3_ASAP7_75t_L g3027 ( 
.A(n_2992),
.Y(n_3027)
);

INVx2_ASAP7_75t_L g3028 ( 
.A(n_2959),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2984),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2983),
.B(n_38),
.Y(n_3030)
);

AND2x2_ASAP7_75t_L g3031 ( 
.A(n_2985),
.B(n_39),
.Y(n_3031)
);

AND2x4_ASAP7_75t_L g3032 ( 
.A(n_2964),
.B(n_39),
.Y(n_3032)
);

INVx2_ASAP7_75t_SL g3033 ( 
.A(n_2954),
.Y(n_3033)
);

AND2x2_ASAP7_75t_L g3034 ( 
.A(n_2985),
.B(n_40),
.Y(n_3034)
);

INVx2_ASAP7_75t_L g3035 ( 
.A(n_2955),
.Y(n_3035)
);

AND2x2_ASAP7_75t_L g3036 ( 
.A(n_2955),
.B(n_40),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2993),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_L g3038 ( 
.A(n_2991),
.B(n_42),
.Y(n_3038)
);

NAND4xp75_ASAP7_75t_SL g3039 ( 
.A(n_2963),
.B(n_44),
.C(n_42),
.D(n_43),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2993),
.Y(n_3040)
);

XNOR2xp5_ASAP7_75t_L g3041 ( 
.A(n_2979),
.B(n_43),
.Y(n_3041)
);

INVxp67_ASAP7_75t_SL g3042 ( 
.A(n_2958),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_2963),
.Y(n_3043)
);

OR2x2_ASAP7_75t_L g3044 ( 
.A(n_2953),
.B(n_44),
.Y(n_3044)
);

OAI22xp33_ASAP7_75t_L g3045 ( 
.A1(n_2958),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_3045)
);

AND2x2_ASAP7_75t_L g3046 ( 
.A(n_2954),
.B(n_47),
.Y(n_3046)
);

XOR2x2_ASAP7_75t_L g3047 ( 
.A(n_2981),
.B(n_48),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_L g3048 ( 
.A(n_2991),
.B(n_2994),
.Y(n_3048)
);

NAND4xp75_ASAP7_75t_L g3049 ( 
.A(n_2994),
.B(n_2967),
.C(n_2973),
.D(n_2951),
.Y(n_3049)
);

NOR3xp33_ASAP7_75t_L g3050 ( 
.A(n_2979),
.B(n_49),
.C(n_50),
.Y(n_3050)
);

INVxp67_ASAP7_75t_SL g3051 ( 
.A(n_2966),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2967),
.Y(n_3052)
);

INVx2_ASAP7_75t_L g3053 ( 
.A(n_2949),
.Y(n_3053)
);

OR2x2_ASAP7_75t_L g3054 ( 
.A(n_2980),
.B(n_50),
.Y(n_3054)
);

AND2x2_ASAP7_75t_L g3055 ( 
.A(n_2952),
.B(n_2961),
.Y(n_3055)
);

INVx2_ASAP7_75t_L g3056 ( 
.A(n_2949),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2960),
.Y(n_3057)
);

INVx2_ASAP7_75t_L g3058 ( 
.A(n_2960),
.Y(n_3058)
);

INVx8_ASAP7_75t_L g3059 ( 
.A(n_2965),
.Y(n_3059)
);

NAND4xp75_ASAP7_75t_L g3060 ( 
.A(n_2965),
.B(n_54),
.C(n_52),
.D(n_53),
.Y(n_3060)
);

AND2x2_ASAP7_75t_L g3061 ( 
.A(n_2969),
.B(n_52),
.Y(n_3061)
);

AOI22xp5_ASAP7_75t_L g3062 ( 
.A1(n_2957),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_L g3063 ( 
.A(n_3026),
.B(n_55),
.Y(n_3063)
);

NAND3x2_ASAP7_75t_L g3064 ( 
.A(n_2998),
.B(n_56),
.C(n_57),
.Y(n_3064)
);

HB1xp67_ASAP7_75t_L g3065 ( 
.A(n_3011),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2997),
.Y(n_3066)
);

INVx2_ASAP7_75t_SL g3067 ( 
.A(n_3059),
.Y(n_3067)
);

AND2x2_ASAP7_75t_L g3068 ( 
.A(n_3015),
.B(n_57),
.Y(n_3068)
);

INVx1_ASAP7_75t_SL g3069 ( 
.A(n_3015),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_L g3070 ( 
.A(n_3007),
.B(n_58),
.Y(n_3070)
);

NOR2xp33_ASAP7_75t_L g3071 ( 
.A(n_3027),
.B(n_59),
.Y(n_3071)
);

AND2x4_ASAP7_75t_L g3072 ( 
.A(n_3013),
.B(n_60),
.Y(n_3072)
);

AND2x2_ASAP7_75t_L g3073 ( 
.A(n_3021),
.B(n_3033),
.Y(n_3073)
);

AOI21xp33_ASAP7_75t_L g3074 ( 
.A1(n_3042),
.A2(n_59),
.B(n_61),
.Y(n_3074)
);

INVx2_ASAP7_75t_L g3075 ( 
.A(n_3020),
.Y(n_3075)
);

OR2x2_ASAP7_75t_L g3076 ( 
.A(n_2996),
.B(n_62),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_3035),
.Y(n_3077)
);

AND2x2_ASAP7_75t_L g3078 ( 
.A(n_3061),
.B(n_62),
.Y(n_3078)
);

INVxp67_ASAP7_75t_L g3079 ( 
.A(n_3018),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_3043),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_3057),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_3057),
.Y(n_3082)
);

AND2x2_ASAP7_75t_L g3083 ( 
.A(n_3009),
.B(n_63),
.Y(n_3083)
);

AND2x2_ASAP7_75t_L g3084 ( 
.A(n_3036),
.B(n_63),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_3029),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_3022),
.B(n_64),
.Y(n_3086)
);

AOI21xp5_ASAP7_75t_L g3087 ( 
.A1(n_3004),
.A2(n_64),
.B(n_65),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_3029),
.Y(n_3088)
);

INVxp67_ASAP7_75t_L g3089 ( 
.A(n_3049),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_3037),
.Y(n_3090)
);

INVx2_ASAP7_75t_L g3091 ( 
.A(n_3025),
.Y(n_3091)
);

INVx2_ASAP7_75t_L g3092 ( 
.A(n_3028),
.Y(n_3092)
);

AND2x2_ASAP7_75t_L g3093 ( 
.A(n_3046),
.B(n_65),
.Y(n_3093)
);

OR2x2_ASAP7_75t_L g3094 ( 
.A(n_3048),
.B(n_3001),
.Y(n_3094)
);

INVxp67_ASAP7_75t_L g3095 ( 
.A(n_3060),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_3037),
.Y(n_3096)
);

NAND2xp5_ASAP7_75t_L g3097 ( 
.A(n_3022),
.B(n_3032),
.Y(n_3097)
);

INVx1_ASAP7_75t_SL g3098 ( 
.A(n_3031),
.Y(n_3098)
);

OR2x2_ASAP7_75t_L g3099 ( 
.A(n_3016),
.B(n_66),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_3040),
.Y(n_3100)
);

AND2x4_ASAP7_75t_L g3101 ( 
.A(n_3032),
.B(n_68),
.Y(n_3101)
);

OR2x2_ASAP7_75t_L g3102 ( 
.A(n_3044),
.B(n_67),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_3040),
.Y(n_3103)
);

INVx1_ASAP7_75t_SL g3104 ( 
.A(n_3034),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_3000),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_3002),
.Y(n_3106)
);

OR2x2_ASAP7_75t_L g3107 ( 
.A(n_3005),
.B(n_67),
.Y(n_3107)
);

OR2x2_ASAP7_75t_L g3108 ( 
.A(n_3003),
.B(n_68),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_3012),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_3014),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_SL g3111 ( 
.A(n_3045),
.B(n_69),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_3050),
.B(n_69),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_3017),
.Y(n_3113)
);

AND2x2_ASAP7_75t_L g3114 ( 
.A(n_3019),
.B(n_70),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_3052),
.Y(n_3115)
);

NOR2xp67_ASAP7_75t_SL g3116 ( 
.A(n_3054),
.B(n_70),
.Y(n_3116)
);

BUFx2_ASAP7_75t_L g3117 ( 
.A(n_3059),
.Y(n_3117)
);

NAND2xp67_ASAP7_75t_L g3118 ( 
.A(n_3010),
.B(n_3055),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_L g3119 ( 
.A(n_3006),
.B(n_71),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_L g3120 ( 
.A(n_3062),
.B(n_71),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_3052),
.Y(n_3121)
);

NAND2x1_ASAP7_75t_SL g3122 ( 
.A(n_3053),
.B(n_72),
.Y(n_3122)
);

AOI22xp5_ASAP7_75t_L g3123 ( 
.A1(n_2995),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_3056),
.Y(n_3124)
);

HB1xp67_ASAP7_75t_L g3125 ( 
.A(n_3058),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_3008),
.Y(n_3126)
);

AND2x2_ASAP7_75t_L g3127 ( 
.A(n_3023),
.B(n_75),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_L g3128 ( 
.A(n_3047),
.B(n_75),
.Y(n_3128)
);

OR2x2_ASAP7_75t_L g3129 ( 
.A(n_3024),
.B(n_77),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_3038),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_3030),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_L g3132 ( 
.A(n_3041),
.B(n_77),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_3051),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_3039),
.Y(n_3134)
);

INVx2_ASAP7_75t_L g3135 ( 
.A(n_2999),
.Y(n_3135)
);

INVxp33_ASAP7_75t_L g3136 ( 
.A(n_3021),
.Y(n_3136)
);

INVx3_ASAP7_75t_L g3137 ( 
.A(n_3020),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2997),
.Y(n_3138)
);

OR2x2_ASAP7_75t_L g3139 ( 
.A(n_2996),
.B(n_78),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2997),
.Y(n_3140)
);

INVx1_ASAP7_75t_SL g3141 ( 
.A(n_3015),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_2997),
.Y(n_3142)
);

INVxp67_ASAP7_75t_L g3143 ( 
.A(n_3007),
.Y(n_3143)
);

OR2x2_ASAP7_75t_L g3144 ( 
.A(n_2996),
.B(n_79),
.Y(n_3144)
);

AND2x2_ASAP7_75t_L g3145 ( 
.A(n_3015),
.B(n_80),
.Y(n_3145)
);

INVx1_ASAP7_75t_L g3146 ( 
.A(n_2997),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_L g3147 ( 
.A(n_3026),
.B(n_80),
.Y(n_3147)
);

NAND2x1p5_ASAP7_75t_L g3148 ( 
.A(n_3021),
.B(n_81),
.Y(n_3148)
);

AND2x2_ASAP7_75t_L g3149 ( 
.A(n_3015),
.B(n_82),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2997),
.Y(n_3150)
);

NOR2x1_ASAP7_75t_L g3151 ( 
.A(n_3007),
.B(n_82),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_2997),
.Y(n_3152)
);

NAND3xp33_ASAP7_75t_L g3153 ( 
.A(n_2995),
.B(n_84),
.C(n_85),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_2997),
.Y(n_3154)
);

INVx2_ASAP7_75t_L g3155 ( 
.A(n_3011),
.Y(n_3155)
);

NAND2x1_ASAP7_75t_L g3156 ( 
.A(n_3011),
.B(n_86),
.Y(n_3156)
);

AOI22xp33_ASAP7_75t_L g3157 ( 
.A1(n_3064),
.A2(n_1518),
.B1(n_1504),
.B2(n_88),
.Y(n_3157)
);

INVx2_ASAP7_75t_L g3158 ( 
.A(n_3148),
.Y(n_3158)
);

AND2x2_ASAP7_75t_L g3159 ( 
.A(n_3069),
.B(n_86),
.Y(n_3159)
);

AOI22xp5_ASAP7_75t_L g3160 ( 
.A1(n_3089),
.A2(n_3153),
.B1(n_3123),
.B2(n_3079),
.Y(n_3160)
);

OAI21xp33_ASAP7_75t_SL g3161 ( 
.A1(n_3119),
.A2(n_87),
.B(n_88),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_3065),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_3125),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_3154),
.Y(n_3164)
);

O2A1O1Ixp33_ASAP7_75t_SL g3165 ( 
.A1(n_3143),
.A2(n_91),
.B(n_89),
.C(n_90),
.Y(n_3165)
);

AOI211xp5_ASAP7_75t_SL g3166 ( 
.A1(n_3066),
.A2(n_92),
.B(n_89),
.C(n_91),
.Y(n_3166)
);

AO21x1_ASAP7_75t_L g3167 ( 
.A1(n_3156),
.A2(n_97),
.B(n_96),
.Y(n_3167)
);

OAI22xp5_ASAP7_75t_L g3168 ( 
.A1(n_3136),
.A2(n_100),
.B1(n_94),
.B2(n_99),
.Y(n_3168)
);

XOR2x2_ASAP7_75t_L g3169 ( 
.A(n_3151),
.B(n_102),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_3154),
.Y(n_3170)
);

AOI22xp33_ASAP7_75t_L g3171 ( 
.A1(n_3135),
.A2(n_1518),
.B1(n_1504),
.B2(n_104),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_3117),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_3073),
.Y(n_3173)
);

INVx4_ASAP7_75t_L g3174 ( 
.A(n_3101),
.Y(n_3174)
);

INVx2_ASAP7_75t_L g3175 ( 
.A(n_3137),
.Y(n_3175)
);

AOI22xp5_ASAP7_75t_L g3176 ( 
.A1(n_3095),
.A2(n_105),
.B1(n_102),
.B2(n_103),
.Y(n_3176)
);

INVxp67_ASAP7_75t_L g3177 ( 
.A(n_3116),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_3141),
.B(n_103),
.Y(n_3178)
);

AOI21xp33_ASAP7_75t_L g3179 ( 
.A1(n_3067),
.A2(n_106),
.B(n_107),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_3084),
.Y(n_3180)
);

XNOR2xp5_ASAP7_75t_L g3181 ( 
.A(n_3098),
.B(n_106),
.Y(n_3181)
);

XNOR2xp5_ASAP7_75t_L g3182 ( 
.A(n_3104),
.B(n_108),
.Y(n_3182)
);

XOR2x2_ASAP7_75t_L g3183 ( 
.A(n_3122),
.B(n_109),
.Y(n_3183)
);

OAI21xp5_ASAP7_75t_L g3184 ( 
.A1(n_3087),
.A2(n_109),
.B(n_113),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_3093),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_3083),
.Y(n_3186)
);

INVx3_ASAP7_75t_L g3187 ( 
.A(n_3137),
.Y(n_3187)
);

OAI21xp33_ASAP7_75t_L g3188 ( 
.A1(n_3118),
.A2(n_114),
.B(n_115),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_3138),
.Y(n_3189)
);

INVxp67_ASAP7_75t_L g3190 ( 
.A(n_3097),
.Y(n_3190)
);

AOI22xp5_ASAP7_75t_L g3191 ( 
.A1(n_3075),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_3191)
);

INVx2_ASAP7_75t_L g3192 ( 
.A(n_3155),
.Y(n_3192)
);

AOI21xp5_ASAP7_75t_L g3193 ( 
.A1(n_3111),
.A2(n_116),
.B(n_117),
.Y(n_3193)
);

AOI211xp5_ASAP7_75t_SL g3194 ( 
.A1(n_3140),
.A2(n_119),
.B(n_117),
.C(n_118),
.Y(n_3194)
);

NAND2x1p5_ASAP7_75t_L g3195 ( 
.A(n_3101),
.B(n_119),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_3142),
.Y(n_3196)
);

OAI21xp5_ASAP7_75t_SL g3197 ( 
.A1(n_3108),
.A2(n_120),
.B(n_121),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_3146),
.Y(n_3198)
);

OAI22xp33_ASAP7_75t_SL g3199 ( 
.A1(n_3150),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.Y(n_3199)
);

AOI21xp33_ASAP7_75t_L g3200 ( 
.A1(n_3094),
.A2(n_123),
.B(n_124),
.Y(n_3200)
);

NAND2xp33_ASAP7_75t_L g3201 ( 
.A(n_3134),
.B(n_125),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_3152),
.Y(n_3202)
);

NAND3xp33_ASAP7_75t_L g3203 ( 
.A(n_3091),
.B(n_125),
.C(n_126),
.Y(n_3203)
);

OAI22xp33_ASAP7_75t_L g3204 ( 
.A1(n_3112),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_3204)
);

OAI211xp5_ASAP7_75t_L g3205 ( 
.A1(n_3074),
.A2(n_130),
.B(n_128),
.C(n_129),
.Y(n_3205)
);

AOI22xp33_ASAP7_75t_L g3206 ( 
.A1(n_3131),
.A2(n_1518),
.B1(n_1504),
.B2(n_133),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_SL g3207 ( 
.A(n_3126),
.B(n_131),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_3115),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_3121),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_3081),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_3082),
.Y(n_3211)
);

OAI22xp5_ASAP7_75t_L g3212 ( 
.A1(n_3128),
.A2(n_134),
.B1(n_131),
.B2(n_132),
.Y(n_3212)
);

INVx2_ASAP7_75t_L g3213 ( 
.A(n_3068),
.Y(n_3213)
);

AOI21xp33_ASAP7_75t_L g3214 ( 
.A1(n_3130),
.A2(n_132),
.B(n_134),
.Y(n_3214)
);

AOI211xp5_ASAP7_75t_L g3215 ( 
.A1(n_3092),
.A2(n_137),
.B(n_135),
.C(n_136),
.Y(n_3215)
);

INVxp67_ASAP7_75t_L g3216 ( 
.A(n_3070),
.Y(n_3216)
);

AOI21xp5_ASAP7_75t_L g3217 ( 
.A1(n_3063),
.A2(n_137),
.B(n_138),
.Y(n_3217)
);

INVx1_ASAP7_75t_L g3218 ( 
.A(n_3086),
.Y(n_3218)
);

OAI21xp5_ASAP7_75t_L g3219 ( 
.A1(n_3120),
.A2(n_138),
.B(n_139),
.Y(n_3219)
);

OAI22xp5_ASAP7_75t_L g3220 ( 
.A1(n_3133),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.Y(n_3220)
);

AOI22xp33_ASAP7_75t_SL g3221 ( 
.A1(n_3077),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_3221)
);

INVx1_ASAP7_75t_L g3222 ( 
.A(n_3078),
.Y(n_3222)
);

OAI21xp5_ASAP7_75t_L g3223 ( 
.A1(n_3080),
.A2(n_142),
.B(n_144),
.Y(n_3223)
);

NOR2xp33_ASAP7_75t_L g3224 ( 
.A(n_3076),
.B(n_145),
.Y(n_3224)
);

NAND4xp25_ASAP7_75t_L g3225 ( 
.A(n_3124),
.B(n_147),
.C(n_145),
.D(n_146),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_3114),
.Y(n_3226)
);

O2A1O1Ixp33_ASAP7_75t_SL g3227 ( 
.A1(n_3147),
.A2(n_3132),
.B(n_3099),
.C(n_3110),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_3102),
.Y(n_3228)
);

INVx1_ASAP7_75t_SL g3229 ( 
.A(n_3145),
.Y(n_3229)
);

OAI21xp33_ASAP7_75t_SL g3230 ( 
.A1(n_3110),
.A2(n_146),
.B(n_148),
.Y(n_3230)
);

O2A1O1Ixp5_ASAP7_75t_L g3231 ( 
.A1(n_3105),
.A2(n_152),
.B(n_149),
.C(n_150),
.Y(n_3231)
);

AOI21xp33_ASAP7_75t_L g3232 ( 
.A1(n_3139),
.A2(n_152),
.B(n_153),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_3149),
.B(n_154),
.Y(n_3233)
);

OAI22xp5_ASAP7_75t_L g3234 ( 
.A1(n_3144),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_3234)
);

NAND2xp5_ASAP7_75t_L g3235 ( 
.A(n_3071),
.B(n_155),
.Y(n_3235)
);

XNOR2xp5_ASAP7_75t_L g3236 ( 
.A(n_3127),
.B(n_157),
.Y(n_3236)
);

INVx2_ASAP7_75t_L g3237 ( 
.A(n_3072),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_3085),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_L g3239 ( 
.A(n_3072),
.B(n_157),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_L g3240 ( 
.A(n_3129),
.B(n_3107),
.Y(n_3240)
);

INVx2_ASAP7_75t_L g3241 ( 
.A(n_3088),
.Y(n_3241)
);

OAI21xp33_ASAP7_75t_SL g3242 ( 
.A1(n_3090),
.A2(n_158),
.B(n_159),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_3096),
.Y(n_3243)
);

INVx2_ASAP7_75t_L g3244 ( 
.A(n_3100),
.Y(n_3244)
);

AOI22xp5_ASAP7_75t_L g3245 ( 
.A1(n_3106),
.A2(n_162),
.B1(n_160),
.B2(n_161),
.Y(n_3245)
);

NAND3xp33_ASAP7_75t_L g3246 ( 
.A(n_3109),
.B(n_3113),
.C(n_3103),
.Y(n_3246)
);

AOI22xp5_ASAP7_75t_L g3247 ( 
.A1(n_3064),
.A2(n_165),
.B1(n_163),
.B2(n_164),
.Y(n_3247)
);

AOI211xp5_ASAP7_75t_L g3248 ( 
.A1(n_3136),
.A2(n_166),
.B(n_164),
.C(n_165),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_3065),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_3065),
.Y(n_3250)
);

OAI21xp33_ASAP7_75t_L g3251 ( 
.A1(n_3089),
.A2(n_166),
.B(n_167),
.Y(n_3251)
);

INVx1_ASAP7_75t_L g3252 ( 
.A(n_3065),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_3065),
.Y(n_3253)
);

INVxp67_ASAP7_75t_L g3254 ( 
.A(n_3151),
.Y(n_3254)
);

AOI22xp5_ASAP7_75t_L g3255 ( 
.A1(n_3064),
.A2(n_171),
.B1(n_167),
.B2(n_169),
.Y(n_3255)
);

OAI22x1_ASAP7_75t_L g3256 ( 
.A1(n_3123),
.A2(n_173),
.B1(n_169),
.B2(n_172),
.Y(n_3256)
);

NAND2xp5_ASAP7_75t_L g3257 ( 
.A(n_3069),
.B(n_172),
.Y(n_3257)
);

NAND2x1p5_ASAP7_75t_L g3258 ( 
.A(n_3151),
.B(n_173),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_3065),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_3065),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_L g3261 ( 
.A(n_3069),
.B(n_174),
.Y(n_3261)
);

OAI22xp5_ASAP7_75t_L g3262 ( 
.A1(n_3064),
.A2(n_176),
.B1(n_174),
.B2(n_175),
.Y(n_3262)
);

OAI31xp33_ASAP7_75t_L g3263 ( 
.A1(n_3153),
.A2(n_177),
.A3(n_175),
.B(n_176),
.Y(n_3263)
);

AOI22xp5_ASAP7_75t_L g3264 ( 
.A1(n_3064),
.A2(n_181),
.B1(n_178),
.B2(n_179),
.Y(n_3264)
);

XNOR2xp5_ASAP7_75t_L g3265 ( 
.A(n_3064),
.B(n_178),
.Y(n_3265)
);

AOI22xp5_ASAP7_75t_L g3266 ( 
.A1(n_3064),
.A2(n_185),
.B1(n_181),
.B2(n_184),
.Y(n_3266)
);

AOI22xp33_ASAP7_75t_L g3267 ( 
.A1(n_3064),
.A2(n_1518),
.B1(n_187),
.B2(n_184),
.Y(n_3267)
);

NOR2x1_ASAP7_75t_L g3268 ( 
.A(n_3119),
.B(n_186),
.Y(n_3268)
);

INVx2_ASAP7_75t_SL g3269 ( 
.A(n_3122),
.Y(n_3269)
);

AOI21xp33_ASAP7_75t_SL g3270 ( 
.A1(n_3143),
.A2(n_186),
.B(n_188),
.Y(n_3270)
);

O2A1O1Ixp33_ASAP7_75t_L g3271 ( 
.A1(n_3143),
.A2(n_190),
.B(n_188),
.C(n_189),
.Y(n_3271)
);

OAI22xp5_ASAP7_75t_L g3272 ( 
.A1(n_3064),
.A2(n_193),
.B1(n_191),
.B2(n_192),
.Y(n_3272)
);

OAI22xp33_ASAP7_75t_L g3273 ( 
.A1(n_3123),
.A2(n_196),
.B1(n_194),
.B2(n_195),
.Y(n_3273)
);

AOI21xp33_ASAP7_75t_L g3274 ( 
.A1(n_3136),
.A2(n_195),
.B(n_197),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_3065),
.Y(n_3275)
);

AOI22xp5_ASAP7_75t_L g3276 ( 
.A1(n_3064),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.Y(n_3276)
);

AOI22xp33_ASAP7_75t_L g3277 ( 
.A1(n_3064),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_3277)
);

OAI21xp5_ASAP7_75t_L g3278 ( 
.A1(n_3064),
.A2(n_201),
.B(n_202),
.Y(n_3278)
);

OAI22xp33_ASAP7_75t_SL g3279 ( 
.A1(n_3143),
.A2(n_204),
.B1(n_202),
.B2(n_203),
.Y(n_3279)
);

AOI211xp5_ASAP7_75t_SL g3280 ( 
.A1(n_3089),
.A2(n_206),
.B(n_204),
.C(n_205),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_3065),
.Y(n_3281)
);

INVx1_ASAP7_75t_SL g3282 ( 
.A(n_3122),
.Y(n_3282)
);

OAI31xp33_ASAP7_75t_L g3283 ( 
.A1(n_3153),
.A2(n_210),
.A3(n_207),
.B(n_208),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_3065),
.Y(n_3284)
);

AOI22xp33_ASAP7_75t_SL g3285 ( 
.A1(n_3064),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.Y(n_3285)
);

INVxp67_ASAP7_75t_SL g3286 ( 
.A(n_3122),
.Y(n_3286)
);

OAI22xp33_ASAP7_75t_L g3287 ( 
.A1(n_3123),
.A2(n_213),
.B1(n_211),
.B2(n_212),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_3069),
.B(n_214),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_3065),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_3065),
.Y(n_3290)
);

AOI22x1_ASAP7_75t_L g3291 ( 
.A1(n_3143),
.A2(n_217),
.B1(n_215),
.B2(n_216),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_3065),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_3065),
.Y(n_3293)
);

INVx2_ASAP7_75t_L g3294 ( 
.A(n_3148),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_3065),
.Y(n_3295)
);

AOI21xp5_ASAP7_75t_L g3296 ( 
.A1(n_3119),
.A2(n_217),
.B(n_218),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_3065),
.Y(n_3297)
);

OAI22xp33_ASAP7_75t_L g3298 ( 
.A1(n_3123),
.A2(n_220),
.B1(n_218),
.B2(n_219),
.Y(n_3298)
);

OAI21xp33_ASAP7_75t_L g3299 ( 
.A1(n_3089),
.A2(n_219),
.B(n_220),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_3065),
.Y(n_3300)
);

OAI22xp5_ASAP7_75t_L g3301 ( 
.A1(n_3064),
.A2(n_224),
.B1(n_222),
.B2(n_223),
.Y(n_3301)
);

AOI22xp5_ASAP7_75t_L g3302 ( 
.A1(n_3064),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.Y(n_3302)
);

NOR2xp33_ASAP7_75t_L g3303 ( 
.A(n_3136),
.B(n_225),
.Y(n_3303)
);

INVxp67_ASAP7_75t_L g3304 ( 
.A(n_3151),
.Y(n_3304)
);

HB1xp67_ASAP7_75t_L g3305 ( 
.A(n_3156),
.Y(n_3305)
);

OAI21xp33_ASAP7_75t_L g3306 ( 
.A1(n_3089),
.A2(n_226),
.B(n_227),
.Y(n_3306)
);

INVx2_ASAP7_75t_L g3307 ( 
.A(n_3148),
.Y(n_3307)
);

INVx2_ASAP7_75t_SL g3308 ( 
.A(n_3122),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3065),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_3069),
.B(n_227),
.Y(n_3310)
);

AOI21xp33_ASAP7_75t_L g3311 ( 
.A1(n_3136),
.A2(n_228),
.B(n_229),
.Y(n_3311)
);

OAI22xp5_ASAP7_75t_L g3312 ( 
.A1(n_3064),
.A2(n_230),
.B1(n_228),
.B2(n_229),
.Y(n_3312)
);

AO22x1_ASAP7_75t_L g3313 ( 
.A1(n_3151),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_3187),
.B(n_231),
.Y(n_3314)
);

INVx2_ASAP7_75t_L g3315 ( 
.A(n_3187),
.Y(n_3315)
);

AOI22xp5_ASAP7_75t_L g3316 ( 
.A1(n_3172),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.Y(n_3316)
);

INVx2_ASAP7_75t_L g3317 ( 
.A(n_3258),
.Y(n_3317)
);

NAND3xp33_ASAP7_75t_L g3318 ( 
.A(n_3254),
.B(n_234),
.C(n_236),
.Y(n_3318)
);

INVx2_ASAP7_75t_SL g3319 ( 
.A(n_3237),
.Y(n_3319)
);

INVx2_ASAP7_75t_SL g3320 ( 
.A(n_3305),
.Y(n_3320)
);

OAI22xp33_ASAP7_75t_L g3321 ( 
.A1(n_3247),
.A2(n_238),
.B1(n_236),
.B2(n_237),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_L g3322 ( 
.A(n_3269),
.B(n_238),
.Y(n_3322)
);

OAI22xp33_ASAP7_75t_L g3323 ( 
.A1(n_3255),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_3323)
);

AOI22xp5_ASAP7_75t_L g3324 ( 
.A1(n_3177),
.A2(n_243),
.B1(n_239),
.B2(n_242),
.Y(n_3324)
);

O2A1O1Ixp33_ASAP7_75t_L g3325 ( 
.A1(n_3304),
.A2(n_245),
.B(n_243),
.C(n_244),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_L g3326 ( 
.A(n_3308),
.B(n_244),
.Y(n_3326)
);

NAND3xp33_ASAP7_75t_L g3327 ( 
.A(n_3160),
.B(n_3174),
.C(n_3280),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_3159),
.Y(n_3328)
);

NOR2xp33_ASAP7_75t_L g3329 ( 
.A(n_3174),
.B(n_246),
.Y(n_3329)
);

AOI22xp5_ASAP7_75t_L g3330 ( 
.A1(n_3201),
.A2(n_3282),
.B1(n_3286),
.B2(n_3229),
.Y(n_3330)
);

OAI21xp33_ASAP7_75t_SL g3331 ( 
.A1(n_3173),
.A2(n_246),
.B(n_247),
.Y(n_3331)
);

AND2x2_ASAP7_75t_L g3332 ( 
.A(n_3158),
.B(n_248),
.Y(n_3332)
);

INVx1_ASAP7_75t_SL g3333 ( 
.A(n_3183),
.Y(n_3333)
);

OAI22xp5_ASAP7_75t_L g3334 ( 
.A1(n_3277),
.A2(n_251),
.B1(n_248),
.B2(n_250),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_3162),
.Y(n_3335)
);

OAI22xp5_ASAP7_75t_L g3336 ( 
.A1(n_3285),
.A2(n_254),
.B1(n_250),
.B2(n_252),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_3249),
.Y(n_3337)
);

INVx1_ASAP7_75t_L g3338 ( 
.A(n_3250),
.Y(n_3338)
);

OAI22xp5_ASAP7_75t_L g3339 ( 
.A1(n_3264),
.A2(n_257),
.B1(n_252),
.B2(n_255),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_3252),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_3253),
.Y(n_3341)
);

AOI211xp5_ASAP7_75t_L g3342 ( 
.A1(n_3313),
.A2(n_259),
.B(n_257),
.C(n_258),
.Y(n_3342)
);

AOI22xp5_ASAP7_75t_L g3343 ( 
.A1(n_3190),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_3343)
);

AOI21xp33_ASAP7_75t_L g3344 ( 
.A1(n_3294),
.A2(n_261),
.B(n_262),
.Y(n_3344)
);

INVx3_ASAP7_75t_L g3345 ( 
.A(n_3195),
.Y(n_3345)
);

OAI22xp5_ASAP7_75t_SL g3346 ( 
.A1(n_3265),
.A2(n_263),
.B1(n_261),
.B2(n_262),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_3175),
.B(n_3166),
.Y(n_3347)
);

INVx1_ASAP7_75t_SL g3348 ( 
.A(n_3169),
.Y(n_3348)
);

AOI21xp33_ASAP7_75t_L g3349 ( 
.A1(n_3307),
.A2(n_264),
.B(n_265),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_L g3350 ( 
.A(n_3194),
.B(n_264),
.Y(n_3350)
);

OR2x2_ASAP7_75t_L g3351 ( 
.A(n_3259),
.B(n_266),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3260),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_L g3353 ( 
.A(n_3275),
.B(n_266),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_L g3354 ( 
.A(n_3281),
.B(n_267),
.Y(n_3354)
);

AOI21xp33_ASAP7_75t_L g3355 ( 
.A1(n_3188),
.A2(n_3289),
.B(n_3284),
.Y(n_3355)
);

AOI22xp5_ASAP7_75t_L g3356 ( 
.A1(n_3262),
.A2(n_269),
.B1(n_267),
.B2(n_268),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3290),
.Y(n_3357)
);

AND2x2_ASAP7_75t_L g3358 ( 
.A(n_3213),
.B(n_269),
.Y(n_3358)
);

OAI22xp5_ASAP7_75t_L g3359 ( 
.A1(n_3266),
.A2(n_3302),
.B1(n_3276),
.B2(n_3267),
.Y(n_3359)
);

INVx2_ASAP7_75t_L g3360 ( 
.A(n_3292),
.Y(n_3360)
);

NOR2xp33_ASAP7_75t_L g3361 ( 
.A(n_3161),
.B(n_270),
.Y(n_3361)
);

NOR2xp33_ASAP7_75t_L g3362 ( 
.A(n_3222),
.B(n_270),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_SL g3363 ( 
.A(n_3167),
.B(n_3279),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_L g3364 ( 
.A(n_3293),
.B(n_271),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_3295),
.Y(n_3365)
);

AOI322xp5_ASAP7_75t_L g3366 ( 
.A1(n_3268),
.A2(n_3309),
.A3(n_3297),
.B1(n_3300),
.B2(n_3299),
.C1(n_3306),
.C2(n_3251),
.Y(n_3366)
);

OAI21xp5_ASAP7_75t_L g3367 ( 
.A1(n_3296),
.A2(n_271),
.B(n_272),
.Y(n_3367)
);

INVx2_ASAP7_75t_SL g3368 ( 
.A(n_3163),
.Y(n_3368)
);

INVx1_ASAP7_75t_L g3369 ( 
.A(n_3178),
.Y(n_3369)
);

OAI211xp5_ASAP7_75t_L g3370 ( 
.A1(n_3263),
.A2(n_274),
.B(n_272),
.C(n_273),
.Y(n_3370)
);

O2A1O1Ixp33_ASAP7_75t_L g3371 ( 
.A1(n_3165),
.A2(n_276),
.B(n_274),
.C(n_275),
.Y(n_3371)
);

INVx2_ASAP7_75t_L g3372 ( 
.A(n_3192),
.Y(n_3372)
);

OR2x2_ASAP7_75t_L g3373 ( 
.A(n_3180),
.B(n_275),
.Y(n_3373)
);

OAI21xp5_ASAP7_75t_L g3374 ( 
.A1(n_3231),
.A2(n_276),
.B(n_277),
.Y(n_3374)
);

INVx1_ASAP7_75t_L g3375 ( 
.A(n_3257),
.Y(n_3375)
);

AND2x2_ASAP7_75t_L g3376 ( 
.A(n_3185),
.B(n_277),
.Y(n_3376)
);

INVx1_ASAP7_75t_SL g3377 ( 
.A(n_3181),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_L g3378 ( 
.A(n_3270),
.B(n_3182),
.Y(n_3378)
);

INVxp67_ASAP7_75t_SL g3379 ( 
.A(n_3268),
.Y(n_3379)
);

OAI32xp33_ASAP7_75t_L g3380 ( 
.A1(n_3230),
.A2(n_280),
.A3(n_278),
.B1(n_279),
.B2(n_281),
.Y(n_3380)
);

OAI221xp5_ASAP7_75t_L g3381 ( 
.A1(n_3283),
.A2(n_280),
.B1(n_278),
.B2(n_279),
.C(n_282),
.Y(n_3381)
);

OAI211xp5_ASAP7_75t_L g3382 ( 
.A1(n_3278),
.A2(n_284),
.B(n_282),
.C(n_283),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_L g3383 ( 
.A(n_3186),
.B(n_284),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_3261),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_L g3385 ( 
.A(n_3226),
.B(n_285),
.Y(n_3385)
);

OAI211xp5_ASAP7_75t_L g3386 ( 
.A1(n_3242),
.A2(n_288),
.B(n_286),
.C(n_287),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3288),
.Y(n_3387)
);

HB1xp67_ASAP7_75t_L g3388 ( 
.A(n_3164),
.Y(n_3388)
);

INVx2_ASAP7_75t_L g3389 ( 
.A(n_3291),
.Y(n_3389)
);

OR2x2_ASAP7_75t_L g3390 ( 
.A(n_3228),
.B(n_286),
.Y(n_3390)
);

INVx1_ASAP7_75t_L g3391 ( 
.A(n_3310),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_3236),
.Y(n_3392)
);

INVx1_ASAP7_75t_SL g3393 ( 
.A(n_3207),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_3272),
.B(n_287),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_3239),
.Y(n_3395)
);

AOI21xp33_ASAP7_75t_L g3396 ( 
.A1(n_3216),
.A2(n_288),
.B(n_289),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_3233),
.Y(n_3397)
);

NOR2xp33_ASAP7_75t_L g3398 ( 
.A(n_3197),
.B(n_289),
.Y(n_3398)
);

INVx1_ASAP7_75t_SL g3399 ( 
.A(n_3240),
.Y(n_3399)
);

INVxp67_ASAP7_75t_L g3400 ( 
.A(n_3303),
.Y(n_3400)
);

AOI22xp5_ASAP7_75t_L g3401 ( 
.A1(n_3301),
.A2(n_3312),
.B1(n_3189),
.B2(n_3198),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_3170),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_3217),
.B(n_290),
.Y(n_3403)
);

AOI21xp33_ASAP7_75t_SL g3404 ( 
.A1(n_3271),
.A2(n_290),
.B(n_291),
.Y(n_3404)
);

AOI221xp5_ASAP7_75t_L g3405 ( 
.A1(n_3227),
.A2(n_294),
.B1(n_292),
.B2(n_293),
.C(n_295),
.Y(n_3405)
);

AND2x2_ASAP7_75t_L g3406 ( 
.A(n_3184),
.B(n_292),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_3196),
.Y(n_3407)
);

INVx2_ASAP7_75t_L g3408 ( 
.A(n_3202),
.Y(n_3408)
);

XNOR2x2_ASAP7_75t_L g3409 ( 
.A(n_3246),
.B(n_294),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3208),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_3209),
.Y(n_3411)
);

AND2x2_ASAP7_75t_L g3412 ( 
.A(n_3218),
.B(n_295),
.Y(n_3412)
);

O2A1O1Ixp33_ASAP7_75t_L g3413 ( 
.A1(n_3199),
.A2(n_298),
.B(n_296),
.C(n_297),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_3210),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_3211),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_3238),
.Y(n_3416)
);

AND2x2_ASAP7_75t_L g3417 ( 
.A(n_3219),
.B(n_299),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_3243),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_3235),
.Y(n_3419)
);

INVx1_ASAP7_75t_L g3420 ( 
.A(n_3241),
.Y(n_3420)
);

NAND2xp33_ASAP7_75t_SL g3421 ( 
.A(n_3256),
.B(n_300),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_3244),
.Y(n_3422)
);

AOI21xp33_ASAP7_75t_SL g3423 ( 
.A1(n_3273),
.A2(n_3298),
.B(n_3287),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_SL g3424 ( 
.A(n_3193),
.B(n_3157),
.Y(n_3424)
);

INVx1_ASAP7_75t_L g3425 ( 
.A(n_3224),
.Y(n_3425)
);

OAI21xp5_ASAP7_75t_L g3426 ( 
.A1(n_3203),
.A2(n_300),
.B(n_302),
.Y(n_3426)
);

INVx2_ASAP7_75t_L g3427 ( 
.A(n_3176),
.Y(n_3427)
);

AOI31xp33_ASAP7_75t_L g3428 ( 
.A1(n_3248),
.A2(n_306),
.A3(n_304),
.B(n_305),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_3220),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_3168),
.Y(n_3430)
);

AND2x2_ASAP7_75t_L g3431 ( 
.A(n_3223),
.B(n_304),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_L g3432 ( 
.A(n_3215),
.B(n_305),
.Y(n_3432)
);

OAI22xp5_ASAP7_75t_L g3433 ( 
.A1(n_3221),
.A2(n_309),
.B1(n_307),
.B2(n_308),
.Y(n_3433)
);

OAI22xp5_ASAP7_75t_L g3434 ( 
.A1(n_3245),
.A2(n_309),
.B1(n_307),
.B2(n_308),
.Y(n_3434)
);

OAI211xp5_ASAP7_75t_L g3435 ( 
.A1(n_3205),
.A2(n_312),
.B(n_310),
.C(n_311),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3234),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_3204),
.B(n_310),
.Y(n_3437)
);

NAND4xp25_ASAP7_75t_L g3438 ( 
.A(n_3200),
.B(n_314),
.C(n_311),
.D(n_312),
.Y(n_3438)
);

OAI22xp5_ASAP7_75t_L g3439 ( 
.A1(n_3191),
.A2(n_317),
.B1(n_315),
.B2(n_316),
.Y(n_3439)
);

AND2x2_ASAP7_75t_L g3440 ( 
.A(n_3377),
.B(n_3232),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_3379),
.Y(n_3441)
);

AND2x2_ASAP7_75t_L g3442 ( 
.A(n_3319),
.B(n_3317),
.Y(n_3442)
);

INVxp67_ASAP7_75t_L g3443 ( 
.A(n_3421),
.Y(n_3443)
);

OR2x2_ASAP7_75t_L g3444 ( 
.A(n_3320),
.B(n_3225),
.Y(n_3444)
);

INVx1_ASAP7_75t_L g3445 ( 
.A(n_3315),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_3347),
.Y(n_3446)
);

AOI22xp33_ASAP7_75t_L g3447 ( 
.A1(n_3327),
.A2(n_3274),
.B1(n_3311),
.B2(n_3212),
.Y(n_3447)
);

INVx1_ASAP7_75t_L g3448 ( 
.A(n_3388),
.Y(n_3448)
);

AOI21xp5_ASAP7_75t_L g3449 ( 
.A1(n_3363),
.A2(n_3214),
.B(n_3179),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_3314),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_L g3451 ( 
.A(n_3348),
.B(n_3171),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_3322),
.Y(n_3452)
);

XNOR2x2_ASAP7_75t_L g3453 ( 
.A(n_3409),
.B(n_3405),
.Y(n_3453)
);

OAI21xp33_ASAP7_75t_L g3454 ( 
.A1(n_3330),
.A2(n_3206),
.B(n_317),
.Y(n_3454)
);

NAND2xp5_ASAP7_75t_L g3455 ( 
.A(n_3333),
.B(n_318),
.Y(n_3455)
);

OR2x2_ASAP7_75t_L g3456 ( 
.A(n_3378),
.B(n_318),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_L g3457 ( 
.A(n_3345),
.B(n_319),
.Y(n_3457)
);

OAI21xp33_ASAP7_75t_L g3458 ( 
.A1(n_3366),
.A2(n_319),
.B(n_320),
.Y(n_3458)
);

AOI21xp5_ASAP7_75t_L g3459 ( 
.A1(n_3371),
.A2(n_320),
.B(n_321),
.Y(n_3459)
);

NOR3xp33_ASAP7_75t_SL g3460 ( 
.A(n_3355),
.B(n_321),
.C(n_323),
.Y(n_3460)
);

NOR2xp33_ASAP7_75t_L g3461 ( 
.A(n_3345),
.B(n_325),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_L g3462 ( 
.A(n_3389),
.B(n_3361),
.Y(n_3462)
);

XOR2x2_ASAP7_75t_L g3463 ( 
.A(n_3336),
.B(n_326),
.Y(n_3463)
);

NOR2xp33_ASAP7_75t_L g3464 ( 
.A(n_3382),
.B(n_326),
.Y(n_3464)
);

AND2x2_ASAP7_75t_L g3465 ( 
.A(n_3328),
.B(n_327),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_L g3466 ( 
.A(n_3342),
.B(n_327),
.Y(n_3466)
);

OAI22xp33_ASAP7_75t_L g3467 ( 
.A1(n_3428),
.A2(n_330),
.B1(n_328),
.B2(n_329),
.Y(n_3467)
);

OAI21xp5_ASAP7_75t_SL g3468 ( 
.A1(n_3401),
.A2(n_328),
.B(n_331),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_3326),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_L g3470 ( 
.A(n_3368),
.B(n_331),
.Y(n_3470)
);

INVxp67_ASAP7_75t_L g3471 ( 
.A(n_3329),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3376),
.Y(n_3472)
);

OAI32xp33_ASAP7_75t_L g3473 ( 
.A1(n_3393),
.A2(n_334),
.A3(n_332),
.B1(n_333),
.B2(n_335),
.Y(n_3473)
);

AOI322xp5_ASAP7_75t_L g3474 ( 
.A1(n_3429),
.A2(n_337),
.A3(n_336),
.B1(n_334),
.B2(n_332),
.C1(n_333),
.C2(n_335),
.Y(n_3474)
);

NOR2xp33_ASAP7_75t_SL g3475 ( 
.A(n_3399),
.B(n_336),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3332),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_3351),
.Y(n_3477)
);

AOI21xp33_ASAP7_75t_SL g3478 ( 
.A1(n_3413),
.A2(n_338),
.B(n_339),
.Y(n_3478)
);

AOI22xp5_ASAP7_75t_L g3479 ( 
.A1(n_3359),
.A2(n_341),
.B1(n_338),
.B2(n_339),
.Y(n_3479)
);

AOI33xp33_ASAP7_75t_L g3480 ( 
.A1(n_3430),
.A2(n_344),
.A3(n_346),
.B1(n_341),
.B2(n_342),
.B3(n_345),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3358),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_3404),
.B(n_3392),
.Y(n_3482)
);

NOR2xp33_ASAP7_75t_L g3483 ( 
.A(n_3386),
.B(n_342),
.Y(n_3483)
);

AOI22xp33_ASAP7_75t_L g3484 ( 
.A1(n_3427),
.A2(n_348),
.B1(n_345),
.B2(n_347),
.Y(n_3484)
);

AOI22xp5_ASAP7_75t_L g3485 ( 
.A1(n_3436),
.A2(n_353),
.B1(n_347),
.B2(n_352),
.Y(n_3485)
);

OAI221xp5_ASAP7_75t_L g3486 ( 
.A1(n_3374),
.A2(n_3337),
.B1(n_3340),
.B2(n_3338),
.C(n_3335),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3373),
.Y(n_3487)
);

NAND2x1p5_ASAP7_75t_L g3488 ( 
.A(n_3372),
.B(n_352),
.Y(n_3488)
);

NOR2xp33_ASAP7_75t_L g3489 ( 
.A(n_3350),
.B(n_353),
.Y(n_3489)
);

OAI22xp5_ASAP7_75t_L g3490 ( 
.A1(n_3356),
.A2(n_356),
.B1(n_354),
.B2(n_355),
.Y(n_3490)
);

AOI221xp5_ASAP7_75t_L g3491 ( 
.A1(n_3423),
.A2(n_359),
.B1(n_354),
.B2(n_358),
.C(n_361),
.Y(n_3491)
);

INVx1_ASAP7_75t_SL g3492 ( 
.A(n_3390),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_L g3493 ( 
.A(n_3404),
.B(n_359),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3353),
.Y(n_3494)
);

AND2x2_ASAP7_75t_L g3495 ( 
.A(n_3406),
.B(n_3417),
.Y(n_3495)
);

HB1xp67_ASAP7_75t_L g3496 ( 
.A(n_3331),
.Y(n_3496)
);

AOI33xp33_ASAP7_75t_L g3497 ( 
.A1(n_3341),
.A2(n_363),
.A3(n_366),
.B1(n_361),
.B2(n_362),
.B3(n_365),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_3398),
.B(n_3360),
.Y(n_3498)
);

OAI21xp5_ASAP7_75t_L g3499 ( 
.A1(n_3370),
.A2(n_362),
.B(n_363),
.Y(n_3499)
);

AND2x2_ASAP7_75t_L g3500 ( 
.A(n_3431),
.B(n_365),
.Y(n_3500)
);

OAI22xp5_ASAP7_75t_L g3501 ( 
.A1(n_3381),
.A2(n_368),
.B1(n_366),
.B2(n_367),
.Y(n_3501)
);

AND2x2_ASAP7_75t_L g3502 ( 
.A(n_3400),
.B(n_369),
.Y(n_3502)
);

INVxp67_ASAP7_75t_L g3503 ( 
.A(n_3362),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_L g3504 ( 
.A(n_3412),
.B(n_371),
.Y(n_3504)
);

INVx2_ASAP7_75t_L g3505 ( 
.A(n_3352),
.Y(n_3505)
);

OAI221xp5_ASAP7_75t_L g3506 ( 
.A1(n_3357),
.A2(n_373),
.B1(n_371),
.B2(n_372),
.C(n_374),
.Y(n_3506)
);

AOI32xp33_ASAP7_75t_L g3507 ( 
.A1(n_3365),
.A2(n_376),
.A3(n_372),
.B1(n_374),
.B2(n_378),
.Y(n_3507)
);

OAI21xp5_ASAP7_75t_L g3508 ( 
.A1(n_3325),
.A2(n_378),
.B(n_379),
.Y(n_3508)
);

INVx1_ASAP7_75t_L g3509 ( 
.A(n_3354),
.Y(n_3509)
);

OAI22xp5_ASAP7_75t_L g3510 ( 
.A1(n_3346),
.A2(n_383),
.B1(n_380),
.B2(n_382),
.Y(n_3510)
);

NAND2xp33_ASAP7_75t_L g3511 ( 
.A(n_3403),
.B(n_382),
.Y(n_3511)
);

A2O1A1Ixp33_ASAP7_75t_L g3512 ( 
.A1(n_3435),
.A2(n_386),
.B(n_384),
.C(n_385),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3408),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3364),
.Y(n_3514)
);

NOR2xp33_ASAP7_75t_L g3515 ( 
.A(n_3438),
.B(n_385),
.Y(n_3515)
);

OR2x2_ASAP7_75t_L g3516 ( 
.A(n_3383),
.B(n_386),
.Y(n_3516)
);

AOI22xp33_ASAP7_75t_L g3517 ( 
.A1(n_3425),
.A2(n_389),
.B1(n_387),
.B2(n_388),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_SL g3518 ( 
.A(n_3321),
.B(n_387),
.Y(n_3518)
);

NOR2xp33_ASAP7_75t_L g3519 ( 
.A(n_3394),
.B(n_389),
.Y(n_3519)
);

NOR2xp33_ASAP7_75t_L g3520 ( 
.A(n_3344),
.B(n_3349),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_3385),
.Y(n_3521)
);

AOI21xp33_ASAP7_75t_L g3522 ( 
.A1(n_3395),
.A2(n_391),
.B(n_392),
.Y(n_3522)
);

INVxp67_ASAP7_75t_SL g3523 ( 
.A(n_3318),
.Y(n_3523)
);

NAND2xp5_ASAP7_75t_L g3524 ( 
.A(n_3323),
.B(n_391),
.Y(n_3524)
);

AOI221xp5_ASAP7_75t_L g3525 ( 
.A1(n_3380),
.A2(n_394),
.B1(n_392),
.B2(n_393),
.C(n_396),
.Y(n_3525)
);

NAND2xp5_ASAP7_75t_L g3526 ( 
.A(n_3369),
.B(n_393),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_L g3527 ( 
.A(n_3375),
.B(n_394),
.Y(n_3527)
);

OR2x2_ASAP7_75t_L g3528 ( 
.A(n_3384),
.B(n_396),
.Y(n_3528)
);

AOI221xp5_ASAP7_75t_L g3529 ( 
.A1(n_3424),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.C(n_400),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_L g3530 ( 
.A(n_3387),
.B(n_397),
.Y(n_3530)
);

OAI22xp5_ASAP7_75t_L g3531 ( 
.A1(n_3432),
.A2(n_401),
.B1(n_399),
.B2(n_400),
.Y(n_3531)
);

NOR2xp33_ASAP7_75t_L g3532 ( 
.A(n_3437),
.B(n_401),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3402),
.Y(n_3533)
);

NAND2x1_ASAP7_75t_L g3534 ( 
.A(n_3420),
.B(n_402),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3407),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3422),
.Y(n_3536)
);

AOI21x1_ASAP7_75t_L g3537 ( 
.A1(n_3410),
.A2(n_402),
.B(n_403),
.Y(n_3537)
);

OAI22xp5_ASAP7_75t_L g3538 ( 
.A1(n_3324),
.A2(n_406),
.B1(n_403),
.B2(n_404),
.Y(n_3538)
);

NAND2x1_ASAP7_75t_SL g3539 ( 
.A(n_3391),
.B(n_404),
.Y(n_3539)
);

AND2x2_ASAP7_75t_L g3540 ( 
.A(n_3367),
.B(n_407),
.Y(n_3540)
);

AOI22xp5_ASAP7_75t_L g3541 ( 
.A1(n_3334),
.A2(n_410),
.B1(n_408),
.B2(n_409),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_3397),
.B(n_409),
.Y(n_3542)
);

AOI21xp33_ASAP7_75t_SL g3543 ( 
.A1(n_3433),
.A2(n_411),
.B(n_412),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3411),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_L g3545 ( 
.A(n_3339),
.B(n_413),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_L g3546 ( 
.A(n_3419),
.B(n_414),
.Y(n_3546)
);

INVx2_ASAP7_75t_L g3547 ( 
.A(n_3414),
.Y(n_3547)
);

OAI22x1_ASAP7_75t_L g3548 ( 
.A1(n_3316),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.Y(n_3548)
);

INVx1_ASAP7_75t_L g3549 ( 
.A(n_3415),
.Y(n_3549)
);

INVxp67_ASAP7_75t_L g3550 ( 
.A(n_3426),
.Y(n_3550)
);

OAI22xp5_ASAP7_75t_L g3551 ( 
.A1(n_3343),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.Y(n_3551)
);

OAI22xp33_ASAP7_75t_L g3552 ( 
.A1(n_3439),
.A2(n_420),
.B1(n_418),
.B2(n_419),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_3434),
.B(n_418),
.Y(n_3553)
);

INVx1_ASAP7_75t_L g3554 ( 
.A(n_3416),
.Y(n_3554)
);

O2A1O1Ixp5_ASAP7_75t_L g3555 ( 
.A1(n_3418),
.A2(n_422),
.B(n_420),
.C(n_421),
.Y(n_3555)
);

INVx1_ASAP7_75t_SL g3556 ( 
.A(n_3396),
.Y(n_3556)
);

AOI22xp5_ASAP7_75t_L g3557 ( 
.A1(n_3421),
.A2(n_424),
.B1(n_422),
.B2(n_423),
.Y(n_3557)
);

A2O1A1Ixp33_ASAP7_75t_L g3558 ( 
.A1(n_3371),
.A2(n_426),
.B(n_423),
.C(n_425),
.Y(n_3558)
);

OR2x2_ASAP7_75t_L g3559 ( 
.A(n_3320),
.B(n_425),
.Y(n_3559)
);

AOI32xp33_ASAP7_75t_L g3560 ( 
.A1(n_3421),
.A2(n_429),
.A3(n_427),
.B1(n_428),
.B2(n_430),
.Y(n_3560)
);

INVx2_ASAP7_75t_L g3561 ( 
.A(n_3345),
.Y(n_3561)
);

AOI21xp33_ASAP7_75t_L g3562 ( 
.A1(n_3379),
.A2(n_427),
.B(n_429),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3379),
.Y(n_3563)
);

AND2x2_ASAP7_75t_L g3564 ( 
.A(n_3377),
.B(n_430),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3379),
.Y(n_3565)
);

AOI21xp33_ASAP7_75t_SL g3566 ( 
.A1(n_3320),
.A2(n_431),
.B(n_432),
.Y(n_3566)
);

AOI32xp33_ASAP7_75t_L g3567 ( 
.A1(n_3421),
.A2(n_435),
.A3(n_432),
.B1(n_433),
.B2(n_436),
.Y(n_3567)
);

OAI222xp33_ASAP7_75t_L g3568 ( 
.A1(n_3363),
.A2(n_437),
.B1(n_439),
.B2(n_433),
.C1(n_436),
.C2(n_438),
.Y(n_3568)
);

INVx1_ASAP7_75t_SL g3569 ( 
.A(n_3421),
.Y(n_3569)
);

HB1xp67_ASAP7_75t_L g3570 ( 
.A(n_3345),
.Y(n_3570)
);

XNOR2x2_ASAP7_75t_L g3571 ( 
.A(n_3409),
.B(n_438),
.Y(n_3571)
);

HB1xp67_ASAP7_75t_L g3572 ( 
.A(n_3345),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3379),
.Y(n_3573)
);

INVx2_ASAP7_75t_L g3574 ( 
.A(n_3345),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_3379),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3320),
.B(n_440),
.Y(n_3576)
);

OAI21xp33_ASAP7_75t_SL g3577 ( 
.A1(n_3379),
.A2(n_442),
.B(n_444),
.Y(n_3577)
);

INVx2_ASAP7_75t_SL g3578 ( 
.A(n_3345),
.Y(n_3578)
);

AOI222xp33_ASAP7_75t_L g3579 ( 
.A1(n_3363),
.A2(n_447),
.B1(n_449),
.B2(n_445),
.C1(n_446),
.C2(n_448),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3320),
.B(n_447),
.Y(n_3580)
);

AOI21xp33_ASAP7_75t_L g3581 ( 
.A1(n_3379),
.A2(n_448),
.B(n_449),
.Y(n_3581)
);

AND2x2_ASAP7_75t_SL g3582 ( 
.A(n_3389),
.B(n_450),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_3379),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3379),
.Y(n_3584)
);

AND2x2_ASAP7_75t_L g3585 ( 
.A(n_3377),
.B(n_450),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3379),
.Y(n_3586)
);

NOR3xp33_ASAP7_75t_L g3587 ( 
.A(n_3327),
.B(n_452),
.C(n_453),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3379),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_L g3589 ( 
.A(n_3320),
.B(n_453),
.Y(n_3589)
);

AOI32xp33_ASAP7_75t_L g3590 ( 
.A1(n_3421),
.A2(n_457),
.A3(n_455),
.B1(n_456),
.B2(n_458),
.Y(n_3590)
);

AOI21xp33_ASAP7_75t_L g3591 ( 
.A1(n_3379),
.A2(n_455),
.B(n_456),
.Y(n_3591)
);

AOI22xp5_ASAP7_75t_L g3592 ( 
.A1(n_3421),
.A2(n_459),
.B1(n_457),
.B2(n_458),
.Y(n_3592)
);

OAI21xp5_ASAP7_75t_L g3593 ( 
.A1(n_3327),
.A2(n_461),
.B(n_462),
.Y(n_3593)
);

AND2x2_ASAP7_75t_L g3594 ( 
.A(n_3377),
.B(n_463),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_3379),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_3320),
.B(n_464),
.Y(n_3596)
);

OAI21xp5_ASAP7_75t_L g3597 ( 
.A1(n_3443),
.A2(n_465),
.B(n_466),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3539),
.Y(n_3598)
);

AOI211xp5_ASAP7_75t_L g3599 ( 
.A1(n_3458),
.A2(n_468),
.B(n_465),
.C(n_467),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_L g3600 ( 
.A(n_3496),
.B(n_467),
.Y(n_3600)
);

NOR3x1_ASAP7_75t_L g3601 ( 
.A(n_3468),
.B(n_468),
.C(n_470),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_L g3602 ( 
.A(n_3569),
.B(n_470),
.Y(n_3602)
);

OAI322xp33_ASAP7_75t_L g3603 ( 
.A1(n_3453),
.A2(n_471),
.A3(n_472),
.B1(n_473),
.B2(n_474),
.C1(n_475),
.C2(n_476),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_SL g3604 ( 
.A(n_3475),
.B(n_475),
.Y(n_3604)
);

NOR3xp33_ASAP7_75t_SL g3605 ( 
.A(n_3486),
.B(n_3449),
.C(n_3482),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_L g3606 ( 
.A(n_3570),
.B(n_476),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_SL g3607 ( 
.A(n_3577),
.B(n_3560),
.Y(n_3607)
);

INVx1_ASAP7_75t_L g3608 ( 
.A(n_3572),
.Y(n_3608)
);

O2A1O1Ixp33_ASAP7_75t_L g3609 ( 
.A1(n_3568),
.A2(n_479),
.B(n_477),
.C(n_478),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_L g3610 ( 
.A(n_3578),
.B(n_477),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_L g3611 ( 
.A(n_3566),
.B(n_479),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3442),
.Y(n_3612)
);

OAI322xp33_ASAP7_75t_L g3613 ( 
.A1(n_3571),
.A2(n_480),
.A3(n_481),
.B1(n_482),
.B2(n_484),
.C1(n_485),
.C2(n_486),
.Y(n_3613)
);

NOR2xp33_ASAP7_75t_SL g3614 ( 
.A(n_3492),
.B(n_481),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3559),
.Y(n_3615)
);

NAND3xp33_ASAP7_75t_SL g3616 ( 
.A(n_3587),
.B(n_485),
.C(n_486),
.Y(n_3616)
);

NAND2xp5_ASAP7_75t_L g3617 ( 
.A(n_3566),
.B(n_487),
.Y(n_3617)
);

NOR4xp75_ASAP7_75t_L g3618 ( 
.A(n_3593),
.B(n_490),
.C(n_487),
.D(n_488),
.Y(n_3618)
);

BUFx2_ASAP7_75t_L g3619 ( 
.A(n_3488),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_3534),
.Y(n_3620)
);

OAI322xp33_ASAP7_75t_L g3621 ( 
.A1(n_3446),
.A2(n_491),
.A3(n_492),
.B1(n_493),
.B2(n_494),
.C1(n_495),
.C2(n_496),
.Y(n_3621)
);

NOR2xp33_ASAP7_75t_L g3622 ( 
.A(n_3478),
.B(n_493),
.Y(n_3622)
);

NAND3xp33_ASAP7_75t_SL g3623 ( 
.A(n_3478),
.B(n_495),
.C(n_496),
.Y(n_3623)
);

AOI221xp5_ASAP7_75t_L g3624 ( 
.A1(n_3447),
.A2(n_501),
.B1(n_497),
.B2(n_500),
.C(n_502),
.Y(n_3624)
);

NOR3xp33_ASAP7_75t_SL g3625 ( 
.A(n_3462),
.B(n_497),
.C(n_501),
.Y(n_3625)
);

AOI221xp5_ASAP7_75t_L g3626 ( 
.A1(n_3550),
.A2(n_504),
.B1(n_502),
.B2(n_503),
.C(n_505),
.Y(n_3626)
);

NAND3xp33_ASAP7_75t_L g3627 ( 
.A(n_3460),
.B(n_504),
.C(n_506),
.Y(n_3627)
);

OR2x2_ASAP7_75t_L g3628 ( 
.A(n_3444),
.B(n_506),
.Y(n_3628)
);

AND2x2_ASAP7_75t_L g3629 ( 
.A(n_3564),
.B(n_507),
.Y(n_3629)
);

NOR3xp33_ASAP7_75t_L g3630 ( 
.A(n_3454),
.B(n_3451),
.C(n_3498),
.Y(n_3630)
);

NOR3x1_ASAP7_75t_L g3631 ( 
.A(n_3499),
.B(n_3508),
.C(n_3523),
.Y(n_3631)
);

NOR3xp33_ASAP7_75t_L g3632 ( 
.A(n_3511),
.B(n_507),
.C(n_508),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3585),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_3594),
.Y(n_3634)
);

NOR2xp33_ASAP7_75t_L g3635 ( 
.A(n_3561),
.B(n_508),
.Y(n_3635)
);

NOR2xp33_ASAP7_75t_L g3636 ( 
.A(n_3574),
.B(n_510),
.Y(n_3636)
);

AND2x2_ASAP7_75t_L g3637 ( 
.A(n_3440),
.B(n_510),
.Y(n_3637)
);

INVx2_ASAP7_75t_L g3638 ( 
.A(n_3582),
.Y(n_3638)
);

INVxp67_ASAP7_75t_L g3639 ( 
.A(n_3483),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3537),
.Y(n_3640)
);

BUFx2_ASAP7_75t_L g3641 ( 
.A(n_3441),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_L g3642 ( 
.A(n_3567),
.B(n_511),
.Y(n_3642)
);

NOR2xp33_ASAP7_75t_L g3643 ( 
.A(n_3467),
.B(n_511),
.Y(n_3643)
);

NAND2xp5_ASAP7_75t_L g3644 ( 
.A(n_3590),
.B(n_512),
.Y(n_3644)
);

AND2x2_ASAP7_75t_L g3645 ( 
.A(n_3495),
.B(n_513),
.Y(n_3645)
);

OAI322xp33_ASAP7_75t_L g3646 ( 
.A1(n_3563),
.A2(n_513),
.A3(n_514),
.B1(n_516),
.B2(n_517),
.C1(n_518),
.C2(n_519),
.Y(n_3646)
);

AND2x2_ASAP7_75t_L g3647 ( 
.A(n_3476),
.B(n_516),
.Y(n_3647)
);

INVx2_ASAP7_75t_L g3648 ( 
.A(n_3500),
.Y(n_3648)
);

NAND2xp5_ASAP7_75t_L g3649 ( 
.A(n_3557),
.B(n_519),
.Y(n_3649)
);

AOI21xp5_ASAP7_75t_L g3650 ( 
.A1(n_3459),
.A2(n_520),
.B(n_521),
.Y(n_3650)
);

NOR2xp67_ASAP7_75t_L g3651 ( 
.A(n_3448),
.B(n_520),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_3592),
.B(n_521),
.Y(n_3652)
);

O2A1O1Ixp5_ASAP7_75t_SL g3653 ( 
.A1(n_3565),
.A2(n_525),
.B(n_522),
.C(n_523),
.Y(n_3653)
);

NOR3x1_ASAP7_75t_L g3654 ( 
.A(n_3455),
.B(n_522),
.C(n_526),
.Y(n_3654)
);

NOR2x1_ASAP7_75t_L g3655 ( 
.A(n_3573),
.B(n_526),
.Y(n_3655)
);

OR2x2_ASAP7_75t_L g3656 ( 
.A(n_3457),
.B(n_528),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_3465),
.Y(n_3657)
);

CKINVDCx5p33_ASAP7_75t_R g3658 ( 
.A(n_3463),
.Y(n_3658)
);

NOR2xp33_ASAP7_75t_L g3659 ( 
.A(n_3472),
.B(n_529),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3596),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_L g3661 ( 
.A(n_3575),
.B(n_529),
.Y(n_3661)
);

INVx1_ASAP7_75t_SL g3662 ( 
.A(n_3493),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_L g3663 ( 
.A(n_3583),
.B(n_530),
.Y(n_3663)
);

OA21x2_ASAP7_75t_L g3664 ( 
.A1(n_3584),
.A2(n_530),
.B(n_531),
.Y(n_3664)
);

NOR3x1_ASAP7_75t_L g3665 ( 
.A(n_3518),
.B(n_531),
.C(n_532),
.Y(n_3665)
);

AOI221xp5_ASAP7_75t_L g3666 ( 
.A1(n_3586),
.A2(n_533),
.B1(n_534),
.B2(n_535),
.C(n_536),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_3576),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3588),
.B(n_533),
.Y(n_3668)
);

CKINVDCx11_ASAP7_75t_R g3669 ( 
.A(n_3445),
.Y(n_3669)
);

INVx2_ASAP7_75t_L g3670 ( 
.A(n_3528),
.Y(n_3670)
);

NAND3xp33_ASAP7_75t_L g3671 ( 
.A(n_3595),
.B(n_535),
.C(n_537),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_L g3672 ( 
.A(n_3461),
.B(n_537),
.Y(n_3672)
);

NAND3xp33_ASAP7_75t_SL g3673 ( 
.A(n_3579),
.B(n_538),
.C(n_539),
.Y(n_3673)
);

AOI211xp5_ASAP7_75t_L g3674 ( 
.A1(n_3543),
.A2(n_541),
.B(n_538),
.C(n_540),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3580),
.Y(n_3675)
);

NOR2xp33_ASAP7_75t_L g3676 ( 
.A(n_3510),
.B(n_540),
.Y(n_3676)
);

O2A1O1Ixp33_ASAP7_75t_L g3677 ( 
.A1(n_3558),
.A2(n_543),
.B(n_541),
.C(n_542),
.Y(n_3677)
);

NAND3xp33_ASAP7_75t_L g3678 ( 
.A(n_3491),
.B(n_542),
.C(n_543),
.Y(n_3678)
);

NOR2xp33_ASAP7_75t_L g3679 ( 
.A(n_3481),
.B(n_544),
.Y(n_3679)
);

OAI21xp33_ASAP7_75t_L g3680 ( 
.A1(n_3520),
.A2(n_544),
.B(n_545),
.Y(n_3680)
);

AOI21xp5_ASAP7_75t_L g3681 ( 
.A1(n_3512),
.A2(n_3589),
.B(n_3466),
.Y(n_3681)
);

NAND3xp33_ASAP7_75t_SL g3682 ( 
.A(n_3556),
.B(n_546),
.C(n_548),
.Y(n_3682)
);

OR2x2_ASAP7_75t_L g3683 ( 
.A(n_3456),
.B(n_546),
.Y(n_3683)
);

OAI322xp33_ASAP7_75t_L g3684 ( 
.A1(n_3536),
.A2(n_549),
.A3(n_550),
.B1(n_551),
.B2(n_553),
.C1(n_554),
.C2(n_555),
.Y(n_3684)
);

HB1xp67_ASAP7_75t_L g3685 ( 
.A(n_3548),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3470),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_3504),
.Y(n_3687)
);

AOI221xp5_ASAP7_75t_L g3688 ( 
.A1(n_3487),
.A2(n_550),
.B1(n_551),
.B2(n_553),
.C(n_554),
.Y(n_3688)
);

NOR2x1_ASAP7_75t_L g3689 ( 
.A(n_3477),
.B(n_555),
.Y(n_3689)
);

NOR3x1_ASAP7_75t_L g3690 ( 
.A(n_3501),
.B(n_556),
.C(n_557),
.Y(n_3690)
);

AOI221xp5_ASAP7_75t_L g3691 ( 
.A1(n_3603),
.A2(n_3613),
.B1(n_3605),
.B2(n_3608),
.C(n_3609),
.Y(n_3691)
);

O2A1O1Ixp5_ASAP7_75t_L g3692 ( 
.A1(n_3607),
.A2(n_3505),
.B(n_3513),
.C(n_3547),
.Y(n_3692)
);

AOI22xp33_ASAP7_75t_L g3693 ( 
.A1(n_3669),
.A2(n_3452),
.B1(n_3469),
.B2(n_3494),
.Y(n_3693)
);

OAI211xp5_ASAP7_75t_L g3694 ( 
.A1(n_3598),
.A2(n_3525),
.B(n_3471),
.C(n_3503),
.Y(n_3694)
);

OAI211xp5_ASAP7_75t_L g3695 ( 
.A1(n_3620),
.A2(n_3535),
.B(n_3549),
.C(n_3544),
.Y(n_3695)
);

NOR3xp33_ASAP7_75t_L g3696 ( 
.A(n_3639),
.B(n_3450),
.C(n_3509),
.Y(n_3696)
);

OAI211xp5_ASAP7_75t_L g3697 ( 
.A1(n_3600),
.A2(n_3554),
.B(n_3479),
.C(n_3533),
.Y(n_3697)
);

NOR3xp33_ASAP7_75t_L g3698 ( 
.A(n_3630),
.B(n_3673),
.C(n_3619),
.Y(n_3698)
);

NOR2xp67_ASAP7_75t_SL g3699 ( 
.A(n_3612),
.B(n_3516),
.Y(n_3699)
);

OAI221xp5_ASAP7_75t_L g3700 ( 
.A1(n_3641),
.A2(n_3507),
.B1(n_3529),
.B2(n_3484),
.C(n_3514),
.Y(n_3700)
);

OAI22xp5_ASAP7_75t_L g3701 ( 
.A1(n_3627),
.A2(n_3485),
.B1(n_3541),
.B2(n_3464),
.Y(n_3701)
);

NOR3xp33_ASAP7_75t_L g3702 ( 
.A(n_3616),
.B(n_3521),
.C(n_3489),
.Y(n_3702)
);

OAI221xp5_ASAP7_75t_L g3703 ( 
.A1(n_3685),
.A2(n_3546),
.B1(n_3542),
.B2(n_3527),
.C(n_3530),
.Y(n_3703)
);

AOI322xp5_ASAP7_75t_L g3704 ( 
.A1(n_3623),
.A2(n_3515),
.A3(n_3540),
.B1(n_3532),
.B2(n_3519),
.C1(n_3524),
.C2(n_3552),
.Y(n_3704)
);

AOI222xp33_ASAP7_75t_L g3705 ( 
.A1(n_3640),
.A2(n_3531),
.B1(n_3490),
.B2(n_3538),
.C1(n_3551),
.C2(n_3545),
.Y(n_3705)
);

NOR2xp33_ASAP7_75t_L g3706 ( 
.A(n_3614),
.B(n_3562),
.Y(n_3706)
);

AOI221xp5_ASAP7_75t_L g3707 ( 
.A1(n_3682),
.A2(n_3473),
.B1(n_3581),
.B2(n_3591),
.C(n_3555),
.Y(n_3707)
);

NAND4xp75_ASAP7_75t_L g3708 ( 
.A(n_3631),
.B(n_3502),
.C(n_3526),
.D(n_3553),
.Y(n_3708)
);

O2A1O1Ixp33_ASAP7_75t_L g3709 ( 
.A1(n_3677),
.A2(n_3522),
.B(n_3506),
.C(n_3517),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_L g3710 ( 
.A(n_3651),
.B(n_3645),
.Y(n_3710)
);

AOI211xp5_ASAP7_75t_SL g3711 ( 
.A1(n_3681),
.A2(n_3480),
.B(n_3474),
.C(n_3497),
.Y(n_3711)
);

OAI21xp33_ASAP7_75t_L g3712 ( 
.A1(n_3658),
.A2(n_556),
.B(n_559),
.Y(n_3712)
);

AOI21xp5_ASAP7_75t_L g3713 ( 
.A1(n_3604),
.A2(n_560),
.B(n_561),
.Y(n_3713)
);

NOR3xp33_ASAP7_75t_L g3714 ( 
.A(n_3638),
.B(n_561),
.C(n_562),
.Y(n_3714)
);

AOI211xp5_ASAP7_75t_L g3715 ( 
.A1(n_3678),
.A2(n_564),
.B(n_562),
.C(n_563),
.Y(n_3715)
);

OAI22xp5_ASAP7_75t_L g3716 ( 
.A1(n_3602),
.A2(n_568),
.B1(n_563),
.B2(n_565),
.Y(n_3716)
);

AOI21xp33_ASAP7_75t_SL g3717 ( 
.A1(n_3622),
.A2(n_3632),
.B(n_3664),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_L g3718 ( 
.A(n_3629),
.B(n_568),
.Y(n_3718)
);

AOI22xp5_ASAP7_75t_L g3719 ( 
.A1(n_3633),
.A2(n_571),
.B1(n_569),
.B2(n_570),
.Y(n_3719)
);

OAI21xp5_ASAP7_75t_L g3720 ( 
.A1(n_3650),
.A2(n_573),
.B(n_574),
.Y(n_3720)
);

INVx2_ASAP7_75t_L g3721 ( 
.A(n_3664),
.Y(n_3721)
);

AOI211xp5_ASAP7_75t_L g3722 ( 
.A1(n_3634),
.A2(n_576),
.B(n_574),
.C(n_575),
.Y(n_3722)
);

AOI21xp5_ASAP7_75t_L g3723 ( 
.A1(n_3611),
.A2(n_575),
.B(n_576),
.Y(n_3723)
);

NAND2xp5_ASAP7_75t_L g3724 ( 
.A(n_3637),
.B(n_579),
.Y(n_3724)
);

NOR2xp67_ASAP7_75t_L g3725 ( 
.A(n_3671),
.B(n_581),
.Y(n_3725)
);

OAI21xp33_ASAP7_75t_L g3726 ( 
.A1(n_3648),
.A2(n_582),
.B(n_583),
.Y(n_3726)
);

AOI211xp5_ASAP7_75t_L g3727 ( 
.A1(n_3597),
.A2(n_3628),
.B(n_3662),
.C(n_3643),
.Y(n_3727)
);

OAI211xp5_ASAP7_75t_L g3728 ( 
.A1(n_3599),
.A2(n_584),
.B(n_582),
.C(n_583),
.Y(n_3728)
);

XNOR2x1_ASAP7_75t_L g3729 ( 
.A(n_3618),
.B(n_585),
.Y(n_3729)
);

NAND3xp33_ASAP7_75t_L g3730 ( 
.A(n_3625),
.B(n_585),
.C(n_586),
.Y(n_3730)
);

AND2x2_ASAP7_75t_L g3731 ( 
.A(n_3657),
.B(n_586),
.Y(n_3731)
);

OAI221xp5_ASAP7_75t_L g3732 ( 
.A1(n_3610),
.A2(n_587),
.B1(n_588),
.B2(n_591),
.C(n_592),
.Y(n_3732)
);

OAI21xp5_ASAP7_75t_SL g3733 ( 
.A1(n_3615),
.A2(n_587),
.B(n_588),
.Y(n_3733)
);

AOI211x1_ASAP7_75t_L g3734 ( 
.A1(n_3606),
.A2(n_593),
.B(n_591),
.C(n_592),
.Y(n_3734)
);

AOI221x1_ASAP7_75t_L g3735 ( 
.A1(n_3661),
.A2(n_593),
.B1(n_594),
.B2(n_595),
.C(n_596),
.Y(n_3735)
);

O2A1O1Ixp33_ASAP7_75t_L g3736 ( 
.A1(n_3617),
.A2(n_3644),
.B(n_3642),
.C(n_3646),
.Y(n_3736)
);

OAI21xp5_ASAP7_75t_L g3737 ( 
.A1(n_3689),
.A2(n_594),
.B(n_595),
.Y(n_3737)
);

OR2x2_ASAP7_75t_L g3738 ( 
.A(n_3683),
.B(n_596),
.Y(n_3738)
);

NOR2xp33_ASAP7_75t_L g3739 ( 
.A(n_3680),
.B(n_597),
.Y(n_3739)
);

AOI322xp5_ASAP7_75t_L g3740 ( 
.A1(n_3655),
.A2(n_597),
.A3(n_598),
.B1(n_599),
.B2(n_600),
.C1(n_601),
.C2(n_602),
.Y(n_3740)
);

AOI21xp5_ASAP7_75t_L g3741 ( 
.A1(n_3663),
.A2(n_3668),
.B(n_3652),
.Y(n_3741)
);

INVxp67_ASAP7_75t_L g3742 ( 
.A(n_3676),
.Y(n_3742)
);

NAND4xp25_ASAP7_75t_L g3743 ( 
.A(n_3665),
.B(n_601),
.C(n_598),
.D(n_599),
.Y(n_3743)
);

OAI211xp5_ASAP7_75t_SL g3744 ( 
.A1(n_3660),
.A2(n_602),
.B(n_603),
.C(n_604),
.Y(n_3744)
);

O2A1O1Ixp33_ASAP7_75t_L g3745 ( 
.A1(n_3621),
.A2(n_603),
.B(n_604),
.C(n_605),
.Y(n_3745)
);

NOR3xp33_ASAP7_75t_L g3746 ( 
.A(n_3667),
.B(n_606),
.C(n_608),
.Y(n_3746)
);

AOI211xp5_ASAP7_75t_SL g3747 ( 
.A1(n_3635),
.A2(n_606),
.B(n_609),
.C(n_610),
.Y(n_3747)
);

NOR2xp33_ASAP7_75t_SL g3748 ( 
.A(n_3684),
.B(n_611),
.Y(n_3748)
);

NOR2xp33_ASAP7_75t_SL g3749 ( 
.A(n_3670),
.B(n_611),
.Y(n_3749)
);

AND2x2_ASAP7_75t_L g3750 ( 
.A(n_3601),
.B(n_614),
.Y(n_3750)
);

AOI211xp5_ASAP7_75t_L g3751 ( 
.A1(n_3636),
.A2(n_614),
.B(n_616),
.C(n_617),
.Y(n_3751)
);

AOI221xp5_ASAP7_75t_SL g3752 ( 
.A1(n_3686),
.A2(n_617),
.B1(n_619),
.B2(n_620),
.C(n_622),
.Y(n_3752)
);

AOI221xp5_ASAP7_75t_L g3753 ( 
.A1(n_3717),
.A2(n_3675),
.B1(n_3687),
.B2(n_3624),
.C(n_3666),
.Y(n_3753)
);

INVx2_ASAP7_75t_L g3754 ( 
.A(n_3721),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3750),
.Y(n_3755)
);

BUFx2_ASAP7_75t_L g3756 ( 
.A(n_3737),
.Y(n_3756)
);

AOI22xp5_ASAP7_75t_L g3757 ( 
.A1(n_3748),
.A2(n_3647),
.B1(n_3674),
.B2(n_3679),
.Y(n_3757)
);

INVx2_ASAP7_75t_L g3758 ( 
.A(n_3738),
.Y(n_3758)
);

OAI22x1_ASAP7_75t_L g3759 ( 
.A1(n_3730),
.A2(n_3659),
.B1(n_3649),
.B2(n_3672),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_3710),
.Y(n_3760)
);

OAI22xp5_ASAP7_75t_L g3761 ( 
.A1(n_3693),
.A2(n_3656),
.B1(n_3688),
.B2(n_3626),
.Y(n_3761)
);

NOR2x1_ASAP7_75t_L g3762 ( 
.A(n_3743),
.B(n_3654),
.Y(n_3762)
);

OAI22xp5_ASAP7_75t_L g3763 ( 
.A1(n_3700),
.A2(n_3742),
.B1(n_3729),
.B2(n_3691),
.Y(n_3763)
);

HB1xp67_ASAP7_75t_L g3764 ( 
.A(n_3725),
.Y(n_3764)
);

AOI221xp5_ASAP7_75t_L g3765 ( 
.A1(n_3701),
.A2(n_3690),
.B1(n_3653),
.B2(n_625),
.C(n_626),
.Y(n_3765)
);

AOI22x1_ASAP7_75t_L g3766 ( 
.A1(n_3705),
.A2(n_3711),
.B1(n_3747),
.B2(n_3723),
.Y(n_3766)
);

AOI31xp33_ASAP7_75t_L g3767 ( 
.A1(n_3727),
.A2(n_619),
.A3(n_622),
.B(n_625),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3731),
.Y(n_3768)
);

AOI22xp33_ASAP7_75t_L g3769 ( 
.A1(n_3698),
.A2(n_626),
.B1(n_627),
.B2(n_628),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_3724),
.Y(n_3770)
);

INVx2_ASAP7_75t_L g3771 ( 
.A(n_3692),
.Y(n_3771)
);

OAI22xp5_ASAP7_75t_SL g3772 ( 
.A1(n_3734),
.A2(n_629),
.B1(n_630),
.B2(n_631),
.Y(n_3772)
);

OAI22x1_ASAP7_75t_L g3773 ( 
.A1(n_3706),
.A2(n_629),
.B1(n_630),
.B2(n_631),
.Y(n_3773)
);

OAI22xp5_ASAP7_75t_L g3774 ( 
.A1(n_3715),
.A2(n_632),
.B1(n_633),
.B2(n_634),
.Y(n_3774)
);

AOI22xp5_ASAP7_75t_L g3775 ( 
.A1(n_3694),
.A2(n_633),
.B1(n_635),
.B2(n_636),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3718),
.Y(n_3776)
);

AO22x2_ASAP7_75t_L g3777 ( 
.A1(n_3708),
.A2(n_636),
.B1(n_637),
.B2(n_638),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3699),
.Y(n_3778)
);

AOI22xp5_ASAP7_75t_L g3779 ( 
.A1(n_3702),
.A2(n_637),
.B1(n_638),
.B2(n_639),
.Y(n_3779)
);

AOI221xp5_ASAP7_75t_L g3780 ( 
.A1(n_3745),
.A2(n_639),
.B1(n_641),
.B2(n_642),
.C(n_643),
.Y(n_3780)
);

INVx1_ASAP7_75t_SL g3781 ( 
.A(n_3749),
.Y(n_3781)
);

INVx2_ASAP7_75t_L g3782 ( 
.A(n_3703),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3726),
.Y(n_3783)
);

INVx1_ASAP7_75t_L g3784 ( 
.A(n_3712),
.Y(n_3784)
);

INVx1_ASAP7_75t_L g3785 ( 
.A(n_3716),
.Y(n_3785)
);

NAND4xp25_ASAP7_75t_SL g3786 ( 
.A(n_3707),
.B(n_641),
.C(n_643),
.D(n_644),
.Y(n_3786)
);

AO22x2_ASAP7_75t_L g3787 ( 
.A1(n_3735),
.A2(n_645),
.B1(n_646),
.B2(n_647),
.Y(n_3787)
);

AOI22xp33_ASAP7_75t_L g3788 ( 
.A1(n_3696),
.A2(n_645),
.B1(n_646),
.B2(n_648),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3739),
.Y(n_3789)
);

AOI211xp5_ASAP7_75t_SL g3790 ( 
.A1(n_3763),
.A2(n_3695),
.B(n_3697),
.C(n_3741),
.Y(n_3790)
);

AOI221xp5_ASAP7_75t_L g3791 ( 
.A1(n_3777),
.A2(n_3709),
.B1(n_3736),
.B2(n_3743),
.C(n_3720),
.Y(n_3791)
);

AOI221xp5_ASAP7_75t_L g3792 ( 
.A1(n_3777),
.A2(n_3728),
.B1(n_3713),
.B2(n_3744),
.C(n_3714),
.Y(n_3792)
);

AOI221xp5_ASAP7_75t_L g3793 ( 
.A1(n_3771),
.A2(n_3733),
.B1(n_3752),
.B2(n_3746),
.C(n_3732),
.Y(n_3793)
);

XOR2xp5_ASAP7_75t_L g3794 ( 
.A(n_3766),
.B(n_3719),
.Y(n_3794)
);

AOI221xp5_ASAP7_75t_SL g3795 ( 
.A1(n_3765),
.A2(n_3722),
.B1(n_3751),
.B2(n_3704),
.C(n_3740),
.Y(n_3795)
);

OAI211xp5_ASAP7_75t_SL g3796 ( 
.A1(n_3753),
.A2(n_648),
.B(n_650),
.C(n_651),
.Y(n_3796)
);

OAI221xp5_ASAP7_75t_L g3797 ( 
.A1(n_3775),
.A2(n_650),
.B1(n_652),
.B2(n_653),
.C(n_655),
.Y(n_3797)
);

NOR2xp33_ASAP7_75t_L g3798 ( 
.A(n_3786),
.B(n_653),
.Y(n_3798)
);

OAI31xp33_ASAP7_75t_L g3799 ( 
.A1(n_3787),
.A2(n_655),
.A3(n_656),
.B(n_657),
.Y(n_3799)
);

OAI211xp5_ASAP7_75t_SL g3800 ( 
.A1(n_3757),
.A2(n_656),
.B(n_657),
.C(n_659),
.Y(n_3800)
);

NAND3x1_ASAP7_75t_L g3801 ( 
.A(n_3762),
.B(n_659),
.C(n_660),
.Y(n_3801)
);

OAI211xp5_ASAP7_75t_SL g3802 ( 
.A1(n_3778),
.A2(n_661),
.B(n_662),
.C(n_663),
.Y(n_3802)
);

AOI222xp33_ASAP7_75t_L g3803 ( 
.A1(n_3754),
.A2(n_661),
.B1(n_665),
.B2(n_666),
.C1(n_667),
.C2(n_668),
.Y(n_3803)
);

OAI21xp5_ASAP7_75t_L g3804 ( 
.A1(n_3761),
.A2(n_668),
.B(n_670),
.Y(n_3804)
);

OAI21xp33_ASAP7_75t_L g3805 ( 
.A1(n_3755),
.A2(n_671),
.B(n_672),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_3787),
.Y(n_3806)
);

AOI211x1_ASAP7_75t_L g3807 ( 
.A1(n_3783),
.A2(n_671),
.B(n_673),
.C(n_675),
.Y(n_3807)
);

OAI221xp5_ASAP7_75t_L g3808 ( 
.A1(n_3780),
.A2(n_673),
.B1(n_675),
.B2(n_676),
.C(n_677),
.Y(n_3808)
);

AOI22xp33_ASAP7_75t_L g3809 ( 
.A1(n_3782),
.A2(n_676),
.B1(n_678),
.B2(n_679),
.Y(n_3809)
);

OAI311xp33_ASAP7_75t_L g3810 ( 
.A1(n_3791),
.A2(n_3793),
.A3(n_3792),
.B1(n_3806),
.C1(n_3784),
.Y(n_3810)
);

OA22x2_ASAP7_75t_L g3811 ( 
.A1(n_3794),
.A2(n_3772),
.B1(n_3781),
.B2(n_3759),
.Y(n_3811)
);

AOI22xp5_ASAP7_75t_L g3812 ( 
.A1(n_3798),
.A2(n_3760),
.B1(n_3768),
.B2(n_3795),
.Y(n_3812)
);

OAI311xp33_ASAP7_75t_L g3813 ( 
.A1(n_3804),
.A2(n_3785),
.A3(n_3789),
.B1(n_3776),
.C1(n_3770),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3801),
.Y(n_3814)
);

NAND2xp5_ASAP7_75t_L g3815 ( 
.A(n_3799),
.B(n_3767),
.Y(n_3815)
);

AOI21xp33_ASAP7_75t_L g3816 ( 
.A1(n_3808),
.A2(n_3764),
.B(n_3758),
.Y(n_3816)
);

OAI211xp5_ASAP7_75t_SL g3817 ( 
.A1(n_3790),
.A2(n_3769),
.B(n_3779),
.C(n_3788),
.Y(n_3817)
);

AOI211xp5_ASAP7_75t_L g3818 ( 
.A1(n_3796),
.A2(n_3800),
.B(n_3774),
.C(n_3797),
.Y(n_3818)
);

O2A1O1Ixp33_ASAP7_75t_L g3819 ( 
.A1(n_3802),
.A2(n_3756),
.B(n_3773),
.C(n_683),
.Y(n_3819)
);

OAI22xp5_ASAP7_75t_L g3820 ( 
.A1(n_3809),
.A2(n_680),
.B1(n_682),
.B2(n_684),
.Y(n_3820)
);

NOR3xp33_ASAP7_75t_L g3821 ( 
.A(n_3805),
.B(n_680),
.C(n_682),
.Y(n_3821)
);

O2A1O1Ixp33_ASAP7_75t_L g3822 ( 
.A1(n_3803),
.A2(n_3807),
.B(n_685),
.C(n_686),
.Y(n_3822)
);

AND2x4_ASAP7_75t_L g3823 ( 
.A(n_3814),
.B(n_3821),
.Y(n_3823)
);

CKINVDCx14_ASAP7_75t_R g3824 ( 
.A(n_3812),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_3811),
.Y(n_3825)
);

NAND2xp5_ASAP7_75t_L g3826 ( 
.A(n_3818),
.B(n_684),
.Y(n_3826)
);

O2A1O1Ixp33_ASAP7_75t_L g3827 ( 
.A1(n_3810),
.A2(n_686),
.B(n_687),
.C(n_688),
.Y(n_3827)
);

INVxp67_ASAP7_75t_L g3828 ( 
.A(n_3815),
.Y(n_3828)
);

INVxp67_ASAP7_75t_L g3829 ( 
.A(n_3820),
.Y(n_3829)
);

OAI211xp5_ASAP7_75t_L g3830 ( 
.A1(n_3816),
.A2(n_687),
.B(n_689),
.C(n_690),
.Y(n_3830)
);

OAI221xp5_ASAP7_75t_SL g3831 ( 
.A1(n_3819),
.A2(n_691),
.B1(n_692),
.B2(n_693),
.C(n_696),
.Y(n_3831)
);

OR2x2_ASAP7_75t_L g3832 ( 
.A(n_3813),
.B(n_692),
.Y(n_3832)
);

OAI21xp5_ASAP7_75t_L g3833 ( 
.A1(n_3827),
.A2(n_3822),
.B(n_3817),
.Y(n_3833)
);

AND3x4_ASAP7_75t_L g3834 ( 
.A(n_3823),
.B(n_693),
.C(n_696),
.Y(n_3834)
);

NAND2xp5_ASAP7_75t_L g3835 ( 
.A(n_3824),
.B(n_697),
.Y(n_3835)
);

AND4x1_ASAP7_75t_L g3836 ( 
.A(n_3825),
.B(n_3826),
.C(n_3831),
.D(n_3832),
.Y(n_3836)
);

NAND4xp25_ASAP7_75t_L g3837 ( 
.A(n_3828),
.B(n_698),
.C(n_699),
.D(n_700),
.Y(n_3837)
);

NOR3xp33_ASAP7_75t_L g3838 ( 
.A(n_3835),
.B(n_3830),
.C(n_3829),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_L g3839 ( 
.A(n_3833),
.B(n_698),
.Y(n_3839)
);

OAI221xp5_ASAP7_75t_R g3840 ( 
.A1(n_3836),
.A2(n_699),
.B1(n_701),
.B2(n_702),
.C(n_704),
.Y(n_3840)
);

XNOR2xp5_ASAP7_75t_L g3841 ( 
.A(n_3838),
.B(n_3834),
.Y(n_3841)
);

AOI211xp5_ASAP7_75t_L g3842 ( 
.A1(n_3841),
.A2(n_3839),
.B(n_3837),
.C(n_3840),
.Y(n_3842)
);

NAND4xp25_ASAP7_75t_L g3843 ( 
.A(n_3842),
.B(n_701),
.C(n_702),
.D(n_704),
.Y(n_3843)
);

A2O1A1Ixp33_ASAP7_75t_L g3844 ( 
.A1(n_3843),
.A2(n_706),
.B(n_707),
.C(n_709),
.Y(n_3844)
);

OAI22xp5_ASAP7_75t_SL g3845 ( 
.A1(n_3844),
.A2(n_707),
.B1(n_709),
.B2(n_710),
.Y(n_3845)
);

INVxp67_ASAP7_75t_SL g3846 ( 
.A(n_3845),
.Y(n_3846)
);

AOI22xp5_ASAP7_75t_L g3847 ( 
.A1(n_3846),
.A2(n_710),
.B1(n_711),
.B2(n_712),
.Y(n_3847)
);

AO21x2_ASAP7_75t_L g3848 ( 
.A1(n_3847),
.A2(n_712),
.B(n_713),
.Y(n_3848)
);

HB1xp67_ASAP7_75t_L g3849 ( 
.A(n_3848),
.Y(n_3849)
);

INVx1_ASAP7_75t_L g3850 ( 
.A(n_3848),
.Y(n_3850)
);

OR2x6_ASAP7_75t_L g3851 ( 
.A(n_3849),
.B(n_713),
.Y(n_3851)
);

AOI21xp5_ASAP7_75t_L g3852 ( 
.A1(n_3851),
.A2(n_3850),
.B(n_716),
.Y(n_3852)
);

AOI211xp5_ASAP7_75t_L g3853 ( 
.A1(n_3852),
.A2(n_715),
.B(n_717),
.C(n_718),
.Y(n_3853)
);


endmodule