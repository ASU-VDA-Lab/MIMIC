module fake_jpeg_3745_n_279 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_38),
.Y(n_55)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_31),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_48),
.Y(n_66)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_33),
.B(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_R g48 ( 
.A(n_33),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_15),
.B1(n_30),
.B2(n_18),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_49),
.A2(n_39),
.B1(n_37),
.B2(n_41),
.Y(n_77)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_54),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_51),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_30),
.B(n_15),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_59),
.C(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

HAxp5_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_29),
.CON(n_56),
.SN(n_56)
);

AOI32xp33_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_29),
.A3(n_17),
.B1(n_34),
.B2(n_35),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_24),
.B1(n_18),
.B2(n_27),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_59),
.A2(n_37),
.B1(n_33),
.B2(n_41),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_27),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_24),
.Y(n_67)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_71),
.Y(n_89)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_75),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_69),
.A2(n_23),
.B(n_26),
.Y(n_91)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_87),
.B1(n_45),
.B2(n_80),
.Y(n_92)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_79),
.B(n_60),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_40),
.B1(n_34),
.B2(n_35),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_64),
.B1(n_62),
.B2(n_60),
.Y(n_103)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_81),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_55),
.B1(n_64),
.B2(n_62),
.Y(n_100)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_52),
.A2(n_37),
.B1(n_41),
.B2(n_42),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_35),
.B(n_34),
.C(n_32),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_46),
.A2(n_61),
.B1(n_65),
.B2(n_50),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_80),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_90),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_55),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_106),
.B(n_67),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_92),
.A2(n_103),
.B1(n_82),
.B2(n_68),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_44),
.C(n_42),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_97),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_55),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_99),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_44),
.C(n_32),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_101),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_75),
.B(n_66),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_100),
.A2(n_108),
.B1(n_81),
.B2(n_83),
.Y(n_134)
);

BUFx12_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_109),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_69),
.A2(n_26),
.B(n_35),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_86),
.Y(n_129)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_111),
.A2(n_115),
.B(n_127),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_112),
.Y(n_143)
);

BUFx12_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_114),
.Y(n_144)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_106),
.A2(n_91),
.B(n_97),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_121),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_119),
.B(n_124),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_94),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_123),
.Y(n_139)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_109),
.B(n_66),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_89),
.B(n_66),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_128),
.A2(n_90),
.B1(n_104),
.B2(n_72),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_133),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_79),
.Y(n_130)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_73),
.Y(n_131)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_88),
.B(n_92),
.Y(n_132)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_78),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_134),
.A2(n_32),
.B1(n_84),
.B2(n_105),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_147),
.B1(n_149),
.B2(n_154),
.Y(n_162)
);

AND2x6_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_122),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_146),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_101),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_125),
.C(n_123),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_110),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_145),
.Y(n_174)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_34),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_128),
.A2(n_72),
.B1(n_96),
.B2(n_110),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_132),
.A2(n_96),
.B1(n_98),
.B2(n_32),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_126),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_114),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_151),
.A2(n_153),
.B1(n_157),
.B2(n_158),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_134),
.A2(n_84),
.B1(n_105),
.B2(n_20),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_115),
.A2(n_25),
.B1(n_29),
.B2(n_17),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_118),
.A2(n_25),
.B1(n_29),
.B2(n_17),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_102),
.B1(n_28),
.B2(n_22),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_122),
.A2(n_102),
.B1(n_28),
.B2(n_2),
.Y(n_159)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_159),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_111),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_165),
.C(n_169),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_144),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_164),
.Y(n_186)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_173),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_143),
.Y(n_164)
);

INVxp67_ASAP7_75t_SL g166 ( 
.A(n_145),
.Y(n_166)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_125),
.Y(n_169)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_126),
.Y(n_171)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_117),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_181),
.Y(n_187)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_178),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_117),
.B(n_133),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_177),
.A2(n_157),
.B(n_112),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_147),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_116),
.Y(n_179)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_179),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_149),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_182),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_113),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_151),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_113),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_154),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_180),
.A2(n_141),
.B1(n_156),
.B2(n_135),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_188),
.A2(n_194),
.B1(n_167),
.B2(n_163),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_168),
.B(n_139),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_195),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_160),
.A2(n_141),
.B1(n_153),
.B2(n_158),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_193),
.Y(n_217)
);

AND2x6_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_159),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_146),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_203),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_201),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_174),
.A2(n_112),
.B(n_28),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_1),
.Y(n_220)
);

MAJx2_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_181),
.C(n_165),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_0),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_204),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_199),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_208),
.Y(n_228)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_162),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_215),
.Y(n_233)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_190),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_212),
.Y(n_231)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_198),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_188),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_213),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_219),
.B1(n_189),
.B2(n_193),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_177),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_176),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_187),
.C(n_4),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_194),
.A2(n_173),
.B1(n_112),
.B2(n_3),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_220),
.A2(n_1),
.B(n_2),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_185),
.B(n_1),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_221),
.B(n_200),
.Y(n_226)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_184),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_2),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_224),
.A2(n_225),
.B(n_236),
.Y(n_248)
);

A2O1A1Ixp33_ASAP7_75t_SL g225 ( 
.A1(n_219),
.A2(n_197),
.B(n_196),
.C(n_203),
.Y(n_225)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_226),
.Y(n_238)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_214),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_227),
.B(n_232),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_229),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_205),
.B(n_195),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_230),
.Y(n_239)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_206),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_218),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_217),
.A2(n_187),
.B(n_4),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_237),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_240),
.B(n_225),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_215),
.C(n_216),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_6),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_206),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_7),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_245),
.B(n_246),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_210),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_14),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_4),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_249),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_250),
.B(n_256),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_239),
.A2(n_225),
.B1(n_236),
.B2(n_231),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_255),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_253),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_242),
.A2(n_225),
.B1(n_228),
.B2(n_235),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_254),
.A2(n_257),
.B(n_243),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_241),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_6),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_248),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_253),
.B(n_240),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_263),
.A2(n_265),
.B(n_266),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_252),
.Y(n_271)
);

AOI31xp33_ASAP7_75t_L g266 ( 
.A1(n_258),
.A2(n_248),
.A3(n_244),
.B(n_10),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_260),
.B(n_259),
.Y(n_267)
);

AO21x1_ASAP7_75t_L g272 ( 
.A1(n_267),
.A2(n_261),
.B(n_9),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_261),
.Y(n_268)
);

A2O1A1Ixp33_ASAP7_75t_L g273 ( 
.A1(n_268),
.A2(n_270),
.B(n_8),
.C(n_9),
.Y(n_273)
);

BUFx24_ASAP7_75t_SL g270 ( 
.A(n_262),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_9),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_272),
.B(n_273),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_274),
.A2(n_269),
.B(n_12),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_276),
.A2(n_275),
.B(n_12),
.Y(n_277)
);

AOI21x1_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_11),
.B(n_12),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_14),
.Y(n_279)
);


endmodule