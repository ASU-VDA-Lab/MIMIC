module fake_jpeg_31450_n_135 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_135);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_22),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_23),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_2),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_40),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_0),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_50),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_65),
.Y(n_72)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_48),
.B(n_1),
.Y(n_66)
);

AO22x1_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_57),
.B1(n_56),
.B2(n_54),
.Y(n_68)
);

AO22x1_ASAP7_75t_SL g67 ( 
.A1(n_61),
.A2(n_53),
.B1(n_44),
.B2(n_48),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_9),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_73),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_64),
.A2(n_54),
.B1(n_53),
.B2(n_44),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_58),
.C(n_66),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_43),
.B(n_52),
.C(n_56),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_74),
.A2(n_10),
.B(n_12),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_49),
.B1(n_57),
.B2(n_56),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_80),
.B1(n_3),
.B2(n_5),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_60),
.A2(n_57),
.B1(n_47),
.B2(n_4),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_78),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_47),
.B1(n_3),
.B2(n_5),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_47),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_82),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_1),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_6),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_86),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_8),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_96),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_68),
.B(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_8),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_90),
.A2(n_92),
.B1(n_95),
.B2(n_93),
.Y(n_99)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_97),
.Y(n_113)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_12),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_93),
.A2(n_70),
.B(n_76),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_99),
.Y(n_120)
);

AND2x6_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_25),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_112),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_90),
.A2(n_26),
.B1(n_41),
.B2(n_38),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_104),
.B1(n_109),
.B2(n_111),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_24),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_114),
.C(n_87),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_42),
.B1(n_21),
.B2(n_27),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_96),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_110),
.B(n_16),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_95),
.A2(n_20),
.B1(n_36),
.B2(n_35),
.Y(n_111)
);

OA21x2_ASAP7_75t_SL g112 ( 
.A1(n_92),
.A2(n_14),
.B(n_15),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_83),
.A2(n_17),
.B(n_18),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_115),
.B(n_117),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_84),
.C(n_19),
.Y(n_117)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_119),
.A2(n_121),
.B(n_114),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_29),
.C(n_30),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_16),
.B1(n_37),
.B2(n_107),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_123),
.A2(n_111),
.B1(n_106),
.B2(n_100),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_126),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_125),
.A2(n_120),
.B(n_98),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_116),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_130),
.B(n_115),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_131),
.B(n_127),
.Y(n_132)
);

AOI322xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_102),
.A3(n_127),
.B1(n_129),
.B2(n_117),
.C1(n_122),
.C2(n_105),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_101),
.C(n_104),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_101),
.Y(n_135)
);


endmodule