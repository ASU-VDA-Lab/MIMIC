module fake_jpeg_29001_n_143 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_143);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

BUFx3_ASAP7_75t_SL g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_24),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_21),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_23),
.Y(n_52)
);

BUFx4f_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_15),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_26),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_0),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_66),
.Y(n_72)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_46),
.B1(n_65),
.B2(n_49),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_37),
.B1(n_51),
.B2(n_54),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_70),
.A2(n_71),
.B1(n_75),
.B2(n_43),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_63),
.A2(n_44),
.B1(n_37),
.B2(n_54),
.Y(n_71)
);

AO22x2_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_46),
.B1(n_51),
.B2(n_48),
.Y(n_73)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_73),
.A2(n_76),
.B1(n_42),
.B2(n_41),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_68),
.A2(n_59),
.B1(n_58),
.B2(n_55),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_64),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_80),
.Y(n_83)
);

CKINVDCx5p33_ASAP7_75t_R g79 ( 
.A(n_64),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_45),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_64),
.Y(n_80)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_94),
.Y(n_108)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_87),
.B(n_3),
.Y(n_105)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_47),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_92),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_72),
.B(n_76),
.C(n_2),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_90),
.B(n_98),
.Y(n_106)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_0),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_96),
.B1(n_99),
.B2(n_1),
.Y(n_103)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_79),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_18),
.B1(n_34),
.B2(n_32),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_74),
.Y(n_101)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_118),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_3),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_112),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_85),
.B(n_4),
.Y(n_112)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_5),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_113),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_121),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_108),
.A2(n_107),
.B(n_106),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

NAND3xp33_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_127),
.C(n_128),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_6),
.Y(n_125)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_117),
.A2(n_12),
.B1(n_14),
.B2(n_16),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_114),
.C(n_117),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_114),
.C(n_123),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_135),
.B(n_136),
.Y(n_138)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_133),
.A2(n_124),
.B(n_122),
.Y(n_137)
);

NAND2xp33_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_137),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_134),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_140),
.B(n_130),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_119),
.B(n_111),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_142),
.B(n_104),
.Y(n_143)
);


endmodule