module fake_aes_7575_n_1033 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_225, n_39, n_1033);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1033;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_383;
wire n_288;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_572;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_975;
wire n_279;
wire n_303;
wire n_968;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_638;
wire n_563;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_1011;
wire n_1025;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1014;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_935;
wire n_427;
wire n_910;
wire n_950;
wire n_460;
wire n_478;
wire n_415;
wire n_482;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_990;
wire n_751;
wire n_800;
wire n_626;
wire n_941;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_475;
wire n_926;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_622;
wire n_549;
wire n_832;
wire n_262;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_446;
wire n_420;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_716;
wire n_653;
wire n_881;
wire n_806;
wire n_539;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_315;
wire n_409;
wire n_363;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_1029;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_811;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_924;
wire n_947;
wire n_912;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_992;
wire n_269;
INVx1_ASAP7_75t_L g262 ( .A(n_71), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g263 ( .A(n_94), .Y(n_263) );
INVxp67_ASAP7_75t_SL g264 ( .A(n_222), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_57), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_235), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_61), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_43), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_169), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_226), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_165), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_123), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_199), .Y(n_273) );
CKINVDCx20_ASAP7_75t_R g274 ( .A(n_180), .Y(n_274) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_14), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_108), .Y(n_276) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_252), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_166), .Y(n_278) );
BUFx2_ASAP7_75t_L g279 ( .A(n_48), .Y(n_279) );
CKINVDCx20_ASAP7_75t_R g280 ( .A(n_238), .Y(n_280) );
CKINVDCx20_ASAP7_75t_R g281 ( .A(n_41), .Y(n_281) );
INVx2_ASAP7_75t_SL g282 ( .A(n_137), .Y(n_282) );
BUFx3_ASAP7_75t_L g283 ( .A(n_40), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_202), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_58), .Y(n_285) );
CKINVDCx20_ASAP7_75t_R g286 ( .A(n_126), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g287 ( .A(n_152), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_259), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_92), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_175), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_221), .Y(n_291) );
CKINVDCx20_ASAP7_75t_R g292 ( .A(n_249), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_215), .Y(n_293) );
BUFx5_ASAP7_75t_L g294 ( .A(n_52), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_174), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_128), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_145), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_79), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_104), .B(n_254), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_187), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_229), .B(n_101), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_56), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_197), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_39), .Y(n_304) );
BUFx3_ASAP7_75t_L g305 ( .A(n_167), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_117), .Y(n_306) );
INVxp67_ASAP7_75t_L g307 ( .A(n_146), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_48), .Y(n_308) );
CKINVDCx20_ASAP7_75t_R g309 ( .A(n_39), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_260), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g311 ( .A(n_53), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_57), .Y(n_312) );
INVxp67_ASAP7_75t_L g313 ( .A(n_210), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_200), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_31), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_213), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_181), .Y(n_317) );
INVxp67_ASAP7_75t_L g318 ( .A(n_220), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_160), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_41), .Y(n_320) );
CKINVDCx20_ASAP7_75t_R g321 ( .A(n_115), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_141), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_256), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_147), .Y(n_324) );
BUFx3_ASAP7_75t_L g325 ( .A(n_77), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_120), .Y(n_326) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_228), .Y(n_327) );
CKINVDCx20_ASAP7_75t_R g328 ( .A(n_230), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_47), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_246), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_255), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_212), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_9), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_21), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_55), .Y(n_335) );
CKINVDCx20_ASAP7_75t_R g336 ( .A(n_25), .Y(n_336) );
INVxp67_ASAP7_75t_SL g337 ( .A(n_17), .Y(n_337) );
CKINVDCx20_ASAP7_75t_R g338 ( .A(n_185), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_5), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_258), .Y(n_340) );
BUFx3_ASAP7_75t_L g341 ( .A(n_82), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_14), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_84), .Y(n_343) );
CKINVDCx20_ASAP7_75t_R g344 ( .A(n_38), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_154), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_22), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_250), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_109), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_234), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_205), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_190), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_211), .Y(n_352) );
INVxp67_ASAP7_75t_SL g353 ( .A(n_36), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_184), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_121), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_203), .Y(n_356) );
BUFx3_ASAP7_75t_L g357 ( .A(n_7), .Y(n_357) );
CKINVDCx20_ASAP7_75t_R g358 ( .A(n_261), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_172), .Y(n_359) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_242), .Y(n_360) );
CKINVDCx20_ASAP7_75t_R g361 ( .A(n_257), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_98), .Y(n_362) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_72), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_12), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_183), .B(n_155), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_105), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_24), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_112), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_103), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_86), .Y(n_370) );
CKINVDCx20_ASAP7_75t_R g371 ( .A(n_171), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_247), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_162), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_135), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_33), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_218), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_214), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_26), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_149), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_251), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_248), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_25), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_21), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_23), .Y(n_384) );
BUFx3_ASAP7_75t_L g385 ( .A(n_12), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_179), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_66), .Y(n_387) );
CKINVDCx16_ASAP7_75t_R g388 ( .A(n_42), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_78), .Y(n_389) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_97), .Y(n_390) );
CKINVDCx16_ASAP7_75t_R g391 ( .A(n_388), .Y(n_391) );
INVx3_ASAP7_75t_L g392 ( .A(n_294), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_275), .Y(n_393) );
INVx4_ASAP7_75t_L g394 ( .A(n_305), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_294), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_294), .Y(n_396) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_327), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_327), .Y(n_398) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_327), .Y(n_399) );
NOR2xp33_ASAP7_75t_SL g400 ( .A(n_278), .B(n_80), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_294), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_294), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_279), .B(n_273), .Y(n_403) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_327), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_360), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_277), .B(n_0), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_360), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_360), .Y(n_408) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_283), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_360), .Y(n_410) );
AND2x4_ASAP7_75t_L g411 ( .A(n_283), .B(n_0), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_294), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_282), .B(n_1), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_294), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_312), .Y(n_415) );
OA21x2_ASAP7_75t_L g416 ( .A1(n_271), .A2(n_83), .B(n_81), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_262), .B(n_1), .Y(n_417) );
AOI22xp5_ASAP7_75t_SL g418 ( .A1(n_281), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_418) );
BUFx2_ASAP7_75t_L g419 ( .A(n_325), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_390), .Y(n_420) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_281), .A2(n_311), .B1(n_336), .B2(n_309), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_390), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_325), .B(n_2), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_390), .Y(n_424) );
BUFx2_ASAP7_75t_L g425 ( .A(n_357), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_390), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_312), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_411), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_411), .Y(n_429) );
NAND2xp5_ASAP7_75t_SL g430 ( .A(n_411), .B(n_271), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_419), .B(n_307), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_423), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_392), .B(n_272), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_419), .B(n_265), .Y(n_434) );
NOR2xp33_ASAP7_75t_SL g435 ( .A(n_400), .B(n_263), .Y(n_435) );
BUFx10_ASAP7_75t_L g436 ( .A(n_393), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_406), .A2(n_274), .B1(n_280), .B2(n_263), .Y(n_437) );
INVx4_ASAP7_75t_L g438 ( .A(n_394), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_425), .Y(n_439) );
AND3x2_ASAP7_75t_L g440 ( .A(n_425), .B(n_353), .C(n_337), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_409), .Y(n_441) );
AND3x2_ASAP7_75t_L g442 ( .A(n_406), .B(n_264), .C(n_267), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_403), .B(n_268), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_391), .A2(n_280), .B1(n_286), .B2(n_274), .Y(n_444) );
INVx3_ASAP7_75t_L g445 ( .A(n_392), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g446 ( .A(n_392), .B(n_272), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_391), .B(n_285), .Y(n_447) );
AND2x6_ASAP7_75t_L g448 ( .A(n_392), .B(n_305), .Y(n_448) );
BUFx3_ASAP7_75t_L g449 ( .A(n_394), .Y(n_449) );
OAI22xp33_ASAP7_75t_L g450 ( .A1(n_421), .A2(n_311), .B1(n_336), .B2(n_309), .Y(n_450) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_397), .Y(n_451) );
INVx5_ASAP7_75t_L g452 ( .A(n_394), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_394), .B(n_313), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_395), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_421), .B(n_302), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_395), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_415), .B(n_357), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_396), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_415), .B(n_318), .Y(n_459) );
INVx3_ASAP7_75t_L g460 ( .A(n_396), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_401), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_417), .A2(n_287), .B1(n_292), .B2(n_286), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_401), .Y(n_463) );
INVxp33_ASAP7_75t_L g464 ( .A(n_413), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_427), .B(n_304), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_402), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_402), .B(n_385), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g468 ( .A1(n_412), .A2(n_292), .B1(n_321), .B2(n_287), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_414), .Y(n_469) );
INVx3_ASAP7_75t_L g470 ( .A(n_414), .Y(n_470) );
OAI22xp33_ASAP7_75t_SL g471 ( .A1(n_418), .A2(n_339), .B1(n_346), .B2(n_320), .Y(n_471) );
INVx4_ASAP7_75t_L g472 ( .A(n_416), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_464), .B(n_284), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_464), .B(n_293), .Y(n_474) );
NOR2x1p5_ASAP7_75t_L g475 ( .A(n_447), .B(n_378), .Y(n_475) );
INVx2_ASAP7_75t_SL g476 ( .A(n_436), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_431), .B(n_297), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_444), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_436), .B(n_443), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_445), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_457), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_465), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_439), .A2(n_328), .B1(n_338), .B2(n_321), .Y(n_483) );
AND2x6_ASAP7_75t_SL g484 ( .A(n_450), .B(n_308), .Y(n_484) );
BUFx12f_ASAP7_75t_L g485 ( .A(n_436), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_434), .B(n_385), .Y(n_486) );
OR2x6_ASAP7_75t_L g487 ( .A(n_432), .B(n_387), .Y(n_487) );
NAND2xp33_ASAP7_75t_SL g488 ( .A(n_428), .B(n_328), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_431), .B(n_306), .Y(n_489) );
INVx2_ASAP7_75t_SL g490 ( .A(n_429), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_460), .B(n_266), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_459), .B(n_315), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_430), .A2(n_416), .B(n_289), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_460), .B(n_269), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_430), .A2(n_333), .B1(n_334), .B2(n_329), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_445), .Y(n_496) );
AND2x6_ASAP7_75t_SL g497 ( .A(n_471), .B(n_335), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_472), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_442), .B(n_342), .Y(n_499) );
BUFx3_ASAP7_75t_L g500 ( .A(n_448), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_470), .B(n_270), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_472), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_472), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_470), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_467), .B(n_314), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_453), .B(n_317), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_453), .B(n_322), .Y(n_507) );
AND3x1_ASAP7_75t_L g508 ( .A(n_437), .B(n_367), .C(n_364), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_433), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_448), .A2(n_375), .B1(n_383), .B2(n_382), .Y(n_510) );
AOI22xp33_ASAP7_75t_SL g511 ( .A1(n_435), .A2(n_344), .B1(n_358), .B2(n_338), .Y(n_511) );
BUFx3_ASAP7_75t_L g512 ( .A(n_448), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_438), .B(n_330), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_456), .Y(n_514) );
CKINVDCx11_ASAP7_75t_R g515 ( .A(n_462), .Y(n_515) );
OR2x6_ASAP7_75t_L g516 ( .A(n_455), .B(n_387), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_456), .B(n_276), .Y(n_517) );
NOR2x2_ASAP7_75t_L g518 ( .A(n_468), .B(n_344), .Y(n_518) );
INVx3_ASAP7_75t_L g519 ( .A(n_438), .Y(n_519) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_440), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_433), .B(n_384), .Y(n_521) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_446), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_461), .A2(n_363), .B1(n_361), .B2(n_358), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_452), .B(n_361), .Y(n_524) );
INVx3_ASAP7_75t_L g525 ( .A(n_449), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_454), .A2(n_295), .B(n_296), .C(n_290), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_458), .A2(n_363), .B1(n_371), .B2(n_369), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_463), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_466), .A2(n_363), .B1(n_371), .B2(n_369), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_469), .A2(n_363), .B1(n_416), .B2(n_300), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_452), .B(n_298), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_451), .B(n_303), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_451), .B(n_3), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_464), .B(n_345), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_457), .Y(n_535) );
INVx1_ASAP7_75t_SL g536 ( .A(n_436), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_436), .B(n_416), .Y(n_537) );
OAI22xp33_ASAP7_75t_L g538 ( .A1(n_468), .A2(n_310), .B1(n_319), .B2(n_316), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_441), .A2(n_324), .B1(n_326), .B2(n_323), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_428), .B(n_331), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_457), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_464), .B(n_348), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_457), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_464), .B(n_349), .Y(n_544) );
OAI22xp5_ASAP7_75t_SL g545 ( .A1(n_437), .A2(n_350), .B1(n_351), .B2(n_340), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_436), .B(n_341), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_436), .Y(n_547) );
INVx5_ASAP7_75t_L g548 ( .A(n_448), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_476), .B(n_352), .Y(n_549) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_490), .A2(n_356), .B(n_362), .C(n_354), .Y(n_550) );
OR2x4_ASAP7_75t_L g551 ( .A(n_542), .B(n_299), .Y(n_551) );
AOI33xp33_ASAP7_75t_L g552 ( .A1(n_482), .A2(n_379), .A3(n_366), .B1(n_368), .B2(n_370), .B3(n_373), .Y(n_552) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_500), .Y(n_553) );
OAI22xp5_ASAP7_75t_SL g554 ( .A1(n_508), .A2(n_377), .B1(n_380), .B2(n_374), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_479), .B(n_4), .Y(n_555) );
O2A1O1Ixp33_ASAP7_75t_L g556 ( .A1(n_526), .A2(n_386), .B(n_389), .C(n_381), .Y(n_556) );
O2A1O1Ixp33_ASAP7_75t_L g557 ( .A1(n_526), .A2(n_289), .B(n_291), .C(n_288), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_498), .A2(n_291), .B(n_288), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_476), .B(n_355), .Y(n_559) );
INVx4_ASAP7_75t_L g560 ( .A(n_485), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_502), .A2(n_343), .B(n_332), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_536), .B(n_359), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_490), .A2(n_365), .B1(n_372), .B2(n_332), .Y(n_563) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_547), .Y(n_564) );
BUFx2_ASAP7_75t_SL g565 ( .A(n_524), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_502), .A2(n_347), .B(n_343), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_503), .A2(n_376), .B(n_347), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_485), .B(n_5), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_503), .A2(n_301), .B(n_398), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_481), .Y(n_570) );
BUFx4f_ASAP7_75t_L g571 ( .A(n_487), .Y(n_571) );
OAI22x1_ASAP7_75t_L g572 ( .A1(n_483), .A2(n_8), .B1(n_6), .B2(n_7), .Y(n_572) );
AND2x4_ASAP7_75t_L g573 ( .A(n_487), .B(n_6), .Y(n_573) );
BUFx2_ASAP7_75t_SL g574 ( .A(n_524), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_473), .B(n_8), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_474), .B(n_9), .Y(n_576) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_515), .Y(n_577) );
AND2x4_ASAP7_75t_L g578 ( .A(n_487), .B(n_10), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_493), .A2(n_405), .B(n_398), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_546), .B(n_10), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_534), .B(n_11), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_545), .A2(n_487), .B1(n_516), .B2(n_488), .Y(n_582) );
A2O1A1Ixp33_ASAP7_75t_L g583 ( .A1(n_528), .A2(n_407), .B(n_408), .C(n_405), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_546), .B(n_11), .Y(n_584) );
BUFx3_ASAP7_75t_L g585 ( .A(n_535), .Y(n_585) );
BUFx2_ASAP7_75t_L g586 ( .A(n_488), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_516), .B(n_13), .Y(n_587) );
NAND3xp33_ASAP7_75t_L g588 ( .A(n_530), .B(n_399), .C(n_397), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_486), .B(n_13), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_541), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_516), .B(n_15), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_543), .Y(n_592) );
BUFx3_ASAP7_75t_L g593 ( .A(n_499), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g594 ( .A(n_515), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_544), .B(n_15), .Y(n_595) );
BUFx3_ASAP7_75t_L g596 ( .A(n_499), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_504), .Y(n_597) );
OAI22x1_ASAP7_75t_L g598 ( .A1(n_518), .A2(n_16), .B1(n_18), .B2(n_19), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_521), .Y(n_599) );
INVx3_ASAP7_75t_L g600 ( .A(n_519), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_511), .B(n_16), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_523), .A2(n_426), .B1(n_424), .B2(n_422), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_527), .A2(n_426), .B1(n_424), .B2(n_422), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_492), .B(n_18), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g605 ( .A1(n_537), .A2(n_410), .B(n_420), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_521), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_520), .B(n_477), .Y(n_607) );
INVx1_ASAP7_75t_SL g608 ( .A(n_537), .Y(n_608) );
INVx4_ASAP7_75t_L g609 ( .A(n_548), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_521), .Y(n_610) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_500), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_492), .B(n_19), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_495), .B(n_20), .Y(n_613) );
BUFx2_ASAP7_75t_L g614 ( .A(n_518), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_489), .B(n_20), .Y(n_615) );
O2A1O1Ixp33_ASAP7_75t_L g616 ( .A1(n_540), .A2(n_22), .B(n_23), .C(n_24), .Y(n_616) );
AND2x4_ASAP7_75t_L g617 ( .A(n_475), .B(n_26), .Y(n_617) );
BUFx2_ASAP7_75t_L g618 ( .A(n_484), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_480), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_480), .Y(n_620) );
O2A1O1Ixp33_ASAP7_75t_L g621 ( .A1(n_517), .A2(n_27), .B(n_28), .C(n_29), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_496), .Y(n_622) );
INVx2_ASAP7_75t_SL g623 ( .A(n_499), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_504), .Y(n_624) );
INVx4_ASAP7_75t_L g625 ( .A(n_512), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_529), .A2(n_404), .B1(n_399), .B2(n_30), .Y(n_626) );
CKINVDCx5p33_ASAP7_75t_R g627 ( .A(n_497), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_510), .A2(n_404), .B1(n_30), .B2(n_31), .Y(n_628) );
INVx3_ASAP7_75t_L g629 ( .A(n_519), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_505), .B(n_28), .Y(n_630) );
NOR2xp67_ASAP7_75t_L g631 ( .A(n_539), .B(n_32), .Y(n_631) );
A2O1A1Ixp33_ASAP7_75t_L g632 ( .A1(n_509), .A2(n_404), .B(n_35), .C(n_36), .Y(n_632) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_513), .B(n_34), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_496), .Y(n_634) );
OR2x6_ASAP7_75t_L g635 ( .A(n_522), .B(n_37), .Y(n_635) );
BUFx2_ASAP7_75t_L g636 ( .A(n_514), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_514), .Y(n_637) );
OR2x6_ASAP7_75t_SL g638 ( .A(n_506), .B(n_42), .Y(n_638) );
O2A1O1Ixp33_ASAP7_75t_L g639 ( .A1(n_491), .A2(n_43), .B(n_44), .C(n_45), .Y(n_639) );
INVx3_ASAP7_75t_L g640 ( .A(n_525), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_507), .B(n_44), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_491), .A2(n_46), .B1(n_49), .B2(n_50), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_494), .A2(n_49), .B1(n_50), .B2(n_51), .Y(n_643) );
AOI21xp5_ASAP7_75t_L g644 ( .A1(n_494), .A2(n_87), .B(n_85), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g645 ( .A1(n_501), .A2(n_89), .B(n_88), .Y(n_645) );
OR2x2_ASAP7_75t_L g646 ( .A(n_533), .B(n_53), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_531), .A2(n_54), .B1(n_55), .B2(n_56), .Y(n_647) );
INVx4_ASAP7_75t_L g648 ( .A(n_531), .Y(n_648) );
AOI21xp5_ASAP7_75t_L g649 ( .A1(n_532), .A2(n_91), .B(n_90), .Y(n_649) );
A2O1A1Ixp33_ASAP7_75t_L g650 ( .A1(n_490), .A2(n_58), .B(n_59), .C(n_60), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_479), .B(n_59), .Y(n_651) );
A2O1A1Ixp33_ASAP7_75t_L g652 ( .A1(n_490), .A2(n_60), .B(n_61), .C(n_62), .Y(n_652) );
OR2x2_ASAP7_75t_L g653 ( .A(n_564), .B(n_62), .Y(n_653) );
OAI21x1_ASAP7_75t_L g654 ( .A1(n_579), .A2(n_176), .B(n_253), .Y(n_654) );
OAI22xp33_ASAP7_75t_L g655 ( .A1(n_571), .A2(n_63), .B1(n_64), .B2(n_65), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_585), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_573), .A2(n_63), .B1(n_64), .B2(n_65), .Y(n_657) );
A2O1A1Ixp33_ASAP7_75t_L g658 ( .A1(n_641), .A2(n_66), .B(n_67), .C(n_68), .Y(n_658) );
OAI221xp5_ASAP7_75t_L g659 ( .A1(n_582), .A2(n_67), .B1(n_68), .B2(n_69), .C(n_70), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_636), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_555), .B(n_69), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_597), .Y(n_662) );
BUFx3_ASAP7_75t_L g663 ( .A(n_560), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_599), .B(n_72), .Y(n_664) );
AO32x2_ASAP7_75t_L g665 ( .A1(n_626), .A2(n_73), .A3(n_74), .B1(n_75), .B2(n_76), .Y(n_665) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_637), .A2(n_182), .B(n_245), .Y(n_666) );
O2A1O1Ixp33_ASAP7_75t_L g667 ( .A1(n_556), .A2(n_73), .B(n_74), .C(n_75), .Y(n_667) );
INVxp67_ASAP7_75t_SL g668 ( .A(n_571), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_573), .A2(n_76), .B1(n_77), .B2(n_93), .Y(n_669) );
A2O1A1Ixp33_ASAP7_75t_L g670 ( .A1(n_557), .A2(n_95), .B(n_96), .C(n_99), .Y(n_670) );
AOI21xp5_ASAP7_75t_L g671 ( .A1(n_588), .A2(n_100), .B(n_102), .Y(n_671) );
AOI22xp33_ASAP7_75t_SL g672 ( .A1(n_578), .A2(n_106), .B1(n_107), .B2(n_110), .Y(n_672) );
CKINVDCx11_ASAP7_75t_R g673 ( .A(n_560), .Y(n_673) );
INVx1_ASAP7_75t_SL g674 ( .A(n_578), .Y(n_674) );
OAI21x1_ASAP7_75t_L g675 ( .A1(n_558), .A2(n_111), .B(n_113), .Y(n_675) );
BUFx6f_ASAP7_75t_L g676 ( .A(n_553), .Y(n_676) );
A2O1A1Ixp33_ASAP7_75t_L g677 ( .A1(n_615), .A2(n_114), .B(n_116), .C(n_118), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_570), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_624), .Y(n_679) );
OAI21x1_ASAP7_75t_L g680 ( .A1(n_561), .A2(n_119), .B(n_122), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_591), .A2(n_554), .B1(n_587), .B2(n_574), .Y(n_681) );
OAI21x1_ASAP7_75t_L g682 ( .A1(n_566), .A2(n_124), .B(n_125), .Y(n_682) );
OAI22xp33_ASAP7_75t_L g683 ( .A1(n_635), .A2(n_127), .B1(n_129), .B2(n_130), .Y(n_683) );
A2O1A1Ixp33_ASAP7_75t_L g684 ( .A1(n_595), .A2(n_131), .B(n_132), .C(n_133), .Y(n_684) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_635), .Y(n_685) );
CKINVDCx11_ASAP7_75t_R g686 ( .A(n_638), .Y(n_686) );
O2A1O1Ixp33_ASAP7_75t_L g687 ( .A1(n_550), .A2(n_134), .B(n_136), .C(n_138), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_590), .Y(n_688) );
AO31x2_ASAP7_75t_L g689 ( .A1(n_632), .A2(n_139), .A3(n_140), .B(n_142), .Y(n_689) );
OAI21x1_ASAP7_75t_L g690 ( .A1(n_567), .A2(n_143), .B(n_144), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_634), .Y(n_691) );
A2O1A1Ixp33_ASAP7_75t_L g692 ( .A1(n_575), .A2(n_148), .B(n_150), .C(n_151), .Y(n_692) );
AND2x4_ASAP7_75t_L g693 ( .A(n_623), .B(n_153), .Y(n_693) );
O2A1O1Ixp33_ASAP7_75t_L g694 ( .A1(n_604), .A2(n_156), .B(n_157), .C(n_158), .Y(n_694) );
NAND2x2_ASAP7_75t_L g695 ( .A(n_598), .B(n_159), .Y(n_695) );
AOI21xp5_ASAP7_75t_L g696 ( .A1(n_619), .A2(n_161), .B(n_163), .Y(n_696) );
BUFx8_ASAP7_75t_L g697 ( .A(n_614), .Y(n_697) );
OAI21x1_ASAP7_75t_L g698 ( .A1(n_569), .A2(n_164), .B(n_168), .Y(n_698) );
AOI21xp5_ASAP7_75t_L g699 ( .A1(n_620), .A2(n_170), .B(n_173), .Y(n_699) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_622), .A2(n_177), .B(n_178), .Y(n_700) );
INVx1_ASAP7_75t_SL g701 ( .A(n_635), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_592), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_608), .A2(n_186), .B1(n_188), .B2(n_189), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_551), .B(n_191), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g705 ( .A1(n_608), .A2(n_192), .B1(n_193), .B2(n_194), .Y(n_705) );
AO31x2_ASAP7_75t_L g706 ( .A1(n_583), .A2(n_195), .A3(n_196), .B(n_198), .Y(n_706) );
INVx1_ASAP7_75t_SL g707 ( .A(n_593), .Y(n_707) );
BUFx2_ASAP7_75t_L g708 ( .A(n_596), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_606), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_651), .A2(n_201), .B1(n_204), .B2(n_206), .Y(n_710) );
BUFx6f_ASAP7_75t_L g711 ( .A(n_553), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_610), .Y(n_712) );
A2O1A1Ixp33_ASAP7_75t_L g713 ( .A1(n_576), .A2(n_207), .B(n_208), .C(n_209), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_612), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_646), .A2(n_216), .B1(n_217), .B2(n_219), .Y(n_715) );
A2O1A1Ixp33_ASAP7_75t_L g716 ( .A1(n_581), .A2(n_223), .B(n_224), .C(n_225), .Y(n_716) );
A2O1A1Ixp33_ASAP7_75t_L g717 ( .A1(n_552), .A2(n_616), .B(n_639), .C(n_621), .Y(n_717) );
O2A1O1Ixp33_ASAP7_75t_SL g718 ( .A1(n_633), .A2(n_227), .B(n_231), .C(n_232), .Y(n_718) );
AO31x2_ASAP7_75t_L g719 ( .A1(n_650), .A2(n_233), .A3(n_236), .B(n_237), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_613), .Y(n_720) );
AO31x2_ASAP7_75t_L g721 ( .A1(n_652), .A2(n_239), .A3(n_240), .B(n_241), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g722 ( .A1(n_630), .A2(n_243), .B(n_244), .Y(n_722) );
OR2x2_ASAP7_75t_L g723 ( .A(n_618), .B(n_554), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_551), .B(n_607), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_565), .A2(n_601), .B1(n_586), .B2(n_617), .Y(n_725) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_563), .A2(n_589), .B1(n_580), .B2(n_584), .Y(n_726) );
AO32x2_ASAP7_75t_L g727 ( .A1(n_602), .A2(n_603), .A3(n_643), .B1(n_642), .B2(n_628), .Y(n_727) );
INVx1_ASAP7_75t_SL g728 ( .A(n_568), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_631), .B(n_562), .Y(n_729) );
NOR2xp33_ASAP7_75t_SL g730 ( .A(n_577), .B(n_594), .Y(n_730) );
AO31x2_ASAP7_75t_L g731 ( .A1(n_572), .A2(n_644), .A3(n_645), .B(n_649), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_617), .A2(n_600), .B1(n_629), .B2(n_640), .Y(n_732) );
AND2x4_ASAP7_75t_L g733 ( .A(n_549), .B(n_559), .Y(n_733) );
A2O1A1Ixp33_ASAP7_75t_L g734 ( .A1(n_647), .A2(n_611), .B(n_627), .C(n_648), .Y(n_734) );
INVxp67_ASAP7_75t_SL g735 ( .A(n_625), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_625), .Y(n_736) );
NOR2xp67_ASAP7_75t_L g737 ( .A(n_609), .B(n_476), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_636), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_585), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_564), .B(n_479), .Y(n_740) );
AND2x4_ASAP7_75t_L g741 ( .A(n_560), .B(n_476), .Y(n_741) );
BUFx12f_ASAP7_75t_L g742 ( .A(n_560), .Y(n_742) );
NOR2xp67_ASAP7_75t_L g743 ( .A(n_573), .B(n_476), .Y(n_743) );
O2A1O1Ixp33_ASAP7_75t_L g744 ( .A1(n_556), .A2(n_526), .B(n_550), .C(n_478), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_585), .Y(n_745) );
BUFx2_ASAP7_75t_L g746 ( .A(n_564), .Y(n_746) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_573), .A2(n_444), .B1(n_479), .B2(n_485), .Y(n_747) );
OAI22xp33_ASAP7_75t_L g748 ( .A1(n_571), .A2(n_444), .B1(n_437), .B2(n_462), .Y(n_748) );
BUFx8_ASAP7_75t_SL g749 ( .A(n_577), .Y(n_749) );
INVx2_ASAP7_75t_L g750 ( .A(n_636), .Y(n_750) );
AOI322xp5_ASAP7_75t_L g751 ( .A1(n_614), .A2(n_450), .A3(n_421), .B1(n_478), .B2(n_582), .C1(n_538), .C2(n_618), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_585), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_573), .A2(n_478), .B1(n_479), .B2(n_545), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_571), .A2(n_578), .B1(n_573), .B2(n_608), .Y(n_754) );
OAI21xp5_ASAP7_75t_L g755 ( .A1(n_605), .A2(n_502), .B(n_498), .Y(n_755) );
AND2x4_ASAP7_75t_L g756 ( .A(n_560), .B(n_476), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_573), .A2(n_478), .B1(n_479), .B2(n_545), .Y(n_757) );
AOI221xp5_ASAP7_75t_L g758 ( .A1(n_554), .A2(n_450), .B1(n_508), .B2(n_538), .C(n_545), .Y(n_758) );
OAI21xp5_ASAP7_75t_L g759 ( .A1(n_605), .A2(n_502), .B(n_498), .Y(n_759) );
A2O1A1Ixp33_ASAP7_75t_L g760 ( .A1(n_641), .A2(n_557), .B(n_615), .C(n_595), .Y(n_760) );
AO31x2_ASAP7_75t_L g761 ( .A1(n_579), .A2(n_493), .A3(n_472), .B(n_632), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_585), .Y(n_762) );
AO221x2_ASAP7_75t_L g763 ( .A1(n_598), .A2(n_450), .B1(n_554), .B2(n_572), .C(n_444), .Y(n_763) );
A2O1A1Ixp33_ASAP7_75t_L g764 ( .A1(n_641), .A2(n_557), .B(n_615), .C(n_595), .Y(n_764) );
AO31x2_ASAP7_75t_L g765 ( .A1(n_579), .A2(n_493), .A3(n_472), .B(n_632), .Y(n_765) );
INVx2_ASAP7_75t_L g766 ( .A(n_678), .Y(n_766) );
AND2x2_ASAP7_75t_L g767 ( .A(n_753), .B(n_757), .Y(n_767) );
HB1xp67_ASAP7_75t_L g768 ( .A(n_746), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g769 ( .A1(n_763), .A2(n_754), .B1(n_758), .B2(n_724), .Y(n_769) );
AOI21xp5_ASAP7_75t_L g770 ( .A1(n_755), .A2(n_759), .B(n_726), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_714), .B(n_720), .Y(n_771) );
AO31x2_ASAP7_75t_L g772 ( .A1(n_717), .A2(n_670), .A3(n_671), .B(n_684), .Y(n_772) );
BUFx6f_ASAP7_75t_L g773 ( .A(n_676), .Y(n_773) );
BUFx6f_ASAP7_75t_L g774 ( .A(n_676), .Y(n_774) );
AO31x2_ASAP7_75t_L g775 ( .A1(n_734), .A2(n_677), .A3(n_692), .B(n_713), .Y(n_775) );
INVx2_ASAP7_75t_SL g776 ( .A(n_742), .Y(n_776) );
OA21x2_ASAP7_75t_L g777 ( .A1(n_654), .A2(n_698), .B(n_690), .Y(n_777) );
OAI21xp33_ASAP7_75t_L g778 ( .A1(n_751), .A2(n_729), .B(n_747), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_688), .B(n_702), .Y(n_779) );
OA21x2_ASAP7_75t_L g780 ( .A1(n_675), .A2(n_680), .B(n_682), .Y(n_780) );
AND2x4_ASAP7_75t_L g781 ( .A(n_743), .B(n_668), .Y(n_781) );
AO31x2_ASAP7_75t_L g782 ( .A1(n_716), .A2(n_715), .A3(n_703), .B(n_705), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_660), .Y(n_783) );
AOI22xp5_ASAP7_75t_L g784 ( .A1(n_763), .A2(n_748), .B1(n_674), .B2(n_681), .Y(n_784) );
OR2x6_ASAP7_75t_L g785 ( .A(n_743), .B(n_663), .Y(n_785) );
HB1xp67_ASAP7_75t_SL g786 ( .A(n_697), .Y(n_786) );
OAI221xp5_ASAP7_75t_L g787 ( .A1(n_725), .A2(n_723), .B1(n_732), .B2(n_701), .C(n_695), .Y(n_787) );
AND2x2_ASAP7_75t_L g788 ( .A(n_738), .B(n_750), .Y(n_788) );
INVx2_ASAP7_75t_L g789 ( .A(n_662), .Y(n_789) );
AND2x4_ASAP7_75t_L g790 ( .A(n_741), .B(n_756), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_709), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_712), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_664), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_653), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_728), .B(n_685), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_656), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_739), .Y(n_797) );
AOI22xp5_ASAP7_75t_L g798 ( .A1(n_659), .A2(n_655), .B1(n_686), .B2(n_657), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_679), .B(n_691), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_745), .Y(n_800) );
INVx1_ASAP7_75t_SL g801 ( .A(n_741), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_661), .B(n_733), .Y(n_802) );
AO22x2_ASAP7_75t_L g803 ( .A1(n_693), .A2(n_752), .B1(n_762), .B2(n_735), .Y(n_803) );
AND2x4_ASAP7_75t_L g804 ( .A(n_756), .B(n_737), .Y(n_804) );
A2O1A1Ixp33_ASAP7_75t_L g805 ( .A1(n_667), .A2(n_704), .B(n_658), .C(n_687), .Y(n_805) );
OR2x6_ASAP7_75t_L g806 ( .A(n_693), .B(n_737), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_697), .A2(n_733), .B1(n_669), .B2(n_708), .Y(n_807) );
AND2x2_ASAP7_75t_L g808 ( .A(n_707), .B(n_665), .Y(n_808) );
OA21x2_ASAP7_75t_L g809 ( .A1(n_722), .A2(n_666), .B(n_700), .Y(n_809) );
OA21x2_ASAP7_75t_L g810 ( .A1(n_696), .A2(n_699), .B(n_710), .Y(n_810) );
OA21x2_ASAP7_75t_L g811 ( .A1(n_761), .A2(n_765), .B(n_736), .Y(n_811) );
OAI21xp5_ASAP7_75t_L g812 ( .A1(n_694), .A2(n_672), .B(n_683), .Y(n_812) );
AO21x2_ASAP7_75t_L g813 ( .A1(n_718), .A2(n_765), .B(n_761), .Y(n_813) );
AND2x2_ASAP7_75t_SL g814 ( .A(n_730), .B(n_711), .Y(n_814) );
INVx4_ASAP7_75t_L g815 ( .A(n_749), .Y(n_815) );
AOI21xp5_ASAP7_75t_L g816 ( .A1(n_731), .A2(n_727), .B(n_689), .Y(n_816) );
AOI22xp33_ASAP7_75t_SL g817 ( .A1(n_665), .A2(n_727), .B1(n_719), .B2(n_721), .Y(n_817) );
INVx2_ASAP7_75t_L g818 ( .A(n_665), .Y(n_818) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_721), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_727), .A2(n_763), .B1(n_758), .B2(n_614), .Y(n_820) );
AOI21xp5_ASAP7_75t_L g821 ( .A1(n_689), .A2(n_764), .B(n_760), .Y(n_821) );
AOI21xp5_ASAP7_75t_L g822 ( .A1(n_706), .A2(n_764), .B(n_760), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_678), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_678), .Y(n_824) );
OR2x2_ASAP7_75t_L g825 ( .A(n_740), .B(n_444), .Y(n_825) );
A2O1A1Ixp33_ASAP7_75t_L g826 ( .A1(n_744), .A2(n_760), .B(n_764), .C(n_641), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_678), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_678), .Y(n_828) );
OAI21xp33_ASAP7_75t_L g829 ( .A1(n_760), .A2(n_764), .B(n_724), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_678), .Y(n_830) );
CKINVDCx6p67_ASAP7_75t_R g831 ( .A(n_673), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_678), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_678), .Y(n_833) );
INVx2_ASAP7_75t_L g834 ( .A(n_678), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_678), .Y(n_835) );
CKINVDCx12_ASAP7_75t_R g836 ( .A(n_673), .Y(n_836) );
BUFx12f_ASAP7_75t_L g837 ( .A(n_673), .Y(n_837) );
INVx2_ASAP7_75t_L g838 ( .A(n_678), .Y(n_838) );
INVx2_ASAP7_75t_L g839 ( .A(n_678), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_714), .B(n_720), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_763), .A2(n_758), .B1(n_614), .B2(n_724), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_763), .A2(n_758), .B1(n_614), .B2(n_724), .Y(n_842) );
AND2x4_ASAP7_75t_L g843 ( .A(n_743), .B(n_668), .Y(n_843) );
AO31x2_ASAP7_75t_L g844 ( .A1(n_760), .A2(n_764), .A3(n_717), .B(n_670), .Y(n_844) );
AOI22xp5_ASAP7_75t_L g845 ( .A1(n_763), .A2(n_754), .B1(n_758), .B2(n_573), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_678), .Y(n_846) );
INVx2_ASAP7_75t_SL g847 ( .A(n_742), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_678), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_714), .B(n_720), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_678), .Y(n_850) );
INVx4_ASAP7_75t_SL g851 ( .A(n_806), .Y(n_851) );
AND2x2_ASAP7_75t_L g852 ( .A(n_829), .B(n_845), .Y(n_852) );
BUFx2_ASAP7_75t_L g853 ( .A(n_803), .Y(n_853) );
AND2x2_ASAP7_75t_L g854 ( .A(n_829), .B(n_845), .Y(n_854) );
NOR2x1_ASAP7_75t_L g855 ( .A(n_806), .B(n_785), .Y(n_855) );
A2O1A1Ixp33_ASAP7_75t_L g856 ( .A1(n_778), .A2(n_784), .B(n_798), .C(n_826), .Y(n_856) );
OR2x6_ASAP7_75t_L g857 ( .A(n_806), .B(n_803), .Y(n_857) );
AO21x2_ASAP7_75t_L g858 ( .A1(n_821), .A2(n_822), .B(n_816), .Y(n_858) );
OR2x6_ASAP7_75t_L g859 ( .A(n_770), .B(n_785), .Y(n_859) );
INVx2_ASAP7_75t_L g860 ( .A(n_811), .Y(n_860) );
AND2x2_ASAP7_75t_L g861 ( .A(n_767), .B(n_789), .Y(n_861) );
AND2x2_ASAP7_75t_L g862 ( .A(n_799), .B(n_766), .Y(n_862) );
OAI22xp33_ASAP7_75t_L g863 ( .A1(n_798), .A2(n_784), .B1(n_769), .B2(n_825), .Y(n_863) );
HB1xp67_ASAP7_75t_L g864 ( .A(n_788), .Y(n_864) );
AND2x2_ASAP7_75t_L g865 ( .A(n_799), .B(n_827), .Y(n_865) );
OR2x6_ASAP7_75t_L g866 ( .A(n_785), .B(n_812), .Y(n_866) );
NOR2xp33_ASAP7_75t_L g867 ( .A(n_778), .B(n_787), .Y(n_867) );
BUFx2_ASAP7_75t_L g868 ( .A(n_773), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_820), .A2(n_841), .B1(n_842), .B2(n_769), .Y(n_869) );
INVxp67_ASAP7_75t_SL g870 ( .A(n_779), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_818), .Y(n_871) );
BUFx2_ASAP7_75t_L g872 ( .A(n_774), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_771), .B(n_840), .Y(n_873) );
OAI22xp5_ASAP7_75t_L g874 ( .A1(n_807), .A2(n_801), .B1(n_771), .B2(n_849), .Y(n_874) );
AND2x4_ASAP7_75t_SL g875 ( .A(n_804), .B(n_790), .Y(n_875) );
INVx4_ASAP7_75t_L g876 ( .A(n_804), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_840), .B(n_849), .Y(n_877) );
AND2x2_ASAP7_75t_L g878 ( .A(n_834), .B(n_838), .Y(n_878) );
NAND3xp33_ASAP7_75t_L g879 ( .A(n_817), .B(n_805), .C(n_812), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_779), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_823), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_824), .Y(n_882) );
AO21x2_ASAP7_75t_L g883 ( .A1(n_813), .A2(n_808), .B(n_802), .Y(n_883) );
INVx2_ASAP7_75t_L g884 ( .A(n_839), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_828), .Y(n_885) );
OR2x2_ASAP7_75t_L g886 ( .A(n_802), .B(n_783), .Y(n_886) );
OAI21xp5_ASAP7_75t_L g887 ( .A1(n_793), .A2(n_794), .B(n_795), .Y(n_887) );
BUFx2_ASAP7_75t_L g888 ( .A(n_774), .Y(n_888) );
AND2x2_ASAP7_75t_L g889 ( .A(n_830), .B(n_850), .Y(n_889) );
INVx2_ASAP7_75t_L g890 ( .A(n_791), .Y(n_890) );
INVx2_ASAP7_75t_SL g891 ( .A(n_814), .Y(n_891) );
OA21x2_ASAP7_75t_L g892 ( .A1(n_792), .A2(n_848), .B(n_846), .Y(n_892) );
AO21x2_ASAP7_75t_L g893 ( .A1(n_832), .A2(n_833), .B(n_835), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_844), .Y(n_894) );
OA21x2_ASAP7_75t_L g895 ( .A1(n_819), .A2(n_844), .B(n_780), .Y(n_895) );
AOI222xp33_ASAP7_75t_L g896 ( .A1(n_837), .A2(n_815), .B1(n_797), .B2(n_800), .C1(n_796), .C2(n_847), .Y(n_896) );
AOI22xp5_ASAP7_75t_L g897 ( .A1(n_781), .A2(n_843), .B1(n_836), .B2(n_786), .Y(n_897) );
AO21x2_ASAP7_75t_L g898 ( .A1(n_777), .A2(n_772), .B(n_775), .Y(n_898) );
AO21x2_ASAP7_75t_L g899 ( .A1(n_772), .A2(n_775), .B(n_782), .Y(n_899) );
INVx3_ASAP7_75t_L g900 ( .A(n_775), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_772), .Y(n_901) );
AND2x2_ASAP7_75t_L g902 ( .A(n_782), .B(n_810), .Y(n_902) );
AO21x2_ASAP7_75t_L g903 ( .A1(n_782), .A2(n_809), .B(n_776), .Y(n_903) );
AND2x2_ASAP7_75t_L g904 ( .A(n_809), .B(n_831), .Y(n_904) );
INVxp67_ASAP7_75t_SL g905 ( .A(n_815), .Y(n_905) );
OR2x6_ASAP7_75t_L g906 ( .A(n_806), .B(n_803), .Y(n_906) );
HB1xp67_ASAP7_75t_L g907 ( .A(n_768), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_871), .Y(n_908) );
AND2x2_ASAP7_75t_L g909 ( .A(n_852), .B(n_854), .Y(n_909) );
AND2x2_ASAP7_75t_L g910 ( .A(n_862), .B(n_865), .Y(n_910) );
INVx2_ASAP7_75t_SL g911 ( .A(n_875), .Y(n_911) );
AND2x4_ASAP7_75t_SL g912 ( .A(n_876), .B(n_857), .Y(n_912) );
AND2x2_ASAP7_75t_L g913 ( .A(n_862), .B(n_865), .Y(n_913) );
INVx2_ASAP7_75t_L g914 ( .A(n_860), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_880), .B(n_870), .Y(n_915) );
AND2x2_ASAP7_75t_L g916 ( .A(n_861), .B(n_903), .Y(n_916) );
OAI31xp33_ASAP7_75t_L g917 ( .A1(n_863), .A2(n_856), .A3(n_874), .B(n_867), .Y(n_917) );
AND2x2_ASAP7_75t_L g918 ( .A(n_903), .B(n_890), .Y(n_918) );
AND2x2_ASAP7_75t_L g919 ( .A(n_890), .B(n_878), .Y(n_919) );
HB1xp67_ASAP7_75t_L g920 ( .A(n_864), .Y(n_920) );
BUFx2_ASAP7_75t_L g921 ( .A(n_857), .Y(n_921) );
AND2x2_ASAP7_75t_L g922 ( .A(n_878), .B(n_889), .Y(n_922) );
AND2x2_ASAP7_75t_SL g923 ( .A(n_853), .B(n_875), .Y(n_923) );
AND2x2_ASAP7_75t_L g924 ( .A(n_904), .B(n_884), .Y(n_924) );
INVx5_ASAP7_75t_SL g925 ( .A(n_857), .Y(n_925) );
INVx5_ASAP7_75t_L g926 ( .A(n_857), .Y(n_926) );
OR2x6_ASAP7_75t_L g927 ( .A(n_906), .B(n_866), .Y(n_927) );
NAND4xp25_ASAP7_75t_L g928 ( .A(n_869), .B(n_896), .C(n_879), .D(n_887), .Y(n_928) );
INVxp67_ASAP7_75t_SL g929 ( .A(n_873), .Y(n_929) );
AND2x2_ASAP7_75t_L g930 ( .A(n_881), .B(n_882), .Y(n_930) );
AND2x2_ASAP7_75t_L g931 ( .A(n_882), .B(n_885), .Y(n_931) );
OR2x2_ASAP7_75t_L g932 ( .A(n_886), .B(n_877), .Y(n_932) );
HB1xp67_ASAP7_75t_L g933 ( .A(n_907), .Y(n_933) );
AND2x2_ASAP7_75t_L g934 ( .A(n_894), .B(n_902), .Y(n_934) );
AND2x4_ASAP7_75t_L g935 ( .A(n_851), .B(n_859), .Y(n_935) );
AND2x2_ASAP7_75t_L g936 ( .A(n_902), .B(n_892), .Y(n_936) );
AND2x2_ASAP7_75t_L g937 ( .A(n_892), .B(n_893), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_892), .Y(n_938) );
AND2x2_ASAP7_75t_L g939 ( .A(n_892), .B(n_893), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_893), .B(n_886), .Y(n_940) );
AND2x4_ASAP7_75t_L g941 ( .A(n_851), .B(n_859), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_908), .Y(n_942) );
AND2x2_ASAP7_75t_L g943 ( .A(n_936), .B(n_900), .Y(n_943) );
AND2x2_ASAP7_75t_L g944 ( .A(n_936), .B(n_900), .Y(n_944) );
AND2x2_ASAP7_75t_L g945 ( .A(n_909), .B(n_899), .Y(n_945) );
AND2x2_ASAP7_75t_L g946 ( .A(n_934), .B(n_899), .Y(n_946) );
NAND3xp33_ASAP7_75t_L g947 ( .A(n_928), .B(n_906), .C(n_897), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g948 ( .A(n_929), .B(n_883), .Y(n_948) );
OR2x2_ASAP7_75t_L g949 ( .A(n_940), .B(n_901), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_934), .B(n_899), .Y(n_950) );
AND2x4_ASAP7_75t_L g951 ( .A(n_935), .B(n_906), .Y(n_951) );
AND2x2_ASAP7_75t_L g952 ( .A(n_916), .B(n_901), .Y(n_952) );
AND2x2_ASAP7_75t_L g953 ( .A(n_916), .B(n_895), .Y(n_953) );
INVx2_ASAP7_75t_L g954 ( .A(n_914), .Y(n_954) );
INVxp67_ASAP7_75t_L g955 ( .A(n_920), .Y(n_955) );
AND2x2_ASAP7_75t_L g956 ( .A(n_937), .B(n_898), .Y(n_956) );
AND2x2_ASAP7_75t_SL g957 ( .A(n_923), .B(n_876), .Y(n_957) );
OR2x2_ASAP7_75t_L g958 ( .A(n_910), .B(n_866), .Y(n_958) );
AND2x2_ASAP7_75t_L g959 ( .A(n_937), .B(n_939), .Y(n_959) );
OR2x2_ASAP7_75t_L g960 ( .A(n_910), .B(n_866), .Y(n_960) );
AND2x2_ASAP7_75t_L g961 ( .A(n_924), .B(n_913), .Y(n_961) );
OR2x2_ASAP7_75t_L g962 ( .A(n_913), .B(n_866), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_922), .B(n_918), .Y(n_963) );
INVx1_ASAP7_75t_SL g964 ( .A(n_933), .Y(n_964) );
OR2x2_ASAP7_75t_L g965 ( .A(n_915), .B(n_858), .Y(n_965) );
OR2x2_ASAP7_75t_L g966 ( .A(n_915), .B(n_858), .Y(n_966) );
AND2x2_ASAP7_75t_L g967 ( .A(n_959), .B(n_927), .Y(n_967) );
AND2x2_ASAP7_75t_L g968 ( .A(n_959), .B(n_943), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_961), .B(n_919), .Y(n_969) );
AND2x2_ASAP7_75t_L g970 ( .A(n_943), .B(n_944), .Y(n_970) );
INVx2_ASAP7_75t_SL g971 ( .A(n_957), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_961), .B(n_919), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_942), .Y(n_973) );
INVx1_ASAP7_75t_L g974 ( .A(n_942), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_964), .B(n_930), .Y(n_975) );
INVx2_ASAP7_75t_L g976 ( .A(n_954), .Y(n_976) );
NAND2xp5_ASAP7_75t_SL g977 ( .A(n_947), .B(n_923), .Y(n_977) );
INVx1_ASAP7_75t_SL g978 ( .A(n_964), .Y(n_978) );
OR2x2_ASAP7_75t_L g979 ( .A(n_963), .B(n_932), .Y(n_979) );
OR2x2_ASAP7_75t_L g980 ( .A(n_963), .B(n_921), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_955), .B(n_930), .Y(n_981) );
NAND2x1p5_ASAP7_75t_L g982 ( .A(n_957), .B(n_855), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_955), .B(n_931), .Y(n_983) );
INVxp67_ASAP7_75t_L g984 ( .A(n_949), .Y(n_984) );
AND2x4_ASAP7_75t_L g985 ( .A(n_951), .B(n_926), .Y(n_985) );
AND2x2_ASAP7_75t_L g986 ( .A(n_945), .B(n_938), .Y(n_986) );
NAND2xp5_ASAP7_75t_SL g987 ( .A(n_977), .B(n_923), .Y(n_987) );
OR2x2_ASAP7_75t_L g988 ( .A(n_979), .B(n_948), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_975), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_984), .B(n_946), .Y(n_990) );
NOR2xp33_ASAP7_75t_L g991 ( .A(n_978), .B(n_928), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_973), .Y(n_992) );
OR2x2_ASAP7_75t_L g993 ( .A(n_969), .B(n_952), .Y(n_993) );
AND2x2_ASAP7_75t_L g994 ( .A(n_968), .B(n_953), .Y(n_994) );
INVxp67_ASAP7_75t_L g995 ( .A(n_981), .Y(n_995) );
AND2x2_ASAP7_75t_L g996 ( .A(n_968), .B(n_953), .Y(n_996) );
OR2x2_ASAP7_75t_L g997 ( .A(n_972), .B(n_952), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_974), .Y(n_998) );
INVx2_ASAP7_75t_L g999 ( .A(n_976), .Y(n_999) );
AND2x2_ASAP7_75t_L g1000 ( .A(n_970), .B(n_953), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g1001 ( .A(n_986), .B(n_950), .Y(n_1001) );
INVx1_ASAP7_75t_L g1002 ( .A(n_983), .Y(n_1002) );
NAND2xp5_ASAP7_75t_L g1003 ( .A(n_986), .B(n_950), .Y(n_1003) );
NAND2xp5_ASAP7_75t_SL g1004 ( .A(n_971), .B(n_926), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_992), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_994), .B(n_970), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_998), .Y(n_1007) );
OAI21xp5_ASAP7_75t_SL g1008 ( .A1(n_987), .A2(n_982), .B(n_917), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_989), .B(n_956), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_1002), .B(n_956), .Y(n_1010) );
INVx1_ASAP7_75t_L g1011 ( .A(n_999), .Y(n_1011) );
OAI322xp33_ASAP7_75t_L g1012 ( .A1(n_991), .A2(n_995), .A3(n_988), .B1(n_987), .B2(n_990), .C1(n_993), .C2(n_997), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_988), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_1013), .Y(n_1014) );
OAI211xp5_ASAP7_75t_L g1015 ( .A1(n_1008), .A2(n_991), .B(n_905), .C(n_917), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g1016 ( .A(n_1006), .B(n_994), .Y(n_1016) );
AOI221xp5_ASAP7_75t_L g1017 ( .A1(n_1012), .A2(n_1000), .B1(n_996), .B2(n_1003), .C(n_1001), .Y(n_1017) );
NAND4xp75_ASAP7_75t_L g1018 ( .A(n_1010), .B(n_855), .C(n_1004), .D(n_891), .Y(n_1018) );
AOI221xp5_ASAP7_75t_L g1019 ( .A1(n_1015), .A2(n_1005), .B1(n_1007), .B2(n_1009), .C(n_1011), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_1016), .B(n_967), .Y(n_1020) );
OAI211xp5_ASAP7_75t_L g1021 ( .A1(n_1017), .A2(n_891), .B(n_926), .C(n_911), .Y(n_1021) );
NOR3xp33_ASAP7_75t_L g1022 ( .A(n_1021), .B(n_1018), .C(n_1014), .Y(n_1022) );
NAND3xp33_ASAP7_75t_SL g1023 ( .A(n_1019), .B(n_980), .C(n_958), .Y(n_1023) );
OR2x2_ASAP7_75t_L g1024 ( .A(n_1023), .B(n_1020), .Y(n_1024) );
NAND3xp33_ASAP7_75t_L g1025 ( .A(n_1022), .B(n_859), .C(n_966), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_1024), .Y(n_1026) );
NOR3x2_ASAP7_75t_L g1027 ( .A(n_1025), .B(n_960), .C(n_962), .Y(n_1027) );
OAI22xp5_ASAP7_75t_SL g1028 ( .A1(n_1026), .A2(n_951), .B1(n_941), .B2(n_935), .Y(n_1028) );
XNOR2xp5_ASAP7_75t_L g1029 ( .A(n_1028), .B(n_1027), .Y(n_1029) );
OAI22xp5_ASAP7_75t_L g1030 ( .A1(n_1029), .A2(n_925), .B1(n_966), .B2(n_965), .Y(n_1030) );
OA21x2_ASAP7_75t_L g1031 ( .A1(n_1030), .A2(n_941), .B(n_985), .Y(n_1031) );
AOI22x1_ASAP7_75t_L g1032 ( .A1(n_1031), .A2(n_872), .B1(n_868), .B2(n_888), .Y(n_1032) );
AOI22xp33_ASAP7_75t_SL g1033 ( .A1(n_1032), .A2(n_912), .B1(n_925), .B2(n_985), .Y(n_1033) );
endmodule