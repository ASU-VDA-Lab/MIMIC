module fake_netlist_5_1778_n_1701 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1701);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1701;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_314;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1543;
wire n_1399;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_48),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_154),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_42),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_79),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_51),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_64),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_68),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_136),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_20),
.Y(n_165)
);

INVxp67_ASAP7_75t_SL g166 ( 
.A(n_70),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_126),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_47),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_48),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_145),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_26),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_21),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_11),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_38),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_86),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_38),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_115),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_42),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_98),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_29),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_83),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_71),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_144),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_53),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_97),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_128),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_10),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_18),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_11),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_112),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_99),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_84),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_1),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_65),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_27),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_139),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_119),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_141),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_49),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_3),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_56),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_150),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_61),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_6),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_3),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_73),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_85),
.Y(n_209)
);

BUFx10_ASAP7_75t_L g210 ( 
.A(n_58),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_63),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_26),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_32),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_140),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_138),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_49),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_153),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_35),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_15),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_89),
.Y(n_220)
);

INVxp67_ASAP7_75t_SL g221 ( 
.A(n_37),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_29),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_34),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_10),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_18),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_23),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_54),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_78),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_67),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_146),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_93),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_15),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_47),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_13),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_132),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_142),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_9),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_147),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_111),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_69),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_94),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_51),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_17),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_152),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_129),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_116),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_53),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_0),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_44),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_103),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_34),
.Y(n_251)
);

INVxp67_ASAP7_75t_SL g252 ( 
.A(n_88),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_105),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_123),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_2),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_6),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_37),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_151),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_95),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_27),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_133),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_82),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_87),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_76),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_57),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_16),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_148),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_14),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_56),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_75),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_7),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_7),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_104),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_40),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_16),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_40),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_25),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_135),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_114),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_33),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_19),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_20),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_77),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_106),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_81),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_50),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_66),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_54),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_22),
.Y(n_289)
);

BUFx10_ASAP7_75t_L g290 ( 
.A(n_137),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_59),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_13),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_1),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_12),
.Y(n_294)
);

BUFx5_ASAP7_75t_L g295 ( 
.A(n_0),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_131),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_30),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_149),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_80),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_8),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_46),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_28),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_25),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_22),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_30),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_110),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_43),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_31),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_127),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_5),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_233),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_295),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_273),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_160),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_158),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_295),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_295),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_2),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_163),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_295),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_162),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_295),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_196),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_295),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_164),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_199),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_183),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_295),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_295),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_167),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_205),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_211),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_248),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_171),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_246),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_183),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_248),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_177),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_229),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_179),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_181),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_184),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_248),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_258),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_213),
.B(n_4),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_248),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_263),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_287),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_248),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_248),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_195),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_287),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_195),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_185),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_233),
.Y(n_355)
);

NOR2xp67_ASAP7_75t_L g356 ( 
.A(n_201),
.B(n_4),
.Y(n_356)
);

INVx2_ASAP7_75t_SL g357 ( 
.A(n_222),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_303),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_298),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_229),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_187),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_172),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_172),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_190),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_188),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_190),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_193),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_197),
.Y(n_368)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_298),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_194),
.B(n_5),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_210),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_197),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_198),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_200),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_303),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_202),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_208),
.Y(n_377)
);

INVxp33_ASAP7_75t_SL g378 ( 
.A(n_225),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_209),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_214),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_228),
.Y(n_381)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_369),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_324),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_333),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_324),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_324),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_369),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_356),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_359),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_333),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_327),
.B(n_222),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_336),
.B(n_339),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_337),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_359),
.Y(n_394)
);

NAND2xp33_ASAP7_75t_L g395 ( 
.A(n_318),
.B(n_201),
.Y(n_395)
);

OA21x2_ASAP7_75t_L g396 ( 
.A1(n_318),
.A2(n_212),
.B(n_202),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_337),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_360),
.B(n_370),
.Y(n_398)
);

CKINVDCx8_ASAP7_75t_R g399 ( 
.A(n_371),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_359),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_312),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_356),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_343),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_343),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_315),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_346),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_346),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_357),
.B(n_276),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_348),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_349),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_378),
.B(n_194),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_369),
.B(n_215),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_352),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_369),
.Y(n_414)
);

INVx6_ASAP7_75t_L g415 ( 
.A(n_371),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_349),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_312),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_350),
.B(n_215),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_316),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_316),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_345),
.B(n_278),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_357),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_317),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_350),
.B(n_230),
.Y(n_424)
);

AND3x2_ASAP7_75t_L g425 ( 
.A(n_358),
.B(n_286),
.C(n_169),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_317),
.B(n_235),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_320),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_320),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_322),
.B(n_276),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_322),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_328),
.Y(n_431)
);

OAI21x1_ASAP7_75t_L g432 ( 
.A1(n_328),
.A2(n_169),
.B(n_157),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_329),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_329),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_311),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_351),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_351),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_353),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_353),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_313),
.B(n_261),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_362),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_362),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_363),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_363),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_364),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_364),
.B(n_366),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_392),
.B(n_321),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_427),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_440),
.B(n_325),
.Y(n_449)
);

INVx5_ASAP7_75t_L g450 ( 
.A(n_417),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_421),
.A2(n_358),
.B1(n_375),
.B2(n_355),
.Y(n_451)
);

AND3x2_ASAP7_75t_L g452 ( 
.A(n_411),
.B(n_375),
.C(n_221),
.Y(n_452)
);

NOR3xp33_ASAP7_75t_L g453 ( 
.A(n_411),
.B(n_421),
.C(n_440),
.Y(n_453)
);

OR2x6_ASAP7_75t_L g454 ( 
.A(n_415),
.B(n_260),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_L g455 ( 
.A1(n_395),
.A2(n_260),
.B1(n_266),
.B2(n_294),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_422),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_385),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_405),
.B(n_330),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_422),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_392),
.B(n_334),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_427),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g462 ( 
.A(n_409),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_409),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_427),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_398),
.B(n_338),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_392),
.A2(n_354),
.B1(n_365),
.B2(n_379),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_395),
.A2(n_266),
.B1(n_294),
.B2(n_307),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_388),
.B(n_340),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_431),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_383),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_385),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_385),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_385),
.Y(n_473)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_383),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_386),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_429),
.B(n_157),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_386),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_431),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_435),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_388),
.B(n_341),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_386),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_398),
.B(n_342),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_386),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_431),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_417),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_433),
.Y(n_486)
);

INVxp33_ASAP7_75t_L g487 ( 
.A(n_435),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_409),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_L g489 ( 
.A1(n_396),
.A2(n_307),
.B1(n_219),
.B2(n_223),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_433),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_401),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_383),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_433),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_401),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_401),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_417),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_402),
.B(n_361),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_402),
.B(n_367),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_426),
.B(n_373),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_434),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_434),
.Y(n_501)
);

AND2x6_ASAP7_75t_L g502 ( 
.A(n_412),
.B(n_298),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_434),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_401),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_423),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_399),
.B(n_374),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_396),
.A2(n_251),
.B1(n_216),
.B2(n_218),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_426),
.B(n_377),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_419),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_419),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_423),
.Y(n_511)
);

INVx5_ASAP7_75t_L g512 ( 
.A(n_417),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_415),
.A2(n_380),
.B1(n_381),
.B2(n_347),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_383),
.Y(n_514)
);

OR2x6_ASAP7_75t_L g515 ( 
.A(n_415),
.B(n_212),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_424),
.B(n_238),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_419),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_399),
.B(n_210),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_424),
.B(n_239),
.Y(n_519)
);

INVx5_ASAP7_75t_L g520 ( 
.A(n_417),
.Y(n_520)
);

BUFx4f_ASAP7_75t_L g521 ( 
.A(n_396),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_423),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_423),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_423),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_408),
.B(n_186),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_423),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_419),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_415),
.A2(n_314),
.B1(n_344),
.B2(n_335),
.Y(n_528)
);

NOR3xp33_ASAP7_75t_L g529 ( 
.A(n_413),
.B(n_161),
.C(n_156),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_428),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_399),
.B(n_210),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_428),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_428),
.Y(n_533)
);

OAI22xp33_ASAP7_75t_L g534 ( 
.A1(n_415),
.A2(n_399),
.B1(n_207),
.B2(n_206),
.Y(n_534)
);

INVx1_ASAP7_75t_SL g535 ( 
.A(n_413),
.Y(n_535)
);

NAND3xp33_ASAP7_75t_SL g536 ( 
.A(n_413),
.B(n_170),
.C(n_159),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_391),
.B(n_319),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_396),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_383),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_428),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_429),
.B(n_366),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_391),
.B(n_210),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_391),
.B(n_323),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_429),
.B(n_173),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_382),
.B(n_241),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_382),
.B(n_244),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_432),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_383),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_396),
.Y(n_549)
);

INVxp67_ASAP7_75t_SL g550 ( 
.A(n_383),
.Y(n_550)
);

NAND2xp33_ASAP7_75t_SL g551 ( 
.A(n_408),
.B(n_174),
.Y(n_551)
);

INVxp67_ASAP7_75t_SL g552 ( 
.A(n_383),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_382),
.B(n_245),
.Y(n_553)
);

BUFx10_ASAP7_75t_L g554 ( 
.A(n_415),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_432),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_383),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_432),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_384),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_408),
.B(n_326),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_432),
.Y(n_560)
);

BUFx10_ASAP7_75t_L g561 ( 
.A(n_415),
.Y(n_561)
);

AND2x6_ASAP7_75t_L g562 ( 
.A(n_412),
.B(n_298),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_412),
.B(n_259),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_443),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_382),
.B(n_250),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_443),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_382),
.B(n_253),
.Y(n_567)
);

NAND2xp33_ASAP7_75t_R g568 ( 
.A(n_396),
.B(n_165),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_382),
.B(n_331),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_412),
.A2(n_247),
.B1(n_216),
.B2(n_308),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_412),
.A2(n_247),
.B1(n_218),
.B2(n_308),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_443),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_412),
.A2(n_249),
.B1(n_219),
.B2(n_304),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_384),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_437),
.B(n_332),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_437),
.B(n_168),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_417),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_384),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_437),
.B(n_175),
.Y(n_579)
);

INVx8_ASAP7_75t_L g580 ( 
.A(n_417),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_390),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_390),
.Y(n_582)
);

OAI22xp33_ASAP7_75t_L g583 ( 
.A1(n_446),
.A2(n_234),
.B1(n_232),
.B2(n_227),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_417),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_425),
.Y(n_585)
);

OR2x6_ASAP7_75t_L g586 ( 
.A(n_446),
.B(n_223),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_390),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_417),
.B(n_254),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_393),
.Y(n_589)
);

INVx4_ASAP7_75t_L g590 ( 
.A(n_420),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_441),
.B(n_259),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_420),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_420),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_393),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_465),
.B(n_425),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_482),
.B(n_420),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_499),
.B(n_508),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_564),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_453),
.A2(n_252),
.B1(n_166),
.B2(n_270),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_516),
.B(n_420),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_568),
.A2(n_262),
.B1(n_284),
.B2(n_283),
.Y(n_601)
);

OAI22xp33_ASAP7_75t_L g602 ( 
.A1(n_447),
.A2(n_240),
.B1(n_236),
.B2(n_231),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_538),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_460),
.B(n_176),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_519),
.B(n_420),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_541),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_541),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_528),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_448),
.B(n_420),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_461),
.B(n_420),
.Y(n_610)
);

OAI221xp5_ASAP7_75t_L g611 ( 
.A1(n_570),
.A2(n_243),
.B1(n_249),
.B2(n_255),
.C(n_272),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_564),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_538),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_464),
.B(n_420),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_484),
.B(n_430),
.Y(n_615)
);

NOR3xp33_ASAP7_75t_SL g616 ( 
.A(n_536),
.B(n_180),
.C(n_178),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_456),
.B(n_182),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_486),
.B(n_430),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_456),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_513),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_549),
.Y(n_621)
);

AND2x6_ASAP7_75t_SL g622 ( 
.A(n_537),
.B(n_243),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_490),
.B(n_430),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_566),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_521),
.B(n_430),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_459),
.B(n_189),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_569),
.A2(n_291),
.B1(n_306),
.B2(n_299),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_493),
.B(n_430),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_500),
.B(n_501),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_497),
.B(n_265),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_503),
.B(n_430),
.Y(n_631)
);

NAND3xp33_ASAP7_75t_L g632 ( 
.A(n_451),
.B(n_242),
.C(n_203),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_566),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_572),
.B(n_430),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_459),
.B(n_498),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_521),
.B(n_430),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_572),
.B(n_430),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_469),
.B(n_441),
.Y(n_638)
);

NOR2xp67_ASAP7_75t_SL g639 ( 
.A(n_549),
.B(n_547),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_574),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_550),
.A2(n_418),
.B(n_414),
.Y(n_641)
);

NOR2xp67_ASAP7_75t_L g642 ( 
.A(n_466),
.B(n_418),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_498),
.B(n_267),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_543),
.B(n_368),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_469),
.B(n_441),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_478),
.B(n_441),
.Y(n_646)
);

O2A1O1Ixp33_ASAP7_75t_L g647 ( 
.A1(n_586),
.A2(n_272),
.B(n_251),
.C(n_304),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_478),
.B(n_441),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_505),
.B(n_441),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_558),
.Y(n_650)
);

BUFx8_ASAP7_75t_L g651 ( 
.A(n_479),
.Y(n_651)
);

NOR2x1p5_ASAP7_75t_L g652 ( 
.A(n_525),
.B(n_224),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_534),
.B(n_296),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_558),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_578),
.Y(n_655)
);

A2O1A1Ixp33_ASAP7_75t_L g656 ( 
.A1(n_521),
.A2(n_236),
.B(n_192),
.C(n_204),
.Y(n_656)
);

NOR2xp67_ASAP7_75t_L g657 ( 
.A(n_559),
.B(n_438),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_575),
.A2(n_231),
.B1(n_192),
.B2(n_204),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_578),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_525),
.B(n_259),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_574),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_581),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_507),
.B(n_298),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_551),
.A2(n_173),
.B1(n_309),
.B2(n_285),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_505),
.B(n_441),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_581),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_582),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_526),
.B(n_441),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_476),
.B(n_544),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_582),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_479),
.Y(n_671)
);

INVxp33_ASAP7_75t_L g672 ( 
.A(n_487),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_449),
.B(n_226),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_587),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_587),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_583),
.B(n_259),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_594),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_594),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_491),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_487),
.B(n_372),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_526),
.B(n_441),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_552),
.B(n_445),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_491),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_489),
.A2(n_255),
.B1(n_309),
.B2(n_264),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_554),
.B(n_298),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_452),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_589),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_476),
.B(n_544),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_511),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_542),
.B(n_237),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_L g691 ( 
.A1(n_515),
.A2(n_454),
.B1(n_544),
.B2(n_455),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_468),
.B(n_290),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_480),
.B(n_256),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_586),
.A2(n_557),
.B1(n_560),
.B2(n_555),
.Y(n_694)
);

INVxp67_ASAP7_75t_L g695 ( 
.A(n_551),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_522),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_523),
.B(n_445),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_518),
.B(n_531),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_524),
.B(n_445),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_576),
.B(n_445),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_547),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_585),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_579),
.B(n_445),
.Y(n_703)
);

NOR3xp33_ASAP7_75t_L g704 ( 
.A(n_462),
.B(n_300),
.C(n_257),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_554),
.B(n_445),
.Y(n_705)
);

INVxp67_ASAP7_75t_L g706 ( 
.A(n_463),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_585),
.B(n_458),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_548),
.B(n_445),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_548),
.B(n_445),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_494),
.Y(n_710)
);

NAND2xp33_ASAP7_75t_L g711 ( 
.A(n_502),
.B(n_217),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_494),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_470),
.B(n_445),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_554),
.B(n_387),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_506),
.B(n_268),
.Y(n_715)
);

OR2x6_ASAP7_75t_L g716 ( 
.A(n_586),
.B(n_217),
.Y(n_716)
);

AND2x4_ASAP7_75t_L g717 ( 
.A(n_586),
.B(n_372),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_561),
.B(n_290),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_555),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_470),
.B(n_387),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_563),
.B(n_269),
.Y(n_721)
);

NAND2xp33_ASAP7_75t_L g722 ( 
.A(n_502),
.B(n_220),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_561),
.B(n_290),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_470),
.B(n_387),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_557),
.Y(n_725)
);

AOI221xp5_ASAP7_75t_L g726 ( 
.A1(n_467),
.A2(n_191),
.B1(n_288),
.B2(n_310),
.C(n_302),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_515),
.B(n_271),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_560),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_492),
.B(n_387),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_492),
.B(n_387),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_492),
.B(n_387),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_514),
.B(n_414),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_561),
.B(n_290),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_515),
.B(n_274),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_571),
.B(n_220),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_495),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_485),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_514),
.B(n_414),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_514),
.B(n_414),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_485),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_495),
.Y(n_741)
);

INVx8_ASAP7_75t_L g742 ( 
.A(n_515),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_573),
.B(n_240),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_539),
.B(n_414),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_504),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_539),
.B(n_414),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_539),
.B(n_393),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_556),
.B(n_397),
.Y(n_748)
);

NAND2xp33_ASAP7_75t_L g749 ( 
.A(n_502),
.B(n_264),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_556),
.B(n_397),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_535),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_529),
.A2(n_285),
.B1(n_279),
.B2(n_444),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_556),
.B(n_397),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_545),
.B(n_275),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_592),
.B(n_403),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_454),
.A2(n_279),
.B1(n_442),
.B2(n_444),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_592),
.B(n_403),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_504),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_454),
.B(n_376),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_592),
.B(n_403),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_546),
.B(n_553),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_509),
.Y(n_762)
);

OAI22xp5_ASAP7_75t_SL g763 ( 
.A1(n_488),
.A2(n_305),
.B1(n_280),
.B2(n_281),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_509),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_588),
.B(n_436),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_597),
.B(n_565),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_644),
.B(n_567),
.Y(n_767)
);

AO21x2_ASAP7_75t_L g768 ( 
.A1(n_625),
.A2(n_591),
.B(n_527),
.Y(n_768)
);

BUFx4f_ASAP7_75t_L g769 ( 
.A(n_751),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_625),
.A2(n_580),
.B(n_474),
.Y(n_770)
);

A2O1A1Ixp33_ASAP7_75t_L g771 ( 
.A1(n_698),
.A2(n_577),
.B(n_540),
.C(n_533),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_672),
.B(n_488),
.Y(n_772)
);

OR2x6_ASAP7_75t_L g773 ( 
.A(n_742),
.B(n_454),
.Y(n_773)
);

NAND3xp33_ASAP7_75t_L g774 ( 
.A(n_726),
.B(n_277),
.C(n_282),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_604),
.B(n_577),
.Y(n_775)
);

A2O1A1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_698),
.A2(n_510),
.B(n_517),
.C(n_530),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_604),
.B(n_754),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_635),
.B(n_590),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_635),
.B(n_590),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_754),
.B(n_510),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_695),
.B(n_590),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_L g782 ( 
.A1(n_636),
.A2(n_517),
.B(n_530),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_657),
.B(n_532),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_606),
.B(n_532),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_636),
.A2(n_580),
.B(n_474),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_642),
.A2(n_502),
.B1(n_562),
.B2(n_593),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_705),
.A2(n_580),
.B(n_593),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_705),
.A2(n_580),
.B(n_593),
.Y(n_788)
);

NAND2x1_ASAP7_75t_L g789 ( 
.A(n_613),
.B(n_485),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_680),
.B(n_376),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_598),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_606),
.B(n_617),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_596),
.A2(n_682),
.B(n_605),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_671),
.B(n_289),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_595),
.A2(n_502),
.B1(n_562),
.B2(n_485),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_617),
.B(n_438),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_613),
.Y(n_797)
);

O2A1O1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_602),
.A2(n_481),
.B(n_477),
.C(n_475),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_613),
.Y(n_799)
);

OAI21xp5_ASAP7_75t_L g800 ( 
.A1(n_761),
.A2(n_472),
.B(n_471),
.Y(n_800)
);

OAI21xp5_ASAP7_75t_L g801 ( 
.A1(n_761),
.A2(n_472),
.B(n_471),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_600),
.A2(n_584),
.B(n_485),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_603),
.B(n_457),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_641),
.A2(n_703),
.B(n_700),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_714),
.A2(n_584),
.B(n_496),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_694),
.A2(n_688),
.B1(n_603),
.B2(n_684),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_595),
.A2(n_562),
.B1(n_502),
.B2(n_496),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_714),
.A2(n_685),
.B(n_765),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_624),
.Y(n_809)
);

NAND2x1p5_ASAP7_75t_L g810 ( 
.A(n_613),
.B(n_496),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_669),
.B(n_438),
.Y(n_811)
);

O2A1O1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_653),
.A2(n_473),
.B(n_483),
.C(n_481),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_707),
.B(n_496),
.Y(n_813)
);

AOI21x1_ASAP7_75t_L g814 ( 
.A1(n_765),
.A2(n_475),
.B(n_457),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_626),
.B(n_439),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_685),
.A2(n_584),
.B(n_496),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_720),
.A2(n_584),
.B(n_450),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_612),
.B(n_473),
.Y(n_818)
);

CKINVDCx8_ASAP7_75t_R g819 ( 
.A(n_622),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_707),
.B(n_292),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_724),
.A2(n_584),
.B(n_450),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_626),
.B(n_293),
.Y(n_822)
);

OAI21xp5_ASAP7_75t_L g823 ( 
.A1(n_634),
.A2(n_483),
.B(n_477),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_673),
.A2(n_439),
.B(n_444),
.C(n_442),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_669),
.A2(n_673),
.B1(n_691),
.B2(n_621),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_633),
.B(n_562),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_637),
.A2(n_562),
.B(n_520),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_640),
.B(n_562),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_661),
.Y(n_829)
);

OAI21xp33_ASAP7_75t_L g830 ( 
.A1(n_693),
.A2(n_297),
.B(n_301),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_674),
.B(n_442),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_729),
.A2(n_520),
.B(n_512),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_730),
.A2(n_732),
.B(n_731),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_738),
.A2(n_520),
.B(n_512),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_662),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_701),
.A2(n_520),
.B(n_512),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_619),
.B(n_607),
.Y(n_837)
);

OAI22xp5_ASAP7_75t_L g838 ( 
.A1(n_694),
.A2(n_410),
.B1(n_404),
.B2(n_406),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_677),
.B(n_442),
.Y(n_839)
);

O2A1O1Ixp5_ASAP7_75t_L g840 ( 
.A1(n_656),
.A2(n_410),
.B(n_407),
.C(n_404),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_662),
.Y(n_841)
);

OAI21xp33_ASAP7_75t_L g842 ( 
.A1(n_693),
.A2(n_439),
.B(n_407),
.Y(n_842)
);

OAI21xp5_ASAP7_75t_L g843 ( 
.A1(n_719),
.A2(n_520),
.B(n_512),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_678),
.B(n_407),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_666),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_687),
.B(n_406),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_739),
.A2(n_512),
.B(n_450),
.Y(n_847)
);

OAI21xp5_ASAP7_75t_L g848 ( 
.A1(n_725),
.A2(n_450),
.B(n_406),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_684),
.B(n_404),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_619),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_621),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_621),
.A2(n_416),
.B1(n_410),
.B2(n_436),
.Y(n_852)
);

O2A1O1Ixp5_ASAP7_75t_L g853 ( 
.A1(n_666),
.A2(n_416),
.B(n_400),
.C(n_394),
.Y(n_853)
);

A2O1A1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_715),
.A2(n_400),
.B(n_394),
.C(n_436),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_744),
.A2(n_746),
.B(n_740),
.Y(n_855)
);

INVxp67_ASAP7_75t_L g856 ( 
.A(n_759),
.Y(n_856)
);

NOR2xp67_ASAP7_75t_L g857 ( 
.A(n_601),
.B(n_72),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_629),
.B(n_436),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_717),
.B(n_436),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_667),
.Y(n_860)
);

OAI21xp5_ASAP7_75t_L g861 ( 
.A1(n_728),
.A2(n_450),
.B(n_400),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_621),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_667),
.B(n_436),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_670),
.B(n_436),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_717),
.B(n_436),
.Y(n_865)
);

AOI22xp5_ASAP7_75t_L g866 ( 
.A1(n_715),
.A2(n_436),
.B1(n_389),
.B2(n_394),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_740),
.A2(n_400),
.B(n_394),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_670),
.B(n_389),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_609),
.A2(n_389),
.B(n_155),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_675),
.B(n_389),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_599),
.A2(n_389),
.B1(n_143),
.B2(n_130),
.Y(n_871)
);

INVxp67_ASAP7_75t_L g872 ( 
.A(n_702),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_675),
.A2(n_389),
.B1(n_125),
.B2(n_124),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_650),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_740),
.A2(n_389),
.B(n_120),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_716),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_689),
.B(n_389),
.Y(n_877)
);

INVx3_ASAP7_75t_L g878 ( 
.A(n_737),
.Y(n_878)
);

OAI21xp33_ASAP7_75t_L g879 ( 
.A1(n_658),
.A2(n_389),
.B(n_9),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_740),
.A2(n_118),
.B(n_117),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_650),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_L g882 ( 
.A1(n_610),
.A2(n_113),
.B(n_109),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_652),
.B(n_8),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_696),
.B(n_12),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_716),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_654),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_654),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_690),
.B(n_14),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_713),
.A2(n_108),
.B(n_107),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_660),
.B(n_17),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_655),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_690),
.B(n_19),
.Y(n_892)
);

O2A1O1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_676),
.A2(n_21),
.B(n_23),
.C(n_24),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_655),
.B(n_24),
.Y(n_894)
);

O2A1O1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_647),
.A2(n_31),
.B(n_32),
.C(n_33),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_708),
.A2(n_102),
.B(n_101),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_L g897 ( 
.A1(n_663),
.A2(n_35),
.B1(n_36),
.B2(n_39),
.Y(n_897)
);

OAI321xp33_ASAP7_75t_L g898 ( 
.A1(n_664),
.A2(n_36),
.A3(n_39),
.B1(n_41),
.B2(n_43),
.C(n_44),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_709),
.A2(n_62),
.B(n_96),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_620),
.B(n_686),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_659),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_721),
.B(n_41),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_727),
.B(n_60),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_747),
.A2(n_74),
.B(n_92),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_742),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_679),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_721),
.A2(n_45),
.B(n_46),
.C(n_50),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_748),
.A2(n_90),
.B(n_91),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_750),
.A2(n_100),
.B(n_52),
.Y(n_909)
);

AOI22xp33_ASAP7_75t_L g910 ( 
.A1(n_663),
.A2(n_55),
.B1(n_45),
.B2(n_52),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_753),
.A2(n_55),
.B(n_618),
.Y(n_911)
);

OAI21xp33_ASAP7_75t_L g912 ( 
.A1(n_632),
.A2(n_643),
.B(n_704),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_614),
.A2(n_628),
.B(n_631),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_727),
.B(n_734),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_734),
.B(n_736),
.Y(n_915)
);

OR2x2_ASAP7_75t_L g916 ( 
.A(n_608),
.B(n_716),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_679),
.B(n_712),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_737),
.Y(n_918)
);

NAND3xp33_ASAP7_75t_L g919 ( 
.A(n_616),
.B(n_752),
.C(n_627),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_615),
.A2(n_623),
.B(n_755),
.Y(n_920)
);

NOR3xp33_ASAP7_75t_L g921 ( 
.A(n_763),
.B(n_692),
.C(n_630),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_683),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_718),
.B(n_723),
.Y(n_923)
);

NOR3xp33_ASAP7_75t_L g924 ( 
.A(n_611),
.B(n_735),
.C(n_743),
.Y(n_924)
);

OAI21xp5_ASAP7_75t_L g925 ( 
.A1(n_638),
.A2(n_645),
.B(n_646),
.Y(n_925)
);

OAI21xp5_ASAP7_75t_L g926 ( 
.A1(n_648),
.A2(n_760),
.B(n_757),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_683),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_710),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_649),
.A2(n_665),
.B(n_668),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_733),
.B(n_764),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_651),
.B(n_758),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_L g932 ( 
.A1(n_710),
.A2(n_762),
.B1(n_736),
.B2(n_712),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_762),
.B(n_745),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_741),
.B(n_681),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_651),
.B(n_756),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_742),
.B(n_697),
.Y(n_936)
);

OR2x6_ASAP7_75t_L g937 ( 
.A(n_699),
.B(n_639),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_711),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_722),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_749),
.B(n_644),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_625),
.A2(n_636),
.B(n_580),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_597),
.B(n_465),
.Y(n_942)
);

CKINVDCx20_ASAP7_75t_R g943 ( 
.A(n_651),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_625),
.A2(n_636),
.B(n_580),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_625),
.A2(n_636),
.B(n_580),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_597),
.B(n_465),
.Y(n_946)
);

OAI21xp33_ASAP7_75t_L g947 ( 
.A1(n_644),
.A2(n_453),
.B(n_411),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_793),
.A2(n_946),
.B(n_777),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_942),
.B(n_792),
.Y(n_949)
);

NAND2x1p5_ASAP7_75t_L g950 ( 
.A(n_862),
.B(n_905),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_769),
.Y(n_951)
);

INVxp33_ASAP7_75t_L g952 ( 
.A(n_772),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_825),
.A2(n_914),
.B1(n_767),
.B2(n_779),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_804),
.A2(n_766),
.B(n_775),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_943),
.Y(n_955)
);

NOR2x1p5_ASAP7_75t_L g956 ( 
.A(n_916),
.B(n_774),
.Y(n_956)
);

NAND2xp33_ASAP7_75t_SL g957 ( 
.A(n_905),
.B(n_888),
.Y(n_957)
);

AO21x1_ASAP7_75t_L g958 ( 
.A1(n_902),
.A2(n_903),
.B(n_822),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_791),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_769),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_808),
.A2(n_780),
.B(n_915),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_796),
.B(n_815),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_947),
.B(n_856),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_837),
.Y(n_964)
);

OAI21x1_ASAP7_75t_L g965 ( 
.A1(n_814),
.A2(n_855),
.B(n_802),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_922),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_829),
.Y(n_967)
);

OR2x2_ASAP7_75t_L g968 ( 
.A(n_856),
.B(n_900),
.Y(n_968)
);

INVx2_ASAP7_75t_SL g969 ( 
.A(n_883),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_905),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_905),
.B(n_850),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_850),
.B(n_811),
.Y(n_972)
);

AOI21x1_ASAP7_75t_L g973 ( 
.A1(n_941),
.A2(n_945),
.B(n_944),
.Y(n_973)
);

OAI21x1_ASAP7_75t_L g974 ( 
.A1(n_833),
.A2(n_805),
.B(n_782),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_822),
.A2(n_820),
.B1(n_921),
.B2(n_923),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_841),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_SL g977 ( 
.A1(n_923),
.A2(n_779),
.B(n_778),
.C(n_813),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_SL g978 ( 
.A(n_900),
.B(n_819),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_860),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_876),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_770),
.A2(n_785),
.B(n_787),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_778),
.B(n_790),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_922),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_806),
.A2(n_771),
.B(n_929),
.Y(n_984)
);

INVxp67_ASAP7_75t_L g985 ( 
.A(n_794),
.Y(n_985)
);

CKINVDCx10_ASAP7_75t_R g986 ( 
.A(n_773),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_912),
.B(n_830),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_813),
.A2(n_800),
.B(n_801),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_892),
.B(n_921),
.Y(n_989)
);

BUFx12f_ASAP7_75t_L g990 ( 
.A(n_773),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_876),
.B(n_885),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_885),
.B(n_890),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_931),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_809),
.Y(n_994)
);

NAND2x1p5_ASAP7_75t_L g995 ( 
.A(n_862),
.B(n_797),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_940),
.B(n_835),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_872),
.B(n_890),
.Y(n_997)
);

NAND2x1p5_ASAP7_75t_L g998 ( 
.A(n_862),
.B(n_797),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_926),
.A2(n_848),
.B(n_920),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_845),
.B(n_781),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_874),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_919),
.A2(n_930),
.B(n_924),
.C(n_879),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_781),
.B(n_784),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_773),
.Y(n_1004)
);

AO21x1_ASAP7_75t_L g1005 ( 
.A1(n_882),
.A2(n_869),
.B(n_871),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_934),
.B(n_886),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_935),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_811),
.B(n_872),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_799),
.Y(n_1009)
);

OR2x6_ASAP7_75t_SL g1010 ( 
.A(n_884),
.B(n_894),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_907),
.A2(n_893),
.B(n_898),
.C(n_895),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_799),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_901),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_851),
.Y(n_1014)
);

BUFx12f_ASAP7_75t_L g1015 ( 
.A(n_938),
.Y(n_1015)
);

OA22x2_ASAP7_75t_L g1016 ( 
.A1(n_795),
.A2(n_807),
.B1(n_936),
.B2(n_786),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_851),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_776),
.A2(n_913),
.B(n_803),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_924),
.A2(n_842),
.B(n_857),
.C(n_911),
.Y(n_1019)
);

O2A1O1Ixp5_ASAP7_75t_SL g1020 ( 
.A1(n_873),
.A2(n_838),
.B(n_928),
.C(n_927),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_788),
.A2(n_858),
.B(n_925),
.Y(n_1021)
);

BUFx12f_ASAP7_75t_L g1022 ( 
.A(n_938),
.Y(n_1022)
);

NOR3xp33_ASAP7_75t_L g1023 ( 
.A(n_859),
.B(n_865),
.C(n_909),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_881),
.Y(n_1024)
);

AOI21x1_ASAP7_75t_L g1025 ( 
.A1(n_863),
.A2(n_864),
.B(n_868),
.Y(n_1025)
);

O2A1O1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_846),
.A2(n_824),
.B(n_844),
.C(n_897),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_887),
.B(n_891),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_906),
.B(n_932),
.Y(n_1028)
);

OAI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_783),
.A2(n_939),
.B1(n_937),
.B2(n_810),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_789),
.A2(n_843),
.B(n_836),
.Y(n_1030)
);

AOI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_897),
.A2(n_910),
.B1(n_849),
.B2(n_938),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_861),
.A2(n_870),
.B(n_823),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_932),
.B(n_917),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_933),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_937),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_939),
.A2(n_937),
.B1(n_810),
.B2(n_938),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_831),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_877),
.A2(n_812),
.B(n_816),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_878),
.B(n_918),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_910),
.A2(n_854),
.B(n_818),
.C(n_839),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_878),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_918),
.B(n_828),
.Y(n_1042)
);

INVxp67_ASAP7_75t_L g1043 ( 
.A(n_826),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_798),
.A2(n_827),
.B(n_853),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_768),
.Y(n_1045)
);

INVx8_ASAP7_75t_L g1046 ( 
.A(n_852),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_853),
.Y(n_1047)
);

O2A1O1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_840),
.A2(n_908),
.B(n_904),
.C(n_889),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_866),
.A2(n_817),
.B1(n_821),
.B2(n_880),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_768),
.B(n_875),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_896),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_840),
.Y(n_1052)
);

NOR2x1_ASAP7_75t_R g1053 ( 
.A(n_899),
.B(n_867),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_832),
.A2(n_834),
.B(n_847),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_793),
.A2(n_946),
.B(n_804),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_777),
.A2(n_942),
.B(n_946),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_791),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_791),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_793),
.A2(n_946),
.B(n_804),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_942),
.B(n_946),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_791),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_942),
.B(n_946),
.Y(n_1062)
);

NOR3xp33_ASAP7_75t_SL g1063 ( 
.A(n_900),
.B(n_620),
.C(n_608),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_942),
.B(n_946),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_942),
.B(n_946),
.Y(n_1065)
);

OR2x6_ASAP7_75t_L g1066 ( 
.A(n_905),
.B(n_742),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_922),
.Y(n_1067)
);

O2A1O1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_777),
.A2(n_942),
.B(n_888),
.C(n_902),
.Y(n_1068)
);

OR2x2_ASAP7_75t_L g1069 ( 
.A(n_946),
.B(n_706),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_793),
.A2(n_946),
.B(n_777),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_850),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_793),
.A2(n_946),
.B(n_777),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_792),
.B(n_644),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_SL g1074 ( 
.A1(n_819),
.A2(n_620),
.B1(n_608),
.B2(n_488),
.Y(n_1074)
);

OR2x2_ASAP7_75t_L g1075 ( 
.A(n_946),
.B(n_706),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_791),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_777),
.A2(n_942),
.B(n_888),
.C(n_902),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_792),
.B(n_644),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_777),
.A2(n_942),
.B(n_946),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_793),
.A2(n_946),
.B(n_777),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_922),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_777),
.A2(n_942),
.B(n_888),
.C(n_902),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_942),
.B(n_946),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_791),
.Y(n_1084)
);

O2A1O1Ixp5_ASAP7_75t_L g1085 ( 
.A1(n_777),
.A2(n_942),
.B(n_888),
.C(n_946),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_905),
.Y(n_1086)
);

INVx1_ASAP7_75t_SL g1087 ( 
.A(n_837),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_793),
.A2(n_946),
.B(n_777),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_922),
.Y(n_1089)
);

AOI21xp33_ASAP7_75t_L g1090 ( 
.A1(n_975),
.A2(n_1077),
.B(n_1068),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_1017),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_965),
.A2(n_1054),
.B(n_973),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1001),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_981),
.A2(n_974),
.B(n_1038),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1055),
.A2(n_1059),
.B(n_948),
.Y(n_1095)
);

NOR2xp67_ASAP7_75t_L g1096 ( 
.A(n_987),
.B(n_1015),
.Y(n_1096)
);

BUFx3_ASAP7_75t_L g1097 ( 
.A(n_960),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_1017),
.Y(n_1098)
);

NOR2xp67_ASAP7_75t_SL g1099 ( 
.A(n_1022),
.B(n_1007),
.Y(n_1099)
);

OA21x2_ASAP7_75t_L g1100 ( 
.A1(n_984),
.A2(n_999),
.B(n_1044),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1013),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1065),
.A2(n_1060),
.B1(n_1064),
.B2(n_1083),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1038),
.A2(n_1018),
.B(n_1025),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_948),
.A2(n_1080),
.B(n_1088),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_1021),
.A2(n_961),
.B(n_1049),
.Y(n_1105)
);

NOR2x1_ASAP7_75t_L g1106 ( 
.A(n_1069),
.B(n_1075),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1060),
.B(n_1062),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_959),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_961),
.A2(n_1032),
.B(n_954),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_1032),
.A2(n_954),
.B(n_999),
.Y(n_1110)
);

O2A1O1Ixp33_ASAP7_75t_SL g1111 ( 
.A1(n_1002),
.A2(n_1019),
.B(n_989),
.C(n_977),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1062),
.A2(n_1064),
.B1(n_1083),
.B2(n_1031),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_985),
.B(n_952),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1070),
.A2(n_1088),
.B(n_1072),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1056),
.B(n_1079),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_1082),
.A2(n_1085),
.B(n_962),
.C(n_953),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_1017),
.Y(n_1117)
);

AO21x1_ASAP7_75t_L g1118 ( 
.A1(n_957),
.A2(n_1080),
.B(n_1072),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1073),
.B(n_1078),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_962),
.B(n_949),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_968),
.B(n_997),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1070),
.A2(n_988),
.B(n_1030),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_1011),
.A2(n_982),
.B(n_1026),
.C(n_963),
.Y(n_1123)
);

AND2x6_ASAP7_75t_L g1124 ( 
.A(n_970),
.B(n_1086),
.Y(n_1124)
);

AO31x2_ASAP7_75t_L g1125 ( 
.A1(n_1052),
.A2(n_1047),
.A3(n_1036),
.B(n_1003),
.Y(n_1125)
);

AO32x2_ASAP7_75t_L g1126 ( 
.A1(n_969),
.A2(n_1020),
.A3(n_1010),
.B1(n_1016),
.B2(n_1045),
.Y(n_1126)
);

INVx4_ASAP7_75t_L g1127 ( 
.A(n_970),
.Y(n_1127)
);

AOI21xp33_ASAP7_75t_L g1128 ( 
.A1(n_982),
.A2(n_1048),
.B(n_1003),
.Y(n_1128)
);

OA21x2_ASAP7_75t_L g1129 ( 
.A1(n_1000),
.A2(n_1050),
.B(n_1033),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_1086),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1040),
.A2(n_1016),
.B(n_1033),
.Y(n_1131)
);

INVx8_ASAP7_75t_L g1132 ( 
.A(n_1066),
.Y(n_1132)
);

AOI221x1_ASAP7_75t_L g1133 ( 
.A1(n_1023),
.A2(n_1000),
.B1(n_992),
.B2(n_1045),
.C(n_996),
.Y(n_1133)
);

INVx3_ASAP7_75t_SL g1134 ( 
.A(n_955),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_951),
.Y(n_1135)
);

HB1xp67_ASAP7_75t_L g1136 ( 
.A(n_964),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1006),
.A2(n_1051),
.B(n_1053),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_1071),
.Y(n_1138)
);

AOI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_978),
.A2(n_956),
.B1(n_1035),
.B2(n_1034),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1006),
.A2(n_996),
.B(n_1028),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1087),
.B(n_1037),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1028),
.A2(n_1061),
.B1(n_1084),
.B2(n_967),
.Y(n_1142)
);

AO21x1_ASAP7_75t_L g1143 ( 
.A1(n_1042),
.A2(n_1039),
.B(n_1076),
.Y(n_1143)
);

OA21x2_ASAP7_75t_L g1144 ( 
.A1(n_1042),
.A2(n_1043),
.B(n_1027),
.Y(n_1144)
);

OAI22x1_ASAP7_75t_L g1145 ( 
.A1(n_993),
.A2(n_980),
.B1(n_991),
.B2(n_971),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1046),
.A2(n_1045),
.B(n_1066),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1063),
.A2(n_1046),
.B(n_1058),
.C(n_1057),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1008),
.B(n_972),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1046),
.A2(n_976),
.B(n_979),
.C(n_994),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1024),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_1004),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1066),
.A2(n_998),
.B(n_995),
.Y(n_1152)
);

O2A1O1Ixp33_ASAP7_75t_SL g1153 ( 
.A1(n_1041),
.A2(n_1089),
.B(n_966),
.C(n_1081),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_990),
.Y(n_1154)
);

BUFx2_ASAP7_75t_R g1155 ( 
.A(n_1009),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_950),
.A2(n_1009),
.B(n_1014),
.Y(n_1156)
);

OAI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_1004),
.A2(n_972),
.B1(n_983),
.B2(n_1067),
.Y(n_1157)
);

OAI22x1_ASAP7_75t_L g1158 ( 
.A1(n_971),
.A2(n_950),
.B1(n_1012),
.B2(n_1014),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1012),
.A2(n_1004),
.B(n_986),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1074),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1055),
.A2(n_1059),
.B(n_948),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1055),
.A2(n_1059),
.B(n_948),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_989),
.A2(n_777),
.B(n_942),
.C(n_822),
.Y(n_1163)
);

O2A1O1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_989),
.A2(n_777),
.B(n_942),
.C(n_822),
.Y(n_1164)
);

OR2x2_ASAP7_75t_L g1165 ( 
.A(n_1069),
.B(n_1075),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_948),
.A2(n_777),
.B(n_1080),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1055),
.A2(n_1059),
.B(n_948),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_SL g1168 ( 
.A1(n_1002),
.A2(n_777),
.B(n_1019),
.C(n_989),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_959),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_948),
.A2(n_777),
.B(n_1080),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_991),
.Y(n_1171)
);

AO31x2_ASAP7_75t_L g1172 ( 
.A1(n_1005),
.A2(n_958),
.A3(n_988),
.B(n_999),
.Y(n_1172)
);

BUFx12f_ASAP7_75t_L g1173 ( 
.A(n_955),
.Y(n_1173)
);

INVx4_ASAP7_75t_L g1174 ( 
.A(n_970),
.Y(n_1174)
);

OR2x6_ASAP7_75t_L g1175 ( 
.A(n_1066),
.B(n_1015),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1073),
.B(n_1078),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_975),
.A2(n_942),
.B(n_1065),
.C(n_777),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1055),
.A2(n_1059),
.B(n_948),
.Y(n_1178)
);

OA21x2_ASAP7_75t_L g1179 ( 
.A1(n_984),
.A2(n_999),
.B(n_1044),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1055),
.A2(n_1059),
.B(n_948),
.Y(n_1180)
);

A2O1A1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_975),
.A2(n_942),
.B(n_1065),
.C(n_777),
.Y(n_1181)
);

NOR2x1_ASAP7_75t_R g1182 ( 
.A(n_993),
.B(n_1007),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_965),
.A2(n_1054),
.B(n_973),
.Y(n_1183)
);

AO31x2_ASAP7_75t_L g1184 ( 
.A1(n_1005),
.A2(n_958),
.A3(n_988),
.B(n_999),
.Y(n_1184)
);

AOI31xp67_ASAP7_75t_L g1185 ( 
.A1(n_975),
.A2(n_989),
.A3(n_1016),
.B(n_903),
.Y(n_1185)
);

AO21x1_ASAP7_75t_L g1186 ( 
.A1(n_1068),
.A2(n_777),
.B(n_1077),
.Y(n_1186)
);

NAND2xp33_ASAP7_75t_L g1187 ( 
.A(n_975),
.B(n_777),
.Y(n_1187)
);

NOR3xp33_ASAP7_75t_L g1188 ( 
.A(n_975),
.B(n_777),
.C(n_822),
.Y(n_1188)
);

AO31x2_ASAP7_75t_L g1189 ( 
.A1(n_1005),
.A2(n_958),
.A3(n_988),
.B(n_999),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1055),
.A2(n_1059),
.B(n_948),
.Y(n_1190)
);

CKINVDCx8_ASAP7_75t_R g1191 ( 
.A(n_986),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1055),
.A2(n_1059),
.B(n_948),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1065),
.B(n_942),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1065),
.B(n_942),
.Y(n_1194)
);

NOR2xp67_ASAP7_75t_L g1195 ( 
.A(n_975),
.B(n_923),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_SL g1196 ( 
.A1(n_953),
.A2(n_1019),
.B(n_1002),
.Y(n_1196)
);

AOI21xp33_ASAP7_75t_SL g1197 ( 
.A1(n_1074),
.A2(n_822),
.B(n_620),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_959),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1055),
.A2(n_1059),
.B(n_948),
.Y(n_1199)
);

NAND2x1p5_ASAP7_75t_L g1200 ( 
.A(n_970),
.B(n_905),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_SL g1201 ( 
.A1(n_975),
.A2(n_1007),
.B1(n_620),
.B2(n_942),
.Y(n_1201)
);

BUFx4f_ASAP7_75t_SL g1202 ( 
.A(n_960),
.Y(n_1202)
);

AOI221x1_ASAP7_75t_L g1203 ( 
.A1(n_953),
.A2(n_777),
.B1(n_1070),
.B2(n_1072),
.C(n_948),
.Y(n_1203)
);

AOI221x1_ASAP7_75t_L g1204 ( 
.A1(n_953),
.A2(n_777),
.B1(n_1070),
.B2(n_1072),
.C(n_948),
.Y(n_1204)
);

AO31x2_ASAP7_75t_L g1205 ( 
.A1(n_1005),
.A2(n_958),
.A3(n_988),
.B(n_999),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1065),
.B(n_942),
.Y(n_1206)
);

OR2x2_ASAP7_75t_L g1207 ( 
.A(n_1069),
.B(n_1075),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_965),
.A2(n_1054),
.B(n_973),
.Y(n_1208)
);

AO31x2_ASAP7_75t_L g1209 ( 
.A1(n_1005),
.A2(n_958),
.A3(n_988),
.B(n_999),
.Y(n_1209)
);

AOI21xp33_ASAP7_75t_L g1210 ( 
.A1(n_975),
.A2(n_777),
.B(n_1068),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_960),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_964),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1065),
.B(n_942),
.Y(n_1213)
);

NOR4xp25_ASAP7_75t_L g1214 ( 
.A(n_1068),
.B(n_1082),
.C(n_1077),
.D(n_898),
.Y(n_1214)
);

AO31x2_ASAP7_75t_L g1215 ( 
.A1(n_1005),
.A2(n_958),
.A3(n_988),
.B(n_999),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_948),
.A2(n_777),
.B(n_1080),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_948),
.A2(n_777),
.B(n_1080),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_965),
.A2(n_1054),
.B(n_973),
.Y(n_1218)
);

AO31x2_ASAP7_75t_L g1219 ( 
.A1(n_1005),
.A2(n_958),
.A3(n_988),
.B(n_999),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_965),
.A2(n_1054),
.B(n_973),
.Y(n_1220)
);

INVxp67_ASAP7_75t_SL g1221 ( 
.A(n_962),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1017),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_965),
.A2(n_1054),
.B(n_973),
.Y(n_1223)
);

AOI221xp5_ASAP7_75t_SL g1224 ( 
.A1(n_1011),
.A2(n_1002),
.B1(n_947),
.B2(n_1062),
.C(n_1060),
.Y(n_1224)
);

AO32x2_ASAP7_75t_L g1225 ( 
.A1(n_953),
.A2(n_1029),
.A3(n_838),
.B1(n_1036),
.B2(n_1049),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1108),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1169),
.Y(n_1227)
);

INVx6_ASAP7_75t_L g1228 ( 
.A(n_1132),
.Y(n_1228)
);

NAND2x1p5_ASAP7_75t_L g1229 ( 
.A(n_1156),
.B(n_1099),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1198),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_SL g1231 ( 
.A1(n_1201),
.A2(n_1194),
.B1(n_1193),
.B2(n_1187),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1188),
.A2(n_1195),
.B1(n_1201),
.B2(n_1210),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1206),
.A2(n_1213),
.B1(n_1177),
.B2(n_1181),
.Y(n_1233)
);

BUFx12f_ASAP7_75t_L g1234 ( 
.A(n_1173),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_SL g1235 ( 
.A1(n_1102),
.A2(n_1112),
.B1(n_1121),
.B2(n_1160),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1093),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1101),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1102),
.B(n_1107),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1195),
.A2(n_1197),
.B1(n_1139),
.B2(n_1106),
.Y(n_1239)
);

INVx3_ASAP7_75t_L g1240 ( 
.A(n_1132),
.Y(n_1240)
);

CKINVDCx11_ASAP7_75t_R g1241 ( 
.A(n_1191),
.Y(n_1241)
);

INVx4_ASAP7_75t_L g1242 ( 
.A(n_1124),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_SL g1243 ( 
.A1(n_1112),
.A2(n_1221),
.B1(n_1115),
.B2(n_1159),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1210),
.A2(n_1090),
.B1(n_1186),
.B2(n_1176),
.Y(n_1244)
);

INVx2_ASAP7_75t_SL g1245 ( 
.A(n_1138),
.Y(n_1245)
);

INVx6_ASAP7_75t_L g1246 ( 
.A(n_1175),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1090),
.A2(n_1113),
.B1(n_1139),
.B2(n_1119),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1120),
.A2(n_1145),
.B1(n_1131),
.B2(n_1137),
.Y(n_1248)
);

INVxp67_ASAP7_75t_SL g1249 ( 
.A(n_1136),
.Y(n_1249)
);

CKINVDCx11_ASAP7_75t_R g1250 ( 
.A(n_1134),
.Y(n_1250)
);

INVx6_ASAP7_75t_L g1251 ( 
.A(n_1175),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1150),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1165),
.A2(n_1207),
.B1(n_1096),
.B2(n_1179),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1163),
.A2(n_1164),
.B1(n_1196),
.B2(n_1149),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1141),
.A2(n_1147),
.B1(n_1123),
.B2(n_1148),
.Y(n_1255)
);

BUFx8_ASAP7_75t_L g1256 ( 
.A(n_1126),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1129),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1125),
.Y(n_1258)
);

BUFx3_ASAP7_75t_L g1259 ( 
.A(n_1211),
.Y(n_1259)
);

OAI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1096),
.A2(n_1175),
.B1(n_1159),
.B2(n_1133),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_1130),
.Y(n_1261)
);

CKINVDCx14_ASAP7_75t_R g1262 ( 
.A(n_1154),
.Y(n_1262)
);

OAI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1212),
.A2(n_1202),
.B1(n_1135),
.B2(n_1146),
.Y(n_1263)
);

INVx5_ASAP7_75t_L g1264 ( 
.A(n_1124),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1224),
.B(n_1168),
.Y(n_1265)
);

AOI22xp5_ASAP7_75t_SL g1266 ( 
.A1(n_1158),
.A2(n_1151),
.B1(n_1152),
.B2(n_1142),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1116),
.A2(n_1155),
.B1(n_1157),
.B2(n_1140),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_1151),
.Y(n_1268)
);

BUFx8_ASAP7_75t_L g1269 ( 
.A(n_1126),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1224),
.B(n_1126),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_SL g1271 ( 
.A1(n_1100),
.A2(n_1170),
.B1(n_1217),
.B2(n_1216),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1130),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_1124),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_1124),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1118),
.A2(n_1128),
.B1(n_1216),
.B2(n_1166),
.Y(n_1275)
);

BUFx10_ASAP7_75t_L g1276 ( 
.A(n_1130),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1128),
.A2(n_1170),
.B1(n_1166),
.B2(n_1143),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1129),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1122),
.A2(n_1144),
.B1(n_1104),
.B2(n_1091),
.Y(n_1279)
);

CKINVDCx11_ASAP7_75t_R g1280 ( 
.A(n_1127),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1214),
.B(n_1111),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1144),
.Y(n_1282)
);

OAI22xp33_ASAP7_75t_SL g1283 ( 
.A1(n_1214),
.A2(n_1185),
.B1(n_1200),
.B2(n_1098),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1225),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1153),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1104),
.A2(n_1222),
.B1(n_1117),
.B2(n_1098),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1222),
.A2(n_1114),
.B1(n_1103),
.B2(n_1110),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1109),
.Y(n_1288)
);

INVx3_ASAP7_75t_L g1289 ( 
.A(n_1127),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1174),
.A2(n_1105),
.B1(n_1162),
.B2(n_1095),
.Y(n_1290)
);

INVx2_ASAP7_75t_SL g1291 ( 
.A(n_1174),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1161),
.A2(n_1199),
.B1(n_1192),
.B2(n_1167),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1178),
.A2(n_1190),
.B1(n_1180),
.B2(n_1094),
.Y(n_1293)
);

OAI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1203),
.A2(n_1204),
.B(n_1208),
.Y(n_1294)
);

OAI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1182),
.A2(n_1225),
.B1(n_1172),
.B2(n_1215),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1184),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1092),
.A2(n_1183),
.B1(n_1223),
.B2(n_1220),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_SL g1298 ( 
.A1(n_1225),
.A2(n_1182),
.B1(n_1184),
.B2(n_1189),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1218),
.A2(n_1189),
.B1(n_1205),
.B2(n_1209),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_1189),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1205),
.Y(n_1301)
);

CKINVDCx11_ASAP7_75t_R g1302 ( 
.A(n_1209),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1215),
.A2(n_1188),
.B1(n_1187),
.B2(n_942),
.Y(n_1303)
);

BUFx2_ASAP7_75t_SL g1304 ( 
.A(n_1219),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1219),
.A2(n_1188),
.B1(n_1187),
.B2(n_942),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1188),
.A2(n_1187),
.B1(n_942),
.B2(n_777),
.Y(n_1306)
);

BUFx2_ASAP7_75t_R g1307 ( 
.A(n_1191),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1108),
.Y(n_1308)
);

BUFx4f_ASAP7_75t_SL g1309 ( 
.A(n_1173),
.Y(n_1309)
);

INVxp67_ASAP7_75t_SL g1310 ( 
.A(n_1136),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1108),
.Y(n_1311)
);

INVx5_ASAP7_75t_L g1312 ( 
.A(n_1124),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1138),
.Y(n_1313)
);

CKINVDCx11_ASAP7_75t_R g1314 ( 
.A(n_1191),
.Y(n_1314)
);

BUFx12f_ASAP7_75t_L g1315 ( 
.A(n_1173),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1193),
.A2(n_1194),
.B1(n_942),
.B2(n_975),
.Y(n_1316)
);

BUFx10_ASAP7_75t_L g1317 ( 
.A(n_1113),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1188),
.A2(n_1187),
.B1(n_942),
.B2(n_777),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1193),
.B(n_1065),
.Y(n_1319)
);

INVxp67_ASAP7_75t_SL g1320 ( 
.A(n_1136),
.Y(n_1320)
);

AOI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1188),
.A2(n_975),
.B1(n_1201),
.B2(n_1194),
.Y(n_1321)
);

BUFx2_ASAP7_75t_SL g1322 ( 
.A(n_1096),
.Y(n_1322)
);

BUFx12f_ASAP7_75t_L g1323 ( 
.A(n_1173),
.Y(n_1323)
);

CKINVDCx6p67_ASAP7_75t_R g1324 ( 
.A(n_1134),
.Y(n_1324)
);

INVx6_ASAP7_75t_L g1325 ( 
.A(n_1132),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1108),
.Y(n_1326)
);

INVx6_ASAP7_75t_L g1327 ( 
.A(n_1132),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1201),
.A2(n_1193),
.B1(n_1194),
.B2(n_942),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1188),
.A2(n_1187),
.B1(n_942),
.B2(n_777),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1188),
.A2(n_1187),
.B1(n_942),
.B2(n_777),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1188),
.A2(n_1187),
.B1(n_942),
.B2(n_777),
.Y(n_1331)
);

OAI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1188),
.A2(n_777),
.B(n_942),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1108),
.Y(n_1333)
);

CKINVDCx11_ASAP7_75t_R g1334 ( 
.A(n_1191),
.Y(n_1334)
);

BUFx8_ASAP7_75t_L g1335 ( 
.A(n_1173),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1097),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_1138),
.Y(n_1337)
);

BUFx2_ASAP7_75t_L g1338 ( 
.A(n_1171),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1257),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1282),
.Y(n_1340)
);

INVx2_ASAP7_75t_SL g1341 ( 
.A(n_1246),
.Y(n_1341)
);

INVxp33_ASAP7_75t_L g1342 ( 
.A(n_1313),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1257),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1294),
.A2(n_1297),
.B(n_1292),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1278),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1270),
.B(n_1298),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1319),
.B(n_1316),
.Y(n_1347)
);

OAI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1332),
.A2(n_1318),
.B(n_1306),
.Y(n_1348)
);

BUFx2_ASAP7_75t_L g1349 ( 
.A(n_1300),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1293),
.A2(n_1290),
.B(n_1287),
.Y(n_1350)
);

AOI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1254),
.A2(n_1281),
.B(n_1285),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1284),
.B(n_1296),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1233),
.B(n_1235),
.Y(n_1353)
);

INVx1_ASAP7_75t_SL g1354 ( 
.A(n_1317),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1301),
.Y(n_1355)
);

CKINVDCx11_ASAP7_75t_R g1356 ( 
.A(n_1241),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1288),
.A2(n_1279),
.B(n_1258),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1270),
.B(n_1284),
.Y(n_1358)
);

INVx2_ASAP7_75t_SL g1359 ( 
.A(n_1246),
.Y(n_1359)
);

AOI22xp5_ASAP7_75t_SL g1360 ( 
.A1(n_1239),
.A2(n_1322),
.B1(n_1255),
.B2(n_1267),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1247),
.B(n_1231),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_1264),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1237),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1304),
.Y(n_1364)
);

AOI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1265),
.A2(n_1238),
.B(n_1252),
.Y(n_1365)
);

BUFx12f_ASAP7_75t_L g1366 ( 
.A(n_1241),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1302),
.Y(n_1367)
);

OAI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1329),
.A2(n_1330),
.B(n_1331),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1236),
.Y(n_1369)
);

AOI21xp33_ASAP7_75t_L g1370 ( 
.A1(n_1321),
.A2(n_1328),
.B(n_1232),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1295),
.B(n_1277),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1275),
.A2(n_1299),
.B(n_1229),
.Y(n_1372)
);

OR2x6_ASAP7_75t_L g1373 ( 
.A(n_1229),
.B(n_1251),
.Y(n_1373)
);

NAND2x1_ASAP7_75t_L g1374 ( 
.A(n_1242),
.B(n_1251),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1271),
.A2(n_1305),
.B(n_1303),
.Y(n_1375)
);

INVxp67_ASAP7_75t_L g1376 ( 
.A(n_1338),
.Y(n_1376)
);

AOI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1226),
.A2(n_1227),
.B(n_1308),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1264),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1244),
.A2(n_1243),
.B(n_1248),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1240),
.B(n_1266),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_1264),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1230),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1311),
.Y(n_1383)
);

OAI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1253),
.A2(n_1260),
.B(n_1286),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1326),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1333),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1283),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1256),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1256),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1249),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1269),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1269),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_SL g1393 ( 
.A1(n_1269),
.A2(n_1228),
.B1(n_1325),
.B2(n_1327),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1310),
.B(n_1320),
.Y(n_1394)
);

BUFx2_ASAP7_75t_L g1395 ( 
.A(n_1263),
.Y(n_1395)
);

BUFx12f_ASAP7_75t_L g1396 ( 
.A(n_1314),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1337),
.B(n_1245),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1317),
.B(n_1245),
.Y(n_1398)
);

NOR2x1_ASAP7_75t_L g1399 ( 
.A(n_1354),
.B(n_1336),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1358),
.B(n_1324),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1361),
.A2(n_1262),
.B1(n_1324),
.B2(n_1268),
.Y(n_1401)
);

OAI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1348),
.A2(n_1291),
.B(n_1262),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1369),
.Y(n_1403)
);

OR2x6_ASAP7_75t_L g1404 ( 
.A(n_1373),
.B(n_1228),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1344),
.A2(n_1289),
.B(n_1312),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_SL g1406 ( 
.A1(n_1347),
.A2(n_1309),
.B1(n_1234),
.B2(n_1323),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_1353),
.B(n_1228),
.Y(n_1407)
);

CKINVDCx10_ASAP7_75t_R g1408 ( 
.A(n_1356),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1367),
.B(n_1268),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1370),
.A2(n_1250),
.B1(n_1315),
.B2(n_1234),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1358),
.B(n_1261),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1346),
.B(n_1261),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_L g1413 ( 
.A(n_1395),
.B(n_1327),
.Y(n_1413)
);

AO21x2_ASAP7_75t_L g1414 ( 
.A1(n_1365),
.A2(n_1274),
.B(n_1273),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1394),
.B(n_1390),
.Y(n_1415)
);

OAI21xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1368),
.A2(n_1291),
.B(n_1289),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1355),
.Y(n_1417)
);

NOR2xp67_ASAP7_75t_L g1418 ( 
.A(n_1398),
.B(n_1323),
.Y(n_1418)
);

OA21x2_ASAP7_75t_L g1419 ( 
.A1(n_1344),
.A2(n_1272),
.B(n_1273),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1366),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1367),
.B(n_1272),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1352),
.B(n_1259),
.Y(n_1422)
);

O2A1O1Ixp33_ASAP7_75t_L g1423 ( 
.A1(n_1379),
.A2(n_1375),
.B(n_1384),
.C(n_1395),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1376),
.B(n_1336),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1360),
.A2(n_1259),
.B(n_1250),
.Y(n_1425)
);

OAI211xp5_ASAP7_75t_SL g1426 ( 
.A1(n_1387),
.A2(n_1280),
.B(n_1334),
.C(n_1314),
.Y(n_1426)
);

AO21x2_ASAP7_75t_L g1427 ( 
.A1(n_1364),
.A2(n_1387),
.B(n_1350),
.Y(n_1427)
);

A2O1A1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1371),
.A2(n_1325),
.B(n_1280),
.C(n_1335),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1371),
.A2(n_1315),
.B1(n_1307),
.B2(n_1335),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1374),
.A2(n_1276),
.B(n_1335),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1383),
.B(n_1334),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_SL g1432 ( 
.A(n_1366),
.B(n_1396),
.Y(n_1432)
);

INVx1_ASAP7_75t_SL g1433 ( 
.A(n_1397),
.Y(n_1433)
);

A2O1A1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1372),
.A2(n_1380),
.B(n_1391),
.C(n_1389),
.Y(n_1434)
);

AOI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1380),
.A2(n_1366),
.B1(n_1396),
.B2(n_1359),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1363),
.Y(n_1436)
);

AO32x2_ASAP7_75t_L g1437 ( 
.A1(n_1341),
.A2(n_1359),
.A3(n_1349),
.B1(n_1355),
.B2(n_1339),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1393),
.A2(n_1342),
.B1(n_1380),
.B2(n_1389),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1351),
.B(n_1380),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1383),
.B(n_1386),
.Y(n_1440)
);

AO21x2_ASAP7_75t_L g1441 ( 
.A1(n_1364),
.A2(n_1350),
.B(n_1357),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1436),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1415),
.B(n_1339),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1403),
.Y(n_1444)
);

INVx4_ASAP7_75t_L g1445 ( 
.A(n_1404),
.Y(n_1445)
);

INVx2_ASAP7_75t_SL g1446 ( 
.A(n_1417),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1423),
.A2(n_1391),
.B1(n_1389),
.B2(n_1392),
.Y(n_1447)
);

OR2x2_ASAP7_75t_SL g1448 ( 
.A(n_1419),
.B(n_1391),
.Y(n_1448)
);

BUFx2_ASAP7_75t_L g1449 ( 
.A(n_1437),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1407),
.B(n_1382),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1437),
.B(n_1339),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1437),
.Y(n_1452)
);

INVxp67_ASAP7_75t_L g1453 ( 
.A(n_1439),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1425),
.A2(n_1396),
.B1(n_1388),
.B2(n_1392),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1410),
.A2(n_1388),
.B1(n_1382),
.B2(n_1385),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_SL g1456 ( 
.A(n_1416),
.B(n_1341),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1441),
.B(n_1343),
.Y(n_1457)
);

NAND3xp33_ASAP7_75t_L g1458 ( 
.A(n_1402),
.B(n_1410),
.C(n_1428),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1427),
.B(n_1345),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1440),
.Y(n_1460)
);

NAND2x1_ASAP7_75t_L g1461 ( 
.A(n_1404),
.B(n_1381),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1419),
.B(n_1411),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1419),
.B(n_1345),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1411),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1439),
.B(n_1340),
.Y(n_1465)
);

AOI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1459),
.A2(n_1418),
.B(n_1377),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1462),
.B(n_1434),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1462),
.B(n_1434),
.Y(n_1468)
);

OAI33xp33_ASAP7_75t_L g1469 ( 
.A1(n_1447),
.A2(n_1429),
.A3(n_1401),
.B1(n_1426),
.B2(n_1431),
.B3(n_1406),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1460),
.B(n_1414),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1460),
.B(n_1414),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1462),
.B(n_1412),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1446),
.Y(n_1473)
);

OR2x6_ASAP7_75t_L g1474 ( 
.A(n_1461),
.B(n_1405),
.Y(n_1474)
);

INVx3_ASAP7_75t_L g1475 ( 
.A(n_1442),
.Y(n_1475)
);

BUFx2_ASAP7_75t_L g1476 ( 
.A(n_1448),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1444),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1451),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1458),
.A2(n_1447),
.B1(n_1407),
.B2(n_1455),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1458),
.A2(n_1433),
.B1(n_1438),
.B2(n_1400),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1448),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1451),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1449),
.B(n_1405),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_1448),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1449),
.B(n_1452),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1444),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1449),
.B(n_1422),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1452),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1446),
.Y(n_1489)
);

BUFx3_ASAP7_75t_L g1490 ( 
.A(n_1461),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1457),
.Y(n_1491)
);

INVx1_ASAP7_75t_SL g1492 ( 
.A(n_1463),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1467),
.B(n_1453),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1473),
.Y(n_1494)
);

INVxp33_ASAP7_75t_L g1495 ( 
.A(n_1480),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1473),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1474),
.B(n_1459),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1477),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1467),
.B(n_1453),
.Y(n_1499)
);

NAND2xp33_ASAP7_75t_SL g1500 ( 
.A(n_1479),
.B(n_1420),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1488),
.B(n_1446),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_1476),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1492),
.B(n_1465),
.Y(n_1503)
);

INVx2_ASAP7_75t_SL g1504 ( 
.A(n_1489),
.Y(n_1504)
);

NAND4xp25_ASAP7_75t_SL g1505 ( 
.A(n_1479),
.B(n_1454),
.C(n_1428),
.D(n_1435),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1467),
.B(n_1468),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1467),
.B(n_1464),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1477),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1475),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1468),
.B(n_1464),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1475),
.Y(n_1511)
);

NAND3xp33_ASAP7_75t_L g1512 ( 
.A(n_1480),
.B(n_1455),
.C(n_1454),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1488),
.B(n_1478),
.Y(n_1513)
);

INVx1_ASAP7_75t_SL g1514 ( 
.A(n_1476),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1477),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1492),
.B(n_1465),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1487),
.B(n_1443),
.Y(n_1517)
);

INVx4_ASAP7_75t_L g1518 ( 
.A(n_1490),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1478),
.B(n_1459),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1486),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1486),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1487),
.B(n_1443),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1486),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1490),
.Y(n_1524)
);

INVx1_ASAP7_75t_SL g1525 ( 
.A(n_1476),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1469),
.B(n_1432),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1495),
.B(n_1450),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1494),
.Y(n_1528)
);

INVx1_ASAP7_75t_SL g1529 ( 
.A(n_1524),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1506),
.B(n_1485),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1494),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1496),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1496),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1513),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1502),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1517),
.B(n_1470),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1498),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1493),
.B(n_1487),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_L g1539 ( 
.A(n_1526),
.B(n_1469),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1506),
.B(n_1485),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1518),
.B(n_1490),
.Y(n_1541)
);

OAI22xp33_ASAP7_75t_SL g1542 ( 
.A1(n_1502),
.A2(n_1481),
.B1(n_1484),
.B2(n_1488),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1498),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1508),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1517),
.B(n_1470),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1508),
.Y(n_1546)
);

INVxp67_ASAP7_75t_L g1547 ( 
.A(n_1512),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1522),
.B(n_1470),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1506),
.B(n_1485),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1513),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_1524),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1493),
.B(n_1485),
.Y(n_1552)
);

AOI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1500),
.A2(n_1469),
.B1(n_1445),
.B2(n_1450),
.Y(n_1553)
);

CKINVDCx20_ASAP7_75t_R g1554 ( 
.A(n_1512),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1493),
.B(n_1490),
.Y(n_1555)
);

NOR2x1p5_ASAP7_75t_SL g1556 ( 
.A(n_1513),
.B(n_1509),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1515),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1522),
.B(n_1471),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1515),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1504),
.Y(n_1560)
);

NAND4xp25_ASAP7_75t_L g1561 ( 
.A(n_1514),
.B(n_1481),
.C(n_1484),
.D(n_1413),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1520),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1499),
.B(n_1472),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1514),
.B(n_1471),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1525),
.Y(n_1565)
);

OR2x6_ASAP7_75t_L g1566 ( 
.A(n_1518),
.B(n_1474),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1499),
.B(n_1490),
.Y(n_1567)
);

INVx2_ASAP7_75t_SL g1568 ( 
.A(n_1504),
.Y(n_1568)
);

INVx2_ASAP7_75t_SL g1569 ( 
.A(n_1568),
.Y(n_1569)
);

OAI21xp33_ASAP7_75t_L g1570 ( 
.A1(n_1547),
.A2(n_1505),
.B(n_1499),
.Y(n_1570)
);

OAI21xp33_ASAP7_75t_SL g1571 ( 
.A1(n_1561),
.A2(n_1525),
.B(n_1505),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1539),
.B(n_1507),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1537),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1543),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1539),
.B(n_1507),
.Y(n_1575)
);

INVx1_ASAP7_75t_SL g1576 ( 
.A(n_1529),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1530),
.B(n_1518),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1544),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1546),
.Y(n_1579)
);

NAND2xp33_ASAP7_75t_SL g1580 ( 
.A(n_1554),
.B(n_1420),
.Y(n_1580)
);

NOR2xp67_ASAP7_75t_SL g1581 ( 
.A(n_1535),
.B(n_1430),
.Y(n_1581)
);

NAND4xp25_ASAP7_75t_L g1582 ( 
.A(n_1553),
.B(n_1518),
.C(n_1481),
.D(n_1484),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1557),
.Y(n_1583)
);

OR2x2_ASAP7_75t_SL g1584 ( 
.A(n_1527),
.B(n_1501),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1530),
.B(n_1540),
.Y(n_1585)
);

NAND3xp33_ASAP7_75t_L g1586 ( 
.A(n_1554),
.B(n_1481),
.C(n_1399),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1559),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1563),
.B(n_1503),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1562),
.Y(n_1589)
);

INVx1_ASAP7_75t_SL g1590 ( 
.A(n_1551),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1568),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1528),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1531),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_SL g1594 ( 
.A(n_1542),
.B(n_1504),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1532),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1565),
.B(n_1507),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1538),
.B(n_1503),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1533),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_SL g1599 ( 
.A(n_1541),
.B(n_1501),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1555),
.B(n_1510),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1540),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1549),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1555),
.B(n_1510),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1585),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1573),
.Y(n_1605)
);

INVx2_ASAP7_75t_SL g1606 ( 
.A(n_1569),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_L g1607 ( 
.A(n_1570),
.B(n_1408),
.Y(n_1607)
);

AOI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1571),
.A2(n_1567),
.B1(n_1541),
.B2(n_1549),
.Y(n_1608)
);

AOI21xp33_ASAP7_75t_L g1609 ( 
.A1(n_1594),
.A2(n_1541),
.B(n_1566),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1577),
.B(n_1567),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1574),
.Y(n_1611)
);

AOI32xp33_ASAP7_75t_L g1612 ( 
.A1(n_1580),
.A2(n_1594),
.A3(n_1576),
.B1(n_1590),
.B2(n_1572),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1578),
.Y(n_1613)
);

OAI21xp33_ASAP7_75t_L g1614 ( 
.A1(n_1582),
.A2(n_1556),
.B(n_1552),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1579),
.Y(n_1615)
);

INVx3_ASAP7_75t_L g1616 ( 
.A(n_1585),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1583),
.Y(n_1617)
);

OAI21xp5_ASAP7_75t_SL g1618 ( 
.A1(n_1586),
.A2(n_1575),
.B(n_1580),
.Y(n_1618)
);

INVx1_ASAP7_75t_SL g1619 ( 
.A(n_1584),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1581),
.B(n_1552),
.Y(n_1620)
);

AOI21xp33_ASAP7_75t_L g1621 ( 
.A1(n_1592),
.A2(n_1566),
.B(n_1560),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1585),
.Y(n_1622)
);

AOI21xp33_ASAP7_75t_L g1623 ( 
.A1(n_1593),
.A2(n_1566),
.B(n_1560),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1569),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1577),
.B(n_1601),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1595),
.B(n_1510),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1587),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1596),
.B(n_1534),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1605),
.Y(n_1629)
);

OAI221xp5_ASAP7_75t_L g1630 ( 
.A1(n_1612),
.A2(n_1599),
.B1(n_1598),
.B2(n_1600),
.C(n_1603),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1616),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1605),
.Y(n_1632)
);

O2A1O1Ixp5_ASAP7_75t_L g1633 ( 
.A1(n_1609),
.A2(n_1599),
.B(n_1591),
.C(n_1550),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1611),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1616),
.B(n_1591),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1616),
.B(n_1602),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1610),
.B(n_1566),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1619),
.B(n_1589),
.Y(n_1638)
);

AOI32xp33_ASAP7_75t_L g1639 ( 
.A1(n_1614),
.A2(n_1483),
.A3(n_1497),
.B1(n_1534),
.B2(n_1550),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1611),
.Y(n_1640)
);

OAI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1608),
.A2(n_1588),
.B1(n_1597),
.B2(n_1474),
.Y(n_1641)
);

OAI31xp33_ASAP7_75t_L g1642 ( 
.A1(n_1618),
.A2(n_1620),
.A3(n_1621),
.B(n_1623),
.Y(n_1642)
);

AO22x1_ASAP7_75t_L g1643 ( 
.A1(n_1607),
.A2(n_1497),
.B1(n_1483),
.B2(n_1492),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1624),
.B(n_1606),
.Y(n_1644)
);

AOI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1604),
.A2(n_1564),
.B(n_1471),
.Y(n_1645)
);

OAI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1604),
.A2(n_1474),
.B1(n_1478),
.B2(n_1482),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1627),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1631),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1635),
.B(n_1622),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1636),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1635),
.B(n_1622),
.Y(n_1651)
);

INVxp67_ASAP7_75t_SL g1652 ( 
.A(n_1644),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1636),
.Y(n_1653)
);

OAI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1630),
.A2(n_1606),
.B1(n_1624),
.B2(n_1627),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1647),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1647),
.Y(n_1656)
);

AOI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1637),
.A2(n_1625),
.B1(n_1610),
.B2(n_1626),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1629),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1632),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1649),
.B(n_1638),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1650),
.Y(n_1661)
);

NOR3xp33_ASAP7_75t_L g1662 ( 
.A(n_1654),
.B(n_1633),
.C(n_1634),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1652),
.B(n_1640),
.Y(n_1663)
);

INVxp67_ASAP7_75t_L g1664 ( 
.A(n_1649),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1651),
.B(n_1642),
.Y(n_1665)
);

OAI21xp33_ASAP7_75t_L g1666 ( 
.A1(n_1657),
.A2(n_1639),
.B(n_1625),
.Y(n_1666)
);

NOR4xp25_ASAP7_75t_L g1667 ( 
.A(n_1654),
.B(n_1613),
.C(n_1615),
.D(n_1617),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1653),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_SL g1669 ( 
.A(n_1664),
.B(n_1651),
.Y(n_1669)
);

OAI211xp5_ASAP7_75t_L g1670 ( 
.A1(n_1662),
.A2(n_1648),
.B(n_1656),
.C(n_1655),
.Y(n_1670)
);

AOI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1666),
.A2(n_1637),
.B1(n_1641),
.B2(n_1659),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1660),
.B(n_1658),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1661),
.Y(n_1673)
);

OAI21xp5_ASAP7_75t_SL g1674 ( 
.A1(n_1671),
.A2(n_1665),
.B(n_1663),
.Y(n_1674)
);

OAI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1669),
.A2(n_1628),
.B1(n_1668),
.B2(n_1645),
.Y(n_1675)
);

OAI21x1_ASAP7_75t_SL g1676 ( 
.A1(n_1673),
.A2(n_1667),
.B(n_1628),
.Y(n_1676)
);

NAND3xp33_ASAP7_75t_L g1677 ( 
.A(n_1670),
.B(n_1643),
.C(n_1646),
.Y(n_1677)
);

NOR3xp33_ASAP7_75t_L g1678 ( 
.A(n_1672),
.B(n_1643),
.C(n_1564),
.Y(n_1678)
);

AOI211xp5_ASAP7_75t_L g1679 ( 
.A1(n_1670),
.A2(n_1409),
.B(n_1421),
.C(n_1545),
.Y(n_1679)
);

NOR2xp67_ASAP7_75t_L g1680 ( 
.A(n_1677),
.B(n_1536),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1675),
.Y(n_1681)
);

NAND4xp75_ASAP7_75t_L g1682 ( 
.A(n_1674),
.B(n_1483),
.C(n_1456),
.D(n_1424),
.Y(n_1682)
);

NOR2x1_ASAP7_75t_L g1683 ( 
.A(n_1676),
.B(n_1501),
.Y(n_1683)
);

AND2x4_ASAP7_75t_L g1684 ( 
.A(n_1678),
.B(n_1558),
.Y(n_1684)
);

NOR3xp33_ASAP7_75t_L g1685 ( 
.A(n_1681),
.B(n_1679),
.C(n_1545),
.Y(n_1685)
);

NAND3xp33_ASAP7_75t_L g1686 ( 
.A(n_1683),
.B(n_1548),
.C(n_1536),
.Y(n_1686)
);

NAND3x1_ASAP7_75t_L g1687 ( 
.A(n_1680),
.B(n_1519),
.C(n_1516),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1687),
.Y(n_1688)
);

OAI22x1_ASAP7_75t_L g1689 ( 
.A1(n_1688),
.A2(n_1684),
.B1(n_1686),
.B2(n_1685),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1689),
.B(n_1682),
.Y(n_1690)
);

INVx2_ASAP7_75t_SL g1691 ( 
.A(n_1690),
.Y(n_1691)
);

OAI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1691),
.A2(n_1548),
.B(n_1558),
.Y(n_1692)
);

AO21x2_ASAP7_75t_L g1693 ( 
.A1(n_1692),
.A2(n_1511),
.B(n_1509),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_SL g1694 ( 
.A1(n_1692),
.A2(n_1497),
.B1(n_1483),
.B2(n_1489),
.Y(n_1694)
);

AOI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1694),
.A2(n_1516),
.B(n_1497),
.Y(n_1695)
);

OA22x2_ASAP7_75t_L g1696 ( 
.A1(n_1693),
.A2(n_1497),
.B1(n_1509),
.B2(n_1511),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1696),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1695),
.Y(n_1698)
);

OAI221xp5_ASAP7_75t_R g1699 ( 
.A1(n_1698),
.A2(n_1511),
.B1(n_1466),
.B2(n_1491),
.C(n_1520),
.Y(n_1699)
);

OAI221xp5_ASAP7_75t_R g1700 ( 
.A1(n_1697),
.A2(n_1466),
.B1(n_1491),
.B2(n_1521),
.C(n_1523),
.Y(n_1700)
);

AOI211xp5_ASAP7_75t_L g1701 ( 
.A1(n_1700),
.A2(n_1699),
.B(n_1362),
.C(n_1378),
.Y(n_1701)
);


endmodule