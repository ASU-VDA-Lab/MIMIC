module fake_jpeg_28611_n_61 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_61);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_61;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_48;
wire n_35;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

INVx2_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_19),
.B(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_1),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_1),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_11),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_11),
.B1(n_15),
.B2(n_17),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_22),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_7),
.B1(n_26),
.B2(n_32),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_30),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_42),
.B(n_43),
.Y(n_46)
);

AND2x6_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_23),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_40),
.C(n_41),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_25),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_27),
.C(n_20),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_31),
.A2(n_26),
.B1(n_14),
.B2(n_21),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_SL g45 ( 
.A(n_40),
.B(n_29),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_39),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_42),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_48),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_52),
.B(n_33),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_51),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_33),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_44),
.B1(n_34),
.B2(n_35),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_44),
.C(n_46),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_54),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_56),
.B(n_57),
.Y(n_59)
);

AOI322xp5_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_7),
.A3(n_30),
.B1(n_34),
.B2(n_35),
.C1(n_55),
.C2(n_51),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_35),
.C(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_59),
.Y(n_61)
);


endmodule