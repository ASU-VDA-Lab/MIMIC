module real_aes_9799_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_1745;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1694;
wire n_1224;
wire n_1639;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1346;
wire n_552;
wire n_1383;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_1666;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1760;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_354;
wire n_1026;
wire n_1756;
wire n_492;
wire n_407;
wire n_1699;
wire n_419;
wire n_730;
wire n_1023;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1172;
wire n_459;
wire n_1689;
wire n_998;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1605;
wire n_1592;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1761;
wire n_1015;
wire n_1375;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1691;
wire n_640;
wire n_1721;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_317;
wire n_1595;
wire n_321;
wire n_1735;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1654;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_344;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_1352;
wire n_394;
wire n_729;
wire n_1323;
wire n_1280;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_1705;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
CKINVDCx5p33_ASAP7_75t_R g624 ( .A(n_0), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_1), .A2(n_281), .B1(n_529), .B2(n_530), .Y(n_528) );
INVx1_ASAP7_75t_L g582 ( .A(n_1), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g1440 ( .A1(n_2), .A2(n_303), .B1(n_1414), .B2(n_1422), .Y(n_1440) );
INVx1_ASAP7_75t_L g1188 ( .A(n_3), .Y(n_1188) );
AOI22xp33_ASAP7_75t_L g1213 ( .A1(n_3), .A2(n_123), .B1(n_1214), .B2(n_1215), .Y(n_1213) );
CKINVDCx5p33_ASAP7_75t_R g523 ( .A(n_4), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_5), .A2(n_181), .B1(n_839), .B2(n_840), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_5), .A2(n_181), .B1(n_855), .B2(n_857), .Y(n_854) );
AOI221xp5_ASAP7_75t_L g1155 ( .A1(n_6), .A2(n_174), .B1(n_562), .B2(n_1102), .C(n_1103), .Y(n_1155) );
OAI22xp33_ASAP7_75t_L g1160 ( .A1(n_6), .A2(n_276), .B1(n_504), .B2(n_1109), .Y(n_1160) );
AOI221xp5_ASAP7_75t_L g968 ( .A1(n_7), .A2(n_24), .B1(n_969), .B2(n_971), .C(n_973), .Y(n_968) );
INVx1_ASAP7_75t_L g1037 ( .A(n_7), .Y(n_1037) );
OAI22xp33_ASAP7_75t_L g410 ( .A1(n_8), .A2(n_85), .B1(n_411), .B2(n_413), .Y(n_410) );
AOI221xp5_ASAP7_75t_L g450 ( .A1(n_8), .A2(n_85), .B1(n_424), .B2(n_451), .C(n_453), .Y(n_450) );
AOI221xp5_ASAP7_75t_L g789 ( .A1(n_9), .A2(n_255), .B1(n_365), .B2(n_383), .C(n_650), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_9), .A2(n_255), .B1(n_532), .B2(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g919 ( .A(n_10), .Y(n_919) );
AOI22xp33_ASAP7_75t_SL g933 ( .A1(n_10), .A2(n_247), .B1(n_693), .B2(n_934), .Y(n_933) );
OAI22xp33_ASAP7_75t_L g1667 ( .A1(n_11), .A2(n_64), .B1(n_1668), .B2(n_1670), .Y(n_1667) );
OAI22xp33_ASAP7_75t_L g1676 ( .A1(n_11), .A2(n_160), .B1(n_327), .B2(n_665), .Y(n_1676) );
CKINVDCx20_ASAP7_75t_R g1079 ( .A(n_12), .Y(n_1079) );
AO22x2_ASAP7_75t_L g815 ( .A1(n_13), .A2(n_816), .B1(n_880), .B2(n_881), .Y(n_815) );
INVxp67_ASAP7_75t_SL g880 ( .A(n_13), .Y(n_880) );
AOI22xp5_ASAP7_75t_L g1441 ( .A1(n_13), .A2(n_260), .B1(n_1430), .B2(n_1436), .Y(n_1441) );
AOI21xp5_ASAP7_75t_L g1198 ( .A1(n_14), .A2(n_376), .B(n_377), .Y(n_1198) );
INVx1_ASAP7_75t_L g1201 ( .A(n_14), .Y(n_1201) );
XNOR2xp5_ASAP7_75t_L g1047 ( .A(n_15), .B(n_1048), .Y(n_1047) );
CKINVDCx16_ASAP7_75t_R g1468 ( .A(n_15), .Y(n_1468) );
INVx1_ASAP7_75t_L g1372 ( .A(n_16), .Y(n_1372) );
AOI22xp33_ASAP7_75t_L g1404 ( .A1(n_16), .A2(n_99), .B1(n_862), .B2(n_864), .Y(n_1404) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_17), .A2(n_309), .B1(n_866), .B2(n_1126), .Y(n_1125) );
INVxp67_ASAP7_75t_SL g1148 ( .A(n_17), .Y(n_1148) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_18), .A2(n_110), .B1(n_955), .B2(n_956), .Y(n_954) );
INVx1_ASAP7_75t_L g1001 ( .A(n_18), .Y(n_1001) );
INVx1_ASAP7_75t_L g1662 ( .A(n_19), .Y(n_1662) );
OAI222xp33_ASAP7_75t_L g1674 ( .A1(n_19), .A2(n_205), .B1(n_289), .B2(n_374), .C1(n_872), .C2(n_1675), .Y(n_1674) );
OAI222xp33_ASAP7_75t_L g608 ( .A1(n_20), .A2(n_62), .B1(n_127), .B2(n_609), .C1(n_614), .C2(n_617), .Y(n_608) );
INVx1_ASAP7_75t_L g651 ( .A(n_20), .Y(n_651) );
CKINVDCx5p33_ASAP7_75t_R g750 ( .A(n_21), .Y(n_750) );
CKINVDCx5p33_ASAP7_75t_R g960 ( .A(n_22), .Y(n_960) );
AOI22xp33_ASAP7_75t_SL g1287 ( .A1(n_23), .A2(n_108), .B1(n_530), .B2(n_537), .Y(n_1287) );
AOI22xp33_ASAP7_75t_L g1293 ( .A1(n_23), .A2(n_108), .B1(n_685), .B2(n_1153), .Y(n_1293) );
INVx1_ASAP7_75t_L g1031 ( .A(n_24), .Y(n_1031) );
AOI221xp5_ASAP7_75t_L g777 ( .A1(n_25), .A2(n_176), .B1(n_562), .B2(n_778), .C(n_779), .Y(n_777) );
INVx1_ASAP7_75t_L g808 ( .A(n_25), .Y(n_808) );
INVx1_ASAP7_75t_L g1274 ( .A(n_26), .Y(n_1274) );
AOI22xp33_ASAP7_75t_L g1291 ( .A1(n_26), .A2(n_292), .B1(n_650), .B2(n_1102), .Y(n_1291) );
CKINVDCx5p33_ASAP7_75t_R g895 ( .A(n_27), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_28), .A2(n_132), .B1(n_539), .B2(n_716), .Y(n_715) );
AOI22xp33_ASAP7_75t_SL g738 ( .A1(n_28), .A2(n_132), .B1(n_739), .B2(n_740), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_29), .A2(n_225), .B1(n_842), .B2(n_843), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_29), .A2(n_225), .B1(n_861), .B2(n_862), .Y(n_860) );
INVx1_ASAP7_75t_L g318 ( .A(n_30), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g1193 ( .A(n_31), .Y(n_1193) );
OAI22xp5_ASAP7_75t_L g1664 ( .A1(n_32), .A2(n_96), .B1(n_1665), .B2(n_1666), .Y(n_1664) );
AOI22xp33_ASAP7_75t_SL g1683 ( .A1(n_32), .A2(n_96), .B1(n_685), .B2(n_1290), .Y(n_1683) );
AOI21xp33_ASAP7_75t_L g1184 ( .A1(n_33), .A2(n_365), .B(n_383), .Y(n_1184) );
INVx1_ASAP7_75t_L g1211 ( .A(n_33), .Y(n_1211) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_34), .A2(n_137), .B1(n_775), .B2(n_776), .Y(n_774) );
INVx1_ASAP7_75t_L g809 ( .A(n_34), .Y(n_809) );
AOI22xp5_ASAP7_75t_L g1413 ( .A1(n_35), .A2(n_135), .B1(n_1414), .B2(n_1422), .Y(n_1413) );
AOI22xp33_ASAP7_75t_L g1454 ( .A1(n_36), .A2(n_196), .B1(n_1426), .B2(n_1455), .Y(n_1454) );
INVx1_ASAP7_75t_L g1226 ( .A(n_37), .Y(n_1226) );
AOI22xp33_ASAP7_75t_L g1259 ( .A1(n_37), .A2(n_191), .B1(n_1102), .B2(n_1254), .Y(n_1259) );
INVx1_ASAP7_75t_L g1321 ( .A(n_38), .Y(n_1321) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_38), .A2(n_249), .B1(n_846), .B2(n_849), .Y(n_1340) );
INVx1_ASAP7_75t_L g1678 ( .A(n_39), .Y(n_1678) );
AOI22xp33_ASAP7_75t_L g1693 ( .A1(n_39), .A2(n_203), .B1(n_866), .B2(n_1126), .Y(n_1693) );
AOI22xp33_ASAP7_75t_L g1253 ( .A1(n_40), .A2(n_128), .B1(n_560), .B2(n_1254), .Y(n_1253) );
AOI22xp33_ASAP7_75t_L g1262 ( .A1(n_40), .A2(n_128), .B1(n_424), .B2(n_693), .Y(n_1262) );
CKINVDCx5p33_ASAP7_75t_R g1192 ( .A(n_41), .Y(n_1192) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_42), .A2(n_213), .B1(n_532), .B2(n_533), .Y(n_531) );
INVx1_ASAP7_75t_L g573 ( .A(n_42), .Y(n_573) );
OAI222xp33_ASAP7_75t_L g1721 ( .A1(n_43), .A2(n_155), .B1(n_246), .B2(n_1722), .C1(n_1723), .C2(n_1724), .Y(n_1721) );
AOI221xp5_ASAP7_75t_L g1756 ( .A1(n_43), .A2(n_155), .B1(n_679), .B2(n_1757), .C(n_1759), .Y(n_1756) );
CKINVDCx5p33_ASAP7_75t_R g1382 ( .A(n_44), .Y(n_1382) );
AOI22xp5_ASAP7_75t_L g1434 ( .A1(n_45), .A2(n_113), .B1(n_1414), .B2(n_1422), .Y(n_1434) );
AO221x2_ASAP7_75t_L g1442 ( .A1(n_46), .A2(n_227), .B1(n_1430), .B2(n_1436), .C(n_1443), .Y(n_1442) );
CKINVDCx16_ASAP7_75t_R g1469 ( .A(n_47), .Y(n_1469) );
INVx1_ASAP7_75t_L g943 ( .A(n_48), .Y(n_943) );
AOI22xp5_ASAP7_75t_SL g1473 ( .A1(n_49), .A2(n_209), .B1(n_1426), .B2(n_1430), .Y(n_1473) );
INVx1_ASAP7_75t_L g1124 ( .A(n_50), .Y(n_1124) );
INVx1_ASAP7_75t_L g1282 ( .A(n_51), .Y(n_1282) );
AOI22xp33_ASAP7_75t_L g1289 ( .A1(n_51), .A2(n_158), .B1(n_677), .B2(n_1290), .Y(n_1289) );
INVx1_ASAP7_75t_L g1100 ( .A(n_52), .Y(n_1100) );
OAI22xp33_ASAP7_75t_L g1108 ( .A1(n_52), .A2(n_107), .B1(n_504), .B2(n_1109), .Y(n_1108) );
INVx1_ASAP7_75t_L g1333 ( .A(n_53), .Y(n_1333) );
AOI22xp33_ASAP7_75t_L g1351 ( .A1(n_53), .A2(n_241), .B1(n_866), .B2(n_1126), .Y(n_1351) );
INVx1_ASAP7_75t_L g1335 ( .A(n_54), .Y(n_1335) );
AOI22xp33_ASAP7_75t_L g1350 ( .A1(n_54), .A2(n_272), .B1(n_864), .B2(n_1349), .Y(n_1350) );
INVx1_ASAP7_75t_L g662 ( .A(n_55), .Y(n_662) );
AOI22xp33_ASAP7_75t_SL g700 ( .A1(n_55), .A2(n_95), .B1(n_424), .B2(n_701), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g1061 ( .A1(n_56), .A2(n_311), .B1(n_866), .B2(n_1062), .Y(n_1061) );
INVx1_ASAP7_75t_L g1086 ( .A(n_56), .Y(n_1086) );
CKINVDCx14_ASAP7_75t_R g1517 ( .A(n_57), .Y(n_1517) );
INVx1_ASAP7_75t_L g356 ( .A(n_58), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g423 ( .A1(n_58), .A2(n_219), .B1(n_424), .B2(n_430), .C(n_436), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g770 ( .A(n_59), .B(n_771), .Y(n_770) );
OAI22xp33_ASAP7_75t_L g890 ( .A1(n_60), .A2(n_278), .B1(n_588), .B2(n_589), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_60), .A2(n_278), .B1(n_724), .B2(n_937), .Y(n_936) );
INVx1_ASAP7_75t_L g1326 ( .A(n_61), .Y(n_1326) );
OAI22xp5_ASAP7_75t_L g1330 ( .A1(n_61), .A2(n_290), .B1(n_871), .B2(n_1303), .Y(n_1330) );
AOI22xp33_ASAP7_75t_SL g673 ( .A1(n_62), .A2(n_265), .B1(n_560), .B2(n_674), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g1251 ( .A1(n_63), .A2(n_171), .B1(n_677), .B2(n_1252), .Y(n_1251) );
AOI22xp33_ASAP7_75t_L g1261 ( .A1(n_63), .A2(n_171), .B1(n_703), .B2(n_862), .Y(n_1261) );
AOI22xp33_ASAP7_75t_L g1684 ( .A1(n_64), .A2(n_122), .B1(n_839), .B2(n_1254), .Y(n_1684) );
AOI22xp33_ASAP7_75t_L g1452 ( .A1(n_65), .A2(n_182), .B1(n_1414), .B2(n_1453), .Y(n_1452) );
CKINVDCx5p33_ASAP7_75t_R g516 ( .A(n_66), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g980 ( .A(n_67), .Y(n_980) );
AOI22xp33_ASAP7_75t_SL g1681 ( .A1(n_68), .A2(n_130), .B1(n_383), .B2(n_1254), .Y(n_1681) );
AOI22xp33_ASAP7_75t_L g1688 ( .A1(n_68), .A2(n_130), .B1(n_864), .B2(n_1689), .Y(n_1688) );
OAI22xp5_ASAP7_75t_L g961 ( .A1(n_69), .A2(n_216), .B1(n_962), .B2(n_965), .Y(n_961) );
OAI221xp5_ASAP7_75t_L g1013 ( .A1(n_69), .A2(n_216), .B1(n_1014), .B2(n_1018), .C(n_1020), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_70), .A2(n_304), .B1(n_451), .B2(n_533), .Y(n_535) );
OAI221xp5_ASAP7_75t_L g569 ( .A1(n_70), .A2(n_411), .B1(n_570), .B2(n_581), .C(n_586), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g1387 ( .A(n_71), .Y(n_1387) );
INVx1_ASAP7_75t_L g1227 ( .A(n_72), .Y(n_1227) );
AOI22xp33_ASAP7_75t_L g1257 ( .A1(n_72), .A2(n_149), .B1(n_677), .B2(n_1258), .Y(n_1257) );
CKINVDCx5p33_ASAP7_75t_R g1057 ( .A(n_73), .Y(n_1057) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_74), .A2(n_221), .B1(n_862), .B2(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g874 ( .A(n_74), .Y(n_874) );
INVx1_ASAP7_75t_L g826 ( .A(n_75), .Y(n_826) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_75), .A2(n_169), .B1(n_871), .B2(n_872), .Y(n_870) );
CKINVDCx14_ASAP7_75t_R g1444 ( .A(n_76), .Y(n_1444) );
CKINVDCx20_ASAP7_75t_R g1119 ( .A(n_77), .Y(n_1119) );
XNOR2x2_ASAP7_75t_L g339 ( .A(n_78), .B(n_340), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_79), .Y(n_382) );
BUFx2_ASAP7_75t_L g421 ( .A(n_80), .Y(n_421) );
BUFx2_ASAP7_75t_L g462 ( .A(n_80), .Y(n_462) );
INVx1_ASAP7_75t_L g476 ( .A(n_80), .Y(n_476) );
OR2x2_ASAP7_75t_L g996 ( .A(n_80), .B(n_396), .Y(n_996) );
AOI22xp33_ASAP7_75t_SL g1682 ( .A1(n_81), .A2(n_211), .B1(n_842), .B2(n_1290), .Y(n_1682) );
AOI22xp33_ASAP7_75t_L g1686 ( .A1(n_81), .A2(n_211), .B1(n_1218), .B2(n_1687), .Y(n_1686) );
INVx1_ASAP7_75t_L g1177 ( .A(n_82), .Y(n_1177) );
AOI22xp33_ASAP7_75t_L g1217 ( .A1(n_82), .A2(n_114), .B1(n_538), .B2(n_1218), .Y(n_1217) );
CKINVDCx5p33_ASAP7_75t_R g1385 ( .A(n_83), .Y(n_1385) );
AOI22xp33_ASAP7_75t_L g1286 ( .A1(n_84), .A2(n_300), .B1(n_424), .B2(n_693), .Y(n_1286) );
AOI22xp33_ASAP7_75t_SL g1294 ( .A1(n_84), .A2(n_300), .B1(n_674), .B2(n_1102), .Y(n_1294) );
CKINVDCx5p33_ASAP7_75t_R g1361 ( .A(n_86), .Y(n_1361) );
AOI22xp33_ASAP7_75t_L g1339 ( .A1(n_87), .A2(n_308), .B1(n_842), .B2(n_843), .Y(n_1339) );
AOI22xp33_ASAP7_75t_SL g1345 ( .A1(n_87), .A2(n_308), .B1(n_1346), .B2(n_1347), .Y(n_1345) );
OAI22xp5_ASAP7_75t_L g1276 ( .A1(n_88), .A2(n_138), .B1(n_617), .B2(n_1277), .Y(n_1276) );
OAI22xp33_ASAP7_75t_L g1302 ( .A1(n_88), .A2(n_138), .B1(n_653), .B2(n_1303), .Y(n_1302) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_89), .Y(n_354) );
INVx1_ASAP7_75t_L g519 ( .A(n_90), .Y(n_519) );
AOI221xp5_ASAP7_75t_L g557 ( .A1(n_90), .A2(n_251), .B1(n_558), .B2(n_560), .C(n_562), .Y(n_557) );
INVx1_ASAP7_75t_L g1323 ( .A(n_91), .Y(n_1323) );
AOI22xp33_ASAP7_75t_L g1341 ( .A1(n_91), .A2(n_103), .B1(n_648), .B2(n_1342), .Y(n_1341) );
AO221x1_ASAP7_75t_L g745 ( .A1(n_92), .A2(n_175), .B1(n_376), .B2(n_377), .C(n_675), .Y(n_745) );
INVx1_ASAP7_75t_L g760 ( .A(n_92), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g976 ( .A1(n_93), .A2(n_237), .B1(n_864), .B2(n_977), .Y(n_976) );
INVx1_ASAP7_75t_L g1038 ( .A(n_93), .Y(n_1038) );
INVx1_ASAP7_75t_L g643 ( .A(n_94), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_94), .A2(n_193), .B1(n_539), .B2(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g647 ( .A(n_95), .Y(n_647) );
XNOR2x2_ASAP7_75t_L g1313 ( .A(n_97), .B(n_1314), .Y(n_1313) );
AO22x2_ASAP7_75t_L g599 ( .A1(n_98), .A2(n_600), .B1(n_601), .B2(n_706), .Y(n_599) );
INVxp67_ASAP7_75t_SL g600 ( .A(n_98), .Y(n_600) );
INVx1_ASAP7_75t_L g1376 ( .A(n_99), .Y(n_1376) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_100), .A2(n_245), .B1(n_693), .B2(n_718), .Y(n_717) );
AOI221xp5_ASAP7_75t_L g741 ( .A1(n_100), .A2(n_245), .B1(n_365), .B2(n_383), .C(n_742), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_101), .A2(n_178), .B1(n_558), .B2(n_560), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_101), .A2(n_178), .B1(n_424), .B2(n_693), .Y(n_692) );
OAI22xp33_ASAP7_75t_L g1076 ( .A1(n_102), .A2(n_170), .B1(n_478), .B2(n_1077), .Y(n_1076) );
INVx1_ASAP7_75t_L g1106 ( .A(n_102), .Y(n_1106) );
INVx1_ASAP7_75t_L g1317 ( .A(n_103), .Y(n_1317) );
INVx1_ASAP7_75t_L g1151 ( .A(n_104), .Y(n_1151) );
OAI22xp33_ASAP7_75t_L g1161 ( .A1(n_104), .A2(n_174), .B1(n_1111), .B2(n_1113), .Y(n_1161) );
XNOR2xp5_ASAP7_75t_L g510 ( .A(n_105), .B(n_511), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_106), .A2(n_145), .B1(n_857), .B2(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g878 ( .A(n_106), .Y(n_878) );
AOI221xp5_ASAP7_75t_L g1101 ( .A1(n_107), .A2(n_262), .B1(n_377), .B2(n_1102), .C(n_1103), .Y(n_1101) );
CKINVDCx5p33_ASAP7_75t_R g902 ( .A(n_109), .Y(n_902) );
INVx1_ASAP7_75t_L g1011 ( .A(n_110), .Y(n_1011) );
OAI222xp33_ASAP7_75t_L g1726 ( .A1(n_111), .A2(n_166), .B1(n_299), .B2(n_1391), .C1(n_1727), .C2(n_1728), .Y(n_1726) );
INVx1_ASAP7_75t_L g1746 ( .A(n_111), .Y(n_1746) );
INVx1_ASAP7_75t_L g1130 ( .A(n_112), .Y(n_1130) );
OAI221xp5_ASAP7_75t_L g1143 ( .A1(n_112), .A2(n_411), .B1(n_586), .B2(n_1144), .C(n_1146), .Y(n_1143) );
INVx1_ASAP7_75t_L g1178 ( .A(n_114), .Y(n_1178) );
INVx1_ASAP7_75t_L g1242 ( .A(n_115), .Y(n_1242) );
AOI22xp33_ASAP7_75t_SL g1264 ( .A1(n_115), .A2(n_274), .B1(n_424), .B2(n_701), .Y(n_1264) );
AOI22xp33_ASAP7_75t_L g1298 ( .A1(n_116), .A2(n_140), .B1(n_539), .B2(n_716), .Y(n_1298) );
INVx1_ASAP7_75t_L g1305 ( .A(n_116), .Y(n_1305) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_117), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_118), .A2(n_173), .B1(n_537), .B2(n_539), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g587 ( .A1(n_118), .A2(n_173), .B1(n_588), .B2(n_589), .Y(n_587) );
INVx1_ASAP7_75t_L g915 ( .A(n_119), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_119), .A2(n_250), .B1(n_537), .B2(n_932), .Y(n_931) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_120), .Y(n_520) );
INVx1_ASAP7_75t_L g1096 ( .A(n_121), .Y(n_1096) );
OAI22xp33_ASAP7_75t_L g1110 ( .A1(n_121), .A2(n_262), .B1(n_1111), .B2(n_1113), .Y(n_1110) );
INVx1_ASAP7_75t_L g1659 ( .A(n_122), .Y(n_1659) );
INVx1_ASAP7_75t_L g1182 ( .A(n_123), .Y(n_1182) );
CKINVDCx5p33_ASAP7_75t_R g1197 ( .A(n_124), .Y(n_1197) );
AOI22xp5_ASAP7_75t_SL g1472 ( .A1(n_125), .A2(n_144), .B1(n_1414), .B2(n_1422), .Y(n_1472) );
AOI221xp5_ASAP7_75t_L g1713 ( .A1(n_126), .A2(n_273), .B1(n_975), .B2(n_1692), .C(n_1714), .Y(n_1713) );
INVx1_ASAP7_75t_L g1755 ( .A(n_126), .Y(n_1755) );
INVx1_ASAP7_75t_L g655 ( .A(n_127), .Y(n_655) );
INVx1_ASAP7_75t_L g1418 ( .A(n_129), .Y(n_1418) );
INVx1_ASAP7_75t_L g1237 ( .A(n_131), .Y(n_1237) );
AOI22xp33_ASAP7_75t_L g1265 ( .A1(n_131), .A2(n_168), .B1(n_495), .B2(n_862), .Y(n_1265) );
CKINVDCx16_ASAP7_75t_R g1465 ( .A(n_133), .Y(n_1465) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_134), .A2(n_268), .B1(n_775), .B2(n_791), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_134), .A2(n_268), .B1(n_438), .B2(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g924 ( .A(n_136), .Y(n_924) );
INVx1_ASAP7_75t_L g805 ( .A(n_137), .Y(n_805) );
INVx1_ASAP7_75t_L g1373 ( .A(n_139), .Y(n_1373) );
AOI221xp5_ASAP7_75t_L g1399 ( .A1(n_139), .A2(n_184), .B1(n_438), .B2(n_1400), .C(n_1402), .Y(n_1399) );
INVx1_ASAP7_75t_L g1306 ( .A(n_140), .Y(n_1306) );
INVx1_ASAP7_75t_L g1419 ( .A(n_141), .Y(n_1419) );
NAND2xp5_ASAP7_75t_L g1424 ( .A(n_141), .B(n_1417), .Y(n_1424) );
AOI221xp5_ASAP7_75t_L g1194 ( .A1(n_142), .A2(n_264), .B1(n_685), .B2(n_1195), .C(n_1196), .Y(n_1194) );
INVx1_ASAP7_75t_L g1204 ( .A(n_142), .Y(n_1204) );
INVx1_ASAP7_75t_L g821 ( .A(n_143), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_143), .A2(n_163), .B1(n_846), .B2(n_849), .Y(n_845) );
INVx1_ASAP7_75t_L g869 ( .A(n_145), .Y(n_869) );
INVx1_ASAP7_75t_L g1363 ( .A(n_146), .Y(n_1363) );
AOI21xp33_ASAP7_75t_L g1396 ( .A1(n_146), .A2(n_722), .B(n_1397), .Y(n_1396) );
INVx2_ASAP7_75t_L g330 ( .A(n_147), .Y(n_330) );
INVx1_ASAP7_75t_L g1364 ( .A(n_148), .Y(n_1364) );
AOI22xp33_ASAP7_75t_L g1395 ( .A1(n_148), .A2(n_201), .B1(n_803), .B2(n_970), .Y(n_1395) );
INVx1_ASAP7_75t_L g1230 ( .A(n_149), .Y(n_1230) );
OAI22xp5_ASAP7_75t_L g1138 ( .A1(n_150), .A2(n_180), .B1(n_1139), .B2(n_1140), .Y(n_1138) );
INVx1_ASAP7_75t_L g1157 ( .A(n_150), .Y(n_1157) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_151), .A2(n_234), .B1(n_685), .B2(n_686), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_151), .A2(n_234), .B1(n_529), .B2(n_539), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_152), .A2(n_305), .B1(n_862), .B2(n_1074), .Y(n_1073) );
OAI22xp5_ASAP7_75t_L g1081 ( .A1(n_152), .A2(n_305), .B1(n_588), .B2(n_589), .Y(n_1081) );
BUFx3_ASAP7_75t_L g428 ( .A(n_153), .Y(n_428) );
INVx1_ASAP7_75t_L g443 ( .A(n_153), .Y(n_443) );
INVx1_ASAP7_75t_L g788 ( .A(n_154), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_154), .A2(n_228), .B1(n_483), .B2(n_488), .Y(n_801) );
CKINVDCx5p33_ASAP7_75t_R g748 ( .A(n_156), .Y(n_748) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_157), .A2(n_284), .B1(n_398), .B2(n_404), .Y(n_397) );
INVx1_ASAP7_75t_L g460 ( .A(n_157), .Y(n_460) );
INVx1_ASAP7_75t_L g1283 ( .A(n_158), .Y(n_1283) );
OAI221xp5_ASAP7_75t_L g1231 ( .A1(n_159), .A2(n_218), .B1(n_617), .B2(n_1232), .C(n_1233), .Y(n_1231) );
INVx1_ASAP7_75t_L g1240 ( .A(n_159), .Y(n_1240) );
AOI22xp33_ASAP7_75t_L g1690 ( .A1(n_160), .A2(n_205), .B1(n_1691), .B2(n_1692), .Y(n_1690) );
INVx1_ASAP7_75t_L g1132 ( .A(n_161), .Y(n_1132) );
OAI211xp5_ASAP7_75t_SL g1149 ( .A1(n_161), .A2(n_413), .B(n_1150), .C(n_1156), .Y(n_1149) );
CKINVDCx5p33_ASAP7_75t_R g728 ( .A(n_162), .Y(n_728) );
INVx1_ASAP7_75t_L g833 ( .A(n_163), .Y(n_833) );
AOI22xp33_ASAP7_75t_SL g723 ( .A1(n_164), .A2(n_310), .B1(n_495), .B2(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g735 ( .A(n_164), .Y(n_735) );
AOI221xp5_ASAP7_75t_L g949 ( .A1(n_165), .A2(n_177), .B1(n_950), .B2(n_951), .C(n_952), .Y(n_949) );
INVx1_ASAP7_75t_L g1008 ( .A(n_165), .Y(n_1008) );
INVx1_ASAP7_75t_L g1737 ( .A(n_166), .Y(n_1737) );
AOI22xp33_ASAP7_75t_L g1712 ( .A1(n_167), .A2(n_261), .B1(n_1136), .B2(n_1346), .Y(n_1712) );
INVx1_ASAP7_75t_L g1744 ( .A(n_167), .Y(n_1744) );
INVx1_ASAP7_75t_L g1238 ( .A(n_168), .Y(n_1238) );
INVx1_ASAP7_75t_L g830 ( .A(n_169), .Y(n_830) );
INVx1_ASAP7_75t_L g1105 ( .A(n_170), .Y(n_1105) );
CKINVDCx5p33_ASAP7_75t_R g896 ( .A(n_172), .Y(n_896) );
INVx1_ASAP7_75t_L g762 ( .A(n_175), .Y(n_762) );
INVx1_ASAP7_75t_L g806 ( .A(n_176), .Y(n_806) );
INVx1_ASAP7_75t_L g1005 ( .A(n_177), .Y(n_1005) );
INVx1_ASAP7_75t_L g448 ( .A(n_179), .Y(n_448) );
INVx1_ASAP7_75t_L g474 ( .A(n_179), .Y(n_474) );
INVx1_ASAP7_75t_L g1158 ( .A(n_180), .Y(n_1158) );
CKINVDCx20_ASAP7_75t_R g1515 ( .A(n_183), .Y(n_1515) );
INVx1_ASAP7_75t_L g1375 ( .A(n_184), .Y(n_1375) );
INVx1_ASAP7_75t_L g785 ( .A(n_185), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_185), .A2(n_223), .B1(n_438), .B2(n_803), .Y(n_802) );
CKINVDCx5p33_ASAP7_75t_R g904 ( .A(n_186), .Y(n_904) );
XOR2x2_ASAP7_75t_L g887 ( .A(n_187), .B(n_888), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_188), .A2(n_288), .B1(n_424), .B2(n_720), .Y(n_719) );
OAI221xp5_ASAP7_75t_L g744 ( .A1(n_188), .A2(n_413), .B1(n_745), .B2(n_746), .C(n_749), .Y(n_744) );
CKINVDCx5p33_ASAP7_75t_R g1280 ( .A(n_189), .Y(n_1280) );
CKINVDCx5p33_ASAP7_75t_R g820 ( .A(n_190), .Y(n_820) );
INVx1_ASAP7_75t_L g1234 ( .A(n_191), .Y(n_1234) );
CKINVDCx5p33_ASAP7_75t_R g1174 ( .A(n_192), .Y(n_1174) );
INVx1_ASAP7_75t_L g640 ( .A(n_193), .Y(n_640) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_194), .Y(n_390) );
OAI221xp5_ASAP7_75t_L g465 ( .A1(n_194), .A2(n_466), .B1(n_477), .B2(n_478), .C(n_482), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g1380 ( .A(n_195), .Y(n_1380) );
CKINVDCx5p33_ASAP7_75t_R g1172 ( .A(n_197), .Y(n_1172) );
AOI221xp5_ASAP7_75t_L g1711 ( .A1(n_198), .A2(n_280), .B1(n_693), .B2(n_1349), .C(n_1397), .Y(n_1711) );
INVx1_ASAP7_75t_L g1742 ( .A(n_198), .Y(n_1742) );
CKINVDCx14_ASAP7_75t_R g1446 ( .A(n_199), .Y(n_1446) );
OAI22xp5_ASAP7_75t_L g781 ( .A1(n_200), .A2(n_214), .B1(n_568), .B2(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g812 ( .A(n_200), .Y(n_812) );
INVx1_ASAP7_75t_L g1359 ( .A(n_201), .Y(n_1359) );
INVx1_ASAP7_75t_L g813 ( .A(n_202), .Y(n_813) );
INVx1_ASAP7_75t_L g1679 ( .A(n_203), .Y(n_1679) );
CKINVDCx5p33_ASAP7_75t_R g900 ( .A(n_204), .Y(n_900) );
CKINVDCx5p33_ASAP7_75t_R g1229 ( .A(n_206), .Y(n_1229) );
CKINVDCx5p33_ASAP7_75t_R g1190 ( .A(n_207), .Y(n_1190) );
AOI22xp33_ASAP7_75t_L g1338 ( .A1(n_208), .A2(n_279), .B1(n_839), .B2(n_840), .Y(n_1338) );
AOI22xp33_ASAP7_75t_SL g1348 ( .A1(n_208), .A2(n_279), .B1(n_855), .B2(n_1349), .Y(n_1348) );
INVx1_ASAP7_75t_L g1072 ( .A(n_210), .Y(n_1072) );
OAI211xp5_ASAP7_75t_SL g1093 ( .A1(n_210), .A2(n_413), .B(n_1094), .C(n_1104), .Y(n_1093) );
INVx1_ASAP7_75t_L g1068 ( .A(n_212), .Y(n_1068) );
OAI221xp5_ASAP7_75t_L g1082 ( .A1(n_212), .A2(n_411), .B1(n_793), .B2(n_1083), .C(n_1091), .Y(n_1082) );
INVx1_ASAP7_75t_L g577 ( .A(n_213), .Y(n_577) );
INVx1_ASAP7_75t_L g811 ( .A(n_214), .Y(n_811) );
INVx1_ASAP7_75t_L g832 ( .A(n_215), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_215), .A2(n_301), .B1(n_839), .B2(n_840), .Y(n_850) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_217), .Y(n_373) );
INVx1_ASAP7_75t_L g1241 ( .A(n_218), .Y(n_1241) );
AOI21xp33_ASAP7_75t_L g361 ( .A1(n_219), .A2(n_362), .B(n_365), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g1056 ( .A(n_220), .Y(n_1056) );
INVx1_ASAP7_75t_L g876 ( .A(n_221), .Y(n_876) );
OAI221xp5_ASAP7_75t_L g891 ( .A1(n_222), .A2(n_413), .B1(n_892), .B2(n_898), .C(n_903), .Y(n_891) );
AOI22xp33_ASAP7_75t_SL g935 ( .A1(n_222), .A2(n_287), .B1(n_451), .B2(n_934), .Y(n_935) );
INVx1_ASAP7_75t_L g786 ( .A(n_223), .Y(n_786) );
INVx1_ASAP7_75t_L g992 ( .A(n_224), .Y(n_992) );
CKINVDCx5p33_ASAP7_75t_R g985 ( .A(n_226), .Y(n_985) );
AOI22xp33_ASAP7_75t_SL g1700 ( .A1(n_227), .A2(n_1701), .B1(n_1705), .B2(n_1761), .Y(n_1700) );
XNOR2x1_ASAP7_75t_L g1707 ( .A(n_227), .B(n_1708), .Y(n_1707) );
INVx1_ASAP7_75t_L g780 ( .A(n_228), .Y(n_780) );
CKINVDCx20_ASAP7_75t_R g1462 ( .A(n_229), .Y(n_1462) );
BUFx3_ASAP7_75t_L g429 ( .A(n_230), .Y(n_429) );
INVx1_ASAP7_75t_L g440 ( .A(n_230), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g1175 ( .A(n_231), .Y(n_1175) );
AO221x2_ASAP7_75t_L g1512 ( .A1(n_232), .A2(n_293), .B1(n_1455), .B2(n_1513), .C(n_1514), .Y(n_1512) );
CKINVDCx5p33_ASAP7_75t_R g727 ( .A(n_233), .Y(n_727) );
AO22x2_ASAP7_75t_L g1222 ( .A1(n_235), .A2(n_1223), .B1(n_1266), .B2(n_1267), .Y(n_1222) );
INVxp67_ASAP7_75t_L g1266 ( .A(n_235), .Y(n_1266) );
AOI22xp5_ASAP7_75t_L g1435 ( .A1(n_235), .A2(n_236), .B1(n_1430), .B2(n_1436), .Y(n_1435) );
INVx1_ASAP7_75t_L g1029 ( .A(n_237), .Y(n_1029) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_238), .Y(n_326) );
INVx1_ASAP7_75t_L g380 ( .A(n_238), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_238), .B(n_295), .Y(n_396) );
AND2x2_ASAP7_75t_L g400 ( .A(n_238), .B(n_367), .Y(n_400) );
CKINVDCx5p33_ASAP7_75t_R g747 ( .A(n_239), .Y(n_747) );
AOI21xp33_ASAP7_75t_L g375 ( .A1(n_240), .A2(n_376), .B(n_377), .Y(n_375) );
INVx1_ASAP7_75t_L g493 ( .A(n_240), .Y(n_493) );
INVx1_ASAP7_75t_L g1332 ( .A(n_241), .Y(n_1332) );
XNOR2xp5_ASAP7_75t_L g1270 ( .A(n_242), .B(n_1271), .Y(n_1270) );
INVx2_ASAP7_75t_L g449 ( .A(n_243), .Y(n_449) );
OR2x2_ASAP7_75t_L g492 ( .A(n_243), .B(n_474), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g989 ( .A(n_244), .Y(n_989) );
INVx1_ASAP7_75t_L g1760 ( .A(n_246), .Y(n_1760) );
INVx1_ASAP7_75t_L g922 ( .A(n_247), .Y(n_922) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_248), .Y(n_348) );
INVx1_ASAP7_75t_L g1318 ( .A(n_249), .Y(n_1318) );
INVx1_ASAP7_75t_L g911 ( .A(n_250), .Y(n_911) );
INVx1_ASAP7_75t_L g517 ( .A(n_251), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_252), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g1715 ( .A1(n_253), .A2(n_275), .B1(n_862), .B2(n_1716), .Y(n_1715) );
INVx1_ASAP7_75t_L g1753 ( .A(n_253), .Y(n_1753) );
INVx1_ASAP7_75t_L g1354 ( .A(n_254), .Y(n_1354) );
AOI22xp5_ASAP7_75t_SL g1425 ( .A1(n_254), .A2(n_258), .B1(n_1426), .B2(n_1430), .Y(n_1425) );
AOI22xp5_ASAP7_75t_L g1652 ( .A1(n_256), .A2(n_1653), .B1(n_1654), .B2(n_1694), .Y(n_1652) );
CKINVDCx5p33_ASAP7_75t_R g1653 ( .A(n_256), .Y(n_1653) );
INVx1_ASAP7_75t_L g631 ( .A(n_257), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_257), .A2(n_270), .B1(n_677), .B2(n_679), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g1296 ( .A1(n_259), .A2(n_283), .B1(n_424), .B2(n_1297), .Y(n_1296) );
INVx1_ASAP7_75t_L g1308 ( .A(n_259), .Y(n_1308) );
INVx1_ASAP7_75t_L g1740 ( .A(n_261), .Y(n_1740) );
AOI22x1_ASAP7_75t_L g708 ( .A1(n_263), .A2(n_709), .B1(n_710), .B2(n_763), .Y(n_708) );
INVxp67_ASAP7_75t_SL g763 ( .A(n_263), .Y(n_763) );
INVx1_ASAP7_75t_L g1202 ( .A(n_264), .Y(n_1202) );
INVx1_ASAP7_75t_L g620 ( .A(n_265), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g1133 ( .A1(n_266), .A2(n_296), .B1(n_1134), .B2(n_1136), .Y(n_1133) );
OAI22xp5_ASAP7_75t_L g1142 ( .A1(n_266), .A2(n_296), .B1(n_398), .B2(n_404), .Y(n_1142) );
INVx1_ASAP7_75t_L g1116 ( .A(n_267), .Y(n_1116) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_269), .Y(n_525) );
INVx1_ASAP7_75t_L g629 ( .A(n_270), .Y(n_629) );
CKINVDCx5p33_ASAP7_75t_R g1384 ( .A(n_271), .Y(n_1384) );
INVx1_ASAP7_75t_L g1329 ( .A(n_272), .Y(n_1329) );
AOI221xp5_ASAP7_75t_L g1751 ( .A1(n_273), .A2(n_275), .B1(n_677), .B2(n_1290), .C(n_1752), .Y(n_1751) );
INVx1_ASAP7_75t_L g1247 ( .A(n_274), .Y(n_1247) );
INVx1_ASAP7_75t_L g1154 ( .A(n_276), .Y(n_1154) );
CKINVDCx5p33_ASAP7_75t_R g1320 ( .A(n_277), .Y(n_1320) );
INVx1_ASAP7_75t_L g1750 ( .A(n_280), .Y(n_1750) );
INVx1_ASAP7_75t_L g583 ( .A(n_281), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g1720 ( .A(n_282), .Y(n_1720) );
INVx1_ASAP7_75t_L g1301 ( .A(n_283), .Y(n_1301) );
INVx1_ASAP7_75t_L g456 ( .A(n_284), .Y(n_456) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_285), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g1421 ( .A(n_285), .B(n_318), .Y(n_1421) );
AND3x2_ASAP7_75t_L g1429 ( .A(n_285), .B(n_318), .C(n_1418), .Y(n_1429) );
INVx2_ASAP7_75t_L g331 ( .A(n_286), .Y(n_331) );
OAI221xp5_ASAP7_75t_L g906 ( .A1(n_287), .A2(n_411), .B1(n_793), .B2(n_907), .C(n_916), .Y(n_906) );
INVx1_ASAP7_75t_L g743 ( .A(n_288), .Y(n_743) );
CKINVDCx5p33_ASAP7_75t_R g1661 ( .A(n_289), .Y(n_1661) );
INVx1_ASAP7_75t_L g1324 ( .A(n_290), .Y(n_1324) );
INVx1_ASAP7_75t_L g544 ( .A(n_291), .Y(n_544) );
INVx1_ASAP7_75t_L g1279 ( .A(n_292), .Y(n_1279) );
OAI221xp5_ASAP7_75t_L g1366 ( .A1(n_294), .A2(n_297), .B1(n_1014), .B2(n_1018), .C(n_1367), .Y(n_1366) );
OAI221xp5_ASAP7_75t_L g1390 ( .A1(n_294), .A2(n_297), .B1(n_965), .B2(n_1391), .C(n_1393), .Y(n_1390) );
INVx1_ASAP7_75t_L g333 ( .A(n_295), .Y(n_333) );
INVx2_ASAP7_75t_L g367 ( .A(n_295), .Y(n_367) );
AO22x2_ASAP7_75t_L g1168 ( .A1(n_298), .A2(n_1169), .B1(n_1219), .B2(n_1220), .Y(n_1168) );
INVxp67_ASAP7_75t_SL g1219 ( .A(n_298), .Y(n_1219) );
INVx1_ASAP7_75t_L g1735 ( .A(n_299), .Y(n_1735) );
INVx1_ASAP7_75t_L g823 ( .A(n_301), .Y(n_823) );
INVx1_ASAP7_75t_L g388 ( .A(n_302), .Y(n_388) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_302), .Y(n_477) );
OAI211xp5_ASAP7_75t_SL g550 ( .A1(n_304), .A2(n_413), .B(n_551), .C(n_564), .Y(n_550) );
INVx1_ASAP7_75t_L g1123 ( .A(n_306), .Y(n_1123) );
CKINVDCx5p33_ASAP7_75t_R g905 ( .A(n_307), .Y(n_905) );
INVxp33_ASAP7_75t_SL g1147 ( .A(n_309), .Y(n_1147) );
INVx1_ASAP7_75t_L g736 ( .A(n_310), .Y(n_736) );
INVx1_ASAP7_75t_L g1090 ( .A(n_311), .Y(n_1090) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_334), .B(n_1406), .Y(n_312) );
INVx2_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_316), .B(n_321), .Y(n_315) );
AND2x4_ASAP7_75t_L g1704 ( .A(n_316), .B(n_322), .Y(n_1704) );
NOR2xp33_ASAP7_75t_SL g316 ( .A(n_317), .B(n_319), .Y(n_316) );
INVx1_ASAP7_75t_SL g1699 ( .A(n_317), .Y(n_1699) );
NAND2xp5_ASAP7_75t_L g1767 ( .A(n_317), .B(n_319), .Y(n_1767) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g1698 ( .A(n_319), .B(n_1699), .Y(n_1698) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_327), .Y(n_322) );
INVxp67_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OR2x6_ASAP7_75t_L g670 ( .A(n_324), .B(n_462), .Y(n_670) );
OR2x2_ASAP7_75t_L g879 ( .A(n_324), .B(n_462), .Y(n_879) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g580 ( .A(n_325), .B(n_333), .Y(n_580) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g365 ( .A(n_326), .B(n_366), .Y(n_365) );
INVx8_ASAP7_75t_L g663 ( .A(n_327), .Y(n_663) );
OR2x6_ASAP7_75t_L g327 ( .A(n_328), .B(n_332), .Y(n_327) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_328), .Y(n_576) );
OR2x6_ASAP7_75t_L g665 ( .A(n_328), .B(n_642), .Y(n_665) );
OR2x2_ASAP7_75t_L g995 ( .A(n_328), .B(n_996), .Y(n_995) );
INVx1_ASAP7_75t_L g1028 ( .A(n_328), .Y(n_1028) );
INVx2_ASAP7_75t_SL g1043 ( .A(n_328), .Y(n_1043) );
INVx2_ASAP7_75t_SL g1371 ( .A(n_328), .Y(n_1371) );
BUFx2_ASAP7_75t_L g1754 ( .A(n_328), .Y(n_1754) );
OAI22xp33_ASAP7_75t_L g1759 ( .A1(n_328), .A2(n_752), .B1(n_1720), .B2(n_1760), .Y(n_1759) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx2_ASAP7_75t_L g347 ( .A(n_330), .Y(n_347) );
AND2x4_ASAP7_75t_L g352 ( .A(n_330), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g360 ( .A(n_330), .Y(n_360) );
AND2x2_ASAP7_75t_L g364 ( .A(n_330), .B(n_331), .Y(n_364) );
INVx1_ASAP7_75t_L g417 ( .A(n_330), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_331), .B(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g353 ( .A(n_331), .Y(n_353) );
INVx1_ASAP7_75t_L g359 ( .A(n_331), .Y(n_359) );
INVx1_ASAP7_75t_L g389 ( .A(n_331), .Y(n_389) );
INVx1_ASAP7_75t_L g403 ( .A(n_331), .Y(n_403) );
AND2x4_ASAP7_75t_L g654 ( .A(n_332), .B(n_389), .Y(n_654) );
INVx2_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g872 ( .A(n_333), .B(n_658), .Y(n_872) );
OR2x2_ASAP7_75t_L g1303 ( .A(n_333), .B(n_658), .Y(n_1303) );
XNOR2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_1163), .Y(n_334) );
XOR2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_764), .Y(n_335) );
XOR2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_596), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_339), .B1(n_509), .B2(n_593), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND4xp25_ASAP7_75t_L g340 ( .A(n_341), .B(n_422), .C(n_486), .D(n_499), .Y(n_340) );
OAI31xp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_397), .A3(n_410), .B(n_418), .Y(n_341) );
OAI221xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_355), .B1(n_368), .B2(n_372), .C(n_381), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_348), .B1(n_349), .B2(n_354), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_344), .A2(n_369), .B1(n_370), .B2(n_371), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_344), .A2(n_582), .B1(n_583), .B2(n_584), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_344), .A2(n_370), .B1(n_747), .B2(n_748), .Y(n_746) );
BUFx2_ASAP7_75t_L g899 ( .A(n_344), .Y(n_899) );
OAI22xp5_ASAP7_75t_L g1146 ( .A1(n_344), .A2(n_844), .B1(n_1147), .B2(n_1148), .Y(n_1146) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g553 ( .A(n_345), .Y(n_553) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g910 ( .A(n_346), .Y(n_910) );
BUFx2_ASAP7_75t_L g1187 ( .A(n_346), .Y(n_1187) );
INVx1_ASAP7_75t_L g392 ( .A(n_347), .Y(n_392) );
AND2x4_ASAP7_75t_L g401 ( .A(n_347), .B(n_402), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g436 ( .A1(n_348), .A2(n_354), .B1(n_437), .B2(n_441), .Y(n_436) );
INVx2_ASAP7_75t_SL g1252 ( .A(n_349), .Y(n_1252) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g370 ( .A(n_350), .Y(n_370) );
INVx2_ASAP7_75t_L g680 ( .A(n_350), .Y(n_680) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_350), .Y(n_776) );
INVx1_ASAP7_75t_L g1089 ( .A(n_350), .Y(n_1089) );
INVx3_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx3_ASAP7_75t_L g688 ( .A(n_351), .Y(n_688) );
BUFx6f_ASAP7_75t_L g914 ( .A(n_351), .Y(n_914) );
INVx3_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g409 ( .A(n_352), .Y(n_409) );
INVx1_ASAP7_75t_L g585 ( .A(n_352), .Y(n_585) );
BUFx6f_ASAP7_75t_L g740 ( .A(n_352), .Y(n_740) );
AND2x4_ASAP7_75t_L g416 ( .A(n_353), .B(n_417), .Y(n_416) );
OAI21xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_357), .B(n_361), .Y(n_355) );
INVx3_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g374 ( .A(n_358), .Y(n_374) );
INVx2_ASAP7_75t_L g386 ( .A(n_358), .Y(n_386) );
BUFx2_ASAP7_75t_L g572 ( .A(n_358), .Y(n_572) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_359), .B(n_360), .Y(n_753) );
INVx1_ASAP7_75t_L g658 ( .A(n_360), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_362), .B(n_548), .Y(n_547) );
BUFx2_ASAP7_75t_L g1102 ( .A(n_362), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1749 ( .A(n_362), .B(n_1004), .Y(n_1749) );
INVx2_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g376 ( .A(n_363), .Y(n_376) );
INVx2_ASAP7_75t_SL g1010 ( .A(n_363), .Y(n_1010) );
INVx3_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_364), .Y(n_384) );
OR2x6_ASAP7_75t_L g1025 ( .A(n_365), .B(n_421), .Y(n_1025) );
INVx1_ASAP7_75t_L g642 ( .A(n_366), .Y(n_642) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g379 ( .A(n_367), .Y(n_379) );
AOI222xp33_ASAP7_75t_L g486 ( .A1(n_369), .A2(n_382), .B1(n_487), .B2(n_493), .C1(n_494), .C2(n_497), .Y(n_486) );
INVx2_ASAP7_75t_L g1290 ( .A(n_370), .Y(n_1290) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_371), .A2(n_373), .B1(n_500), .B2(n_503), .Y(n_499) );
OAI21xp33_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_374), .B(n_375), .Y(n_372) );
OAI221xp5_ASAP7_75t_L g1091 ( .A1(n_374), .A2(n_578), .B1(n_1056), .B2(n_1057), .C(n_1092), .Y(n_1091) );
OAI21xp5_ASAP7_75t_SL g1196 ( .A1(n_374), .A2(n_1197), .B(n_1198), .Y(n_1196) );
BUFx3_ASAP7_75t_L g839 ( .A(n_376), .Y(n_839) );
BUFx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g563 ( .A(n_378), .Y(n_563) );
OR2x6_ASAP7_75t_L g682 ( .A(n_378), .B(n_475), .Y(n_682) );
NAND2x1p5_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
INVx1_ASAP7_75t_L g660 ( .A(n_379), .Y(n_660) );
A2O1A1Ixp33_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_383), .B(n_385), .C(n_393), .Y(n_381) );
INVx1_ASAP7_75t_L g1343 ( .A(n_383), .Y(n_1343) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x4_ASAP7_75t_L g412 ( .A(n_384), .B(n_400), .Y(n_412) );
INVx3_ASAP7_75t_L g561 ( .A(n_384), .Y(n_561) );
BUFx2_ASAP7_75t_L g778 ( .A(n_384), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
OR2x2_ASAP7_75t_L g586 ( .A(n_386), .B(n_394), .Y(n_586) );
OR2x6_ASAP7_75t_L g793 ( .A(n_386), .B(n_394), .Y(n_793) );
INVx1_ASAP7_75t_L g918 ( .A(n_386), .Y(n_918) );
AOI22xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_389), .B1(n_390), .B2(n_391), .Y(n_387) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_389), .Y(n_566) );
INVx1_ASAP7_75t_L g756 ( .A(n_389), .Y(n_756) );
NAND2x1p5_ASAP7_75t_L g1019 ( .A(n_391), .B(n_1017), .Y(n_1019) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OR2x6_ASAP7_75t_L g568 ( .A(n_392), .B(n_394), .Y(n_568) );
A2O1A1Ixp33_ASAP7_75t_L g749 ( .A1(n_393), .A2(n_560), .B(n_750), .C(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g548 ( .A(n_394), .Y(n_548) );
INVx1_ASAP7_75t_L g783 ( .A(n_394), .Y(n_783) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx3_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx3_ASAP7_75t_L g588 ( .A(n_399), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_399), .A2(n_405), .B1(n_735), .B2(n_736), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_399), .A2(n_405), .B1(n_785), .B2(n_786), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g1176 ( .A1(n_399), .A2(n_405), .B1(n_1177), .B2(n_1178), .Y(n_1176) );
AND2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
INVx2_ASAP7_75t_L g407 ( .A(n_400), .Y(n_407) );
AND2x4_ASAP7_75t_L g1004 ( .A(n_400), .B(n_476), .Y(n_1004) );
AND2x4_ASAP7_75t_L g641 ( .A(n_401), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g678 ( .A(n_401), .Y(n_678) );
BUFx2_ASAP7_75t_L g685 ( .A(n_401), .Y(n_685) );
BUFx6f_ASAP7_75t_L g739 ( .A(n_401), .Y(n_739) );
BUFx6f_ASAP7_75t_L g775 ( .A(n_401), .Y(n_775) );
BUFx2_ASAP7_75t_L g842 ( .A(n_401), .Y(n_842) );
BUFx6f_ASAP7_75t_L g848 ( .A(n_401), .Y(n_848) );
INVx1_ASAP7_75t_L g1758 ( .A(n_401), .Y(n_1758) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx3_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx3_ASAP7_75t_L g589 ( .A(n_405), .Y(n_589) );
AND2x4_ASAP7_75t_L g405 ( .A(n_406), .B(n_408), .Y(n_405) );
AND2x4_ASAP7_75t_L g414 ( .A(n_406), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g556 ( .A(n_408), .Y(n_556) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g791 ( .A(n_409), .Y(n_791) );
CKINVDCx6p67_ASAP7_75t_R g411 ( .A(n_412), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_412), .A2(n_738), .B1(n_741), .B2(n_743), .Y(n_737) );
AOI221xp5_ASAP7_75t_L g787 ( .A1(n_412), .A2(n_788), .B1(n_789), .B2(n_790), .C(n_792), .Y(n_787) );
AOI222xp33_ASAP7_75t_L g1171 ( .A1(n_412), .A2(n_414), .B1(n_1172), .B2(n_1173), .C1(n_1174), .C2(n_1175), .Y(n_1171) );
INVx8_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AOI221xp5_ASAP7_75t_SL g773 ( .A1(n_414), .A2(n_774), .B1(n_777), .B2(n_780), .C(n_781), .Y(n_773) );
INVx1_ASAP7_75t_L g559 ( .A(n_415), .Y(n_559) );
BUFx3_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx6f_ASAP7_75t_L g650 ( .A(n_416), .Y(n_650) );
AND2x4_ASAP7_75t_L g667 ( .A(n_416), .B(n_668), .Y(n_667) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_416), .Y(n_675) );
BUFx3_ASAP7_75t_L g742 ( .A(n_416), .Y(n_742) );
BUFx2_ASAP7_75t_L g1245 ( .A(n_416), .Y(n_1245) );
INVx1_ASAP7_75t_L g794 ( .A(n_418), .Y(n_794) );
OAI31xp33_ASAP7_75t_L g1141 ( .A1(n_418), .A2(n_1142), .A3(n_1143), .B(n_1149), .Y(n_1141) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NOR2xp67_ASAP7_75t_L g546 ( .A(n_419), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OR2x6_ASAP7_75t_L g445 ( .A(n_420), .B(n_446), .Y(n_445) );
BUFx2_ASAP7_75t_L g592 ( .A(n_420), .Y(n_592) );
AND2x4_ASAP7_75t_L g690 ( .A(n_420), .B(n_580), .Y(n_690) );
OR2x2_ASAP7_75t_L g697 ( .A(n_420), .B(n_698), .Y(n_697) );
OR2x2_ASAP7_75t_L g714 ( .A(n_420), .B(n_446), .Y(n_714) );
AND2x4_ASAP7_75t_L g837 ( .A(n_420), .B(n_580), .Y(n_837) );
OAI31xp33_ASAP7_75t_L g889 ( .A1(n_420), .A2(n_890), .A3(n_891), .B(n_906), .Y(n_889) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx2_ASAP7_75t_L g637 ( .A(n_421), .Y(n_637) );
AOI221xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_444), .B1(n_450), .B2(n_461), .C(n_465), .Y(n_422) );
INVx3_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g800 ( .A(n_425), .Y(n_800) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND2x4_ASAP7_75t_L g604 ( .A(n_426), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g731 ( .A(n_426), .Y(n_731) );
BUFx6f_ASAP7_75t_L g825 ( .A(n_426), .Y(n_825) );
BUFx6f_ASAP7_75t_L g859 ( .A(n_426), .Y(n_859) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_427), .Y(n_484) );
AND2x2_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
INVx2_ASAP7_75t_L g434 ( .A(n_428), .Y(n_434) );
AND2x4_ASAP7_75t_L g439 ( .A(n_428), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g435 ( .A(n_429), .Y(n_435) );
AND2x4_ASAP7_75t_L g442 ( .A(n_429), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g1716 ( .A(n_431), .Y(n_1716) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_432), .Y(n_452) );
INVx2_ASAP7_75t_L g623 ( .A(n_432), .Y(n_623) );
INVx2_ASAP7_75t_L g694 ( .A(n_432), .Y(n_694) );
INVx1_ASAP7_75t_L g701 ( .A(n_432), .Y(n_701) );
INVx2_ASAP7_75t_SL g722 ( .A(n_432), .Y(n_722) );
INVx2_ASAP7_75t_L g856 ( .A(n_432), .Y(n_856) );
INVx6_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g489 ( .A(n_433), .Y(n_489) );
AND2x2_ASAP7_75t_L g498 ( .A(n_433), .B(n_472), .Y(n_498) );
BUFx2_ASAP7_75t_L g532 ( .A(n_433), .Y(n_532) );
AND2x4_ASAP7_75t_L g625 ( .A(n_433), .B(n_626), .Y(n_625) );
AND2x4_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
INVx1_ASAP7_75t_L g481 ( .A(n_434), .Y(n_481) );
INVx1_ASAP7_75t_L g469 ( .A(n_435), .Y(n_469) );
INVx1_ASAP7_75t_L g955 ( .A(n_437), .Y(n_955) );
INVx1_ASAP7_75t_L g1687 ( .A(n_437), .Y(n_1687) );
INVx2_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
BUFx3_ASAP7_75t_L g861 ( .A(n_438), .Y(n_861) );
AND2x4_ASAP7_75t_L g958 ( .A(n_438), .B(n_959), .Y(n_958) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_439), .Y(n_455) );
INVx2_ASAP7_75t_SL g496 ( .A(n_439), .Y(n_496) );
BUFx2_ASAP7_75t_L g529 ( .A(n_439), .Y(n_529) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_439), .Y(n_538) );
AND2x6_ASAP7_75t_L g630 ( .A(n_439), .B(n_606), .Y(n_630) );
BUFx2_ASAP7_75t_L g703 ( .A(n_439), .Y(n_703) );
BUFx6f_ASAP7_75t_L g970 ( .A(n_439), .Y(n_970) );
BUFx3_ASAP7_75t_L g1135 ( .A(n_439), .Y(n_1135) );
HB1xp67_ASAP7_75t_L g1714 ( .A(n_439), .Y(n_1714) );
INVx1_ASAP7_75t_L g508 ( .A(n_440), .Y(n_508) );
INVx1_ASAP7_75t_L g1126 ( .A(n_441), .Y(n_1126) );
INVx1_ASAP7_75t_L g1218 ( .A(n_441), .Y(n_1218) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g459 ( .A(n_442), .Y(n_459) );
INVx1_ASAP7_75t_L g502 ( .A(n_442), .Y(n_502) );
BUFx6f_ASAP7_75t_L g633 ( .A(n_442), .Y(n_633) );
BUFx6f_ASAP7_75t_L g803 ( .A(n_442), .Y(n_803) );
INVx1_ASAP7_75t_L g507 ( .A(n_443), .Y(n_507) );
AOI33xp33_ASAP7_75t_L g527 ( .A1(n_444), .A2(n_528), .A3(n_531), .B1(n_535), .B2(n_536), .B3(n_540), .Y(n_527) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g853 ( .A(n_445), .Y(n_853) );
CKINVDCx5p33_ASAP7_75t_R g930 ( .A(n_445), .Y(n_930) );
OAI22xp5_ASAP7_75t_SL g1051 ( .A1(n_445), .A2(n_1052), .B1(n_1064), .B2(n_1065), .Y(n_1051) );
OAI22xp5_ASAP7_75t_SL g1121 ( .A1(n_445), .A2(n_1122), .B1(n_1127), .B2(n_1129), .Y(n_1121) );
OAI22xp5_ASAP7_75t_L g1209 ( .A1(n_445), .A2(n_1127), .B1(n_1210), .B2(n_1216), .Y(n_1209) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g698 ( .A(n_447), .Y(n_698) );
INVx2_ASAP7_75t_SL g975 ( .A(n_447), .Y(n_975) );
BUFx3_ASAP7_75t_L g1403 ( .A(n_447), .Y(n_1403) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
AND2x4_ASAP7_75t_L g463 ( .A(n_448), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g636 ( .A(n_448), .Y(n_636) );
INVx2_ASAP7_75t_L g464 ( .A(n_449), .Y(n_464) );
INVx1_ASAP7_75t_L g607 ( .A(n_449), .Y(n_607) );
INVx1_ASAP7_75t_L g611 ( .A(n_449), .Y(n_611) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_449), .Y(n_627) );
INVx4_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g951 ( .A(n_452), .Y(n_951) );
INVx2_ASAP7_75t_L g1297 ( .A(n_452), .Y(n_1297) );
OAI22xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_456), .B1(n_457), .B2(n_460), .Y(n_453) );
INVx1_ASAP7_75t_L g937 ( .A(n_454), .Y(n_937) );
INVx1_ASAP7_75t_L g1214 ( .A(n_454), .Y(n_1214) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g530 ( .A(n_457), .Y(n_530) );
INVx1_ASAP7_75t_L g539 ( .A(n_457), .Y(n_539) );
INVx2_ASAP7_75t_SL g932 ( .A(n_457), .Y(n_932) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_L g957 ( .A(n_458), .Y(n_957) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g991 ( .A(n_459), .B(n_492), .Y(n_991) );
AOI33xp33_ASAP7_75t_L g852 ( .A1(n_461), .A2(n_853), .A3(n_854), .B1(n_860), .B2(n_863), .B3(n_865), .Y(n_852) );
INVx4_ASAP7_75t_L g1064 ( .A(n_461), .Y(n_1064) );
BUFx4f_ASAP7_75t_L g1128 ( .A(n_461), .Y(n_1128) );
BUFx4f_ASAP7_75t_L g1352 ( .A(n_461), .Y(n_1352) );
AOI33xp33_ASAP7_75t_L g1685 ( .A1(n_461), .A2(n_853), .A3(n_1686), .B1(n_1688), .B2(n_1690), .B3(n_1693), .Y(n_1685) );
AND2x4_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
AND2x4_ASAP7_75t_L g497 ( .A(n_462), .B(n_498), .Y(n_497) );
AND2x4_ASAP7_75t_L g540 ( .A(n_462), .B(n_463), .Y(n_540) );
INVx2_ASAP7_75t_L g953 ( .A(n_463), .Y(n_953) );
CKINVDCx5p33_ASAP7_75t_R g1397 ( .A(n_463), .Y(n_1397) );
AND2x4_ASAP7_75t_L g472 ( .A(n_464), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g524 ( .A(n_466), .Y(n_524) );
INVx2_ASAP7_75t_L g726 ( .A(n_466), .Y(n_726) );
INVx1_ASAP7_75t_L g928 ( .A(n_466), .Y(n_928) );
HB1xp67_ASAP7_75t_L g1077 ( .A(n_466), .Y(n_1077) );
NAND2x1p5_ASAP7_75t_L g466 ( .A(n_467), .B(n_470), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g964 ( .A(n_468), .Y(n_964) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g613 ( .A(n_469), .Y(n_613) );
INVx2_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
OR2x6_ASAP7_75t_L g478 ( .A(n_471), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g485 ( .A(n_471), .Y(n_485) );
OR2x2_ASAP7_75t_L g1140 ( .A(n_471), .B(n_479), .Y(n_1140) );
NAND2x1p5_ASAP7_75t_L g471 ( .A(n_472), .B(n_475), .Y(n_471) );
AND2x4_ASAP7_75t_L g963 ( .A(n_472), .B(n_964), .Y(n_963) );
AND2x2_ASAP7_75t_L g966 ( .A(n_472), .B(n_480), .Y(n_966) );
INVx1_ASAP7_75t_L g983 ( .A(n_472), .Y(n_983) );
AND2x4_ASAP7_75t_L g1392 ( .A(n_472), .B(n_964), .Y(n_1392) );
BUFx2_ASAP7_75t_L g1718 ( .A(n_472), .Y(n_1718) );
AND2x4_ASAP7_75t_L g1729 ( .A(n_472), .B(n_480), .Y(n_1729) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OR2x2_ASAP7_75t_L g491 ( .A(n_476), .B(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g526 ( .A(n_478), .Y(n_526) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
BUFx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND2x6_ASAP7_75t_L g618 ( .A(n_481), .B(n_607), .Y(n_618) );
INVx1_ASAP7_75t_L g542 ( .A(n_482), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_485), .Y(n_482) );
HB1xp67_ASAP7_75t_L g1215 ( .A(n_483), .Y(n_1215) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_SL g534 ( .A(n_484), .Y(n_534) );
BUFx4f_ASAP7_75t_L g718 ( .A(n_484), .Y(n_718) );
AND2x4_ASAP7_75t_L g979 ( .A(n_484), .B(n_959), .Y(n_979) );
INVx1_ASAP7_75t_L g1207 ( .A(n_484), .Y(n_1207) );
BUFx3_ASAP7_75t_L g1689 ( .A(n_484), .Y(n_1689) );
AND2x4_ASAP7_75t_L g1717 ( .A(n_484), .B(n_1718), .Y(n_1717) );
AND2x2_ASAP7_75t_L g729 ( .A(n_485), .B(n_730), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_487), .A2(n_494), .B1(n_519), .B2(n_520), .Y(n_518) );
AOI222xp33_ASAP7_75t_L g759 ( .A1(n_487), .A2(n_497), .B1(n_500), .B2(n_747), .C1(n_750), .C2(n_760), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g807 ( .A1(n_487), .A2(n_494), .B1(n_808), .B2(n_809), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_487), .A2(n_494), .B1(n_896), .B2(n_900), .Y(n_940) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_490), .Y(n_487) );
INVx2_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g864 ( .A(n_489), .Y(n_864) );
AND2x2_ASAP7_75t_L g494 ( .A(n_490), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OR2x6_ASAP7_75t_L g501 ( .A(n_491), .B(n_502), .Y(n_501) );
OR2x6_ASAP7_75t_L g504 ( .A(n_491), .B(n_505), .Y(n_504) );
OR2x2_ASAP7_75t_L g1109 ( .A(n_491), .B(n_502), .Y(n_1109) );
OR2x2_ASAP7_75t_L g1111 ( .A(n_491), .B(n_1112), .Y(n_1111) );
OR2x2_ASAP7_75t_L g1113 ( .A(n_491), .B(n_1114), .Y(n_1113) );
INVx2_ASAP7_75t_L g959 ( .A(n_492), .Y(n_959) );
OR2x2_ASAP7_75t_L g987 ( .A(n_492), .B(n_988), .Y(n_987) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_494), .A2(n_503), .B1(n_748), .B2(n_762), .Y(n_761) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g716 ( .A(n_496), .Y(n_716) );
OR2x6_ASAP7_75t_L g545 ( .A(n_497), .B(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g997 ( .A(n_497), .Y(n_997) );
INVx2_ASAP7_75t_L g1727 ( .A(n_498), .Y(n_1727) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_500), .A2(n_503), .B1(n_516), .B2(n_517), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g804 ( .A1(n_500), .A2(n_503), .B1(n_805), .B2(n_806), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_500), .A2(n_503), .B1(n_895), .B2(n_902), .Y(n_939) );
CKINVDCx6p67_ASAP7_75t_R g500 ( .A(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g798 ( .A(n_502), .Y(n_798) );
CKINVDCx6p67_ASAP7_75t_R g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g616 ( .A(n_506), .Y(n_616) );
BUFx4f_ASAP7_75t_L g1060 ( .A(n_506), .Y(n_1060) );
INVx1_ASAP7_75t_L g1071 ( .A(n_506), .Y(n_1071) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
OR2x2_ASAP7_75t_L g988 ( .A(n_507), .B(n_508), .Y(n_988) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g595 ( .A(n_510), .Y(n_595) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NAND3xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_543), .C(n_549), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_521), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_518), .Y(n_514) );
OAI221xp5_ASAP7_75t_L g551 ( .A1(n_516), .A2(n_520), .B1(n_552), .B2(n_554), .C(n_557), .Y(n_551) );
NAND3xp33_ASAP7_75t_L g521 ( .A(n_522), .B(n_527), .C(n_541), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_524), .B1(n_525), .B2(n_526), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_523), .A2(n_525), .B1(n_565), .B2(n_567), .Y(n_564) );
INVx1_ASAP7_75t_L g1139 ( .A(n_524), .Y(n_1139) );
AOI221xp5_ASAP7_75t_L g725 ( .A1(n_526), .A2(n_726), .B1(n_727), .B2(n_728), .C(n_729), .Y(n_725) );
AOI221xp5_ASAP7_75t_L g810 ( .A1(n_526), .A2(n_726), .B1(n_729), .B2(n_811), .C(n_812), .Y(n_810) );
AOI22xp5_ASAP7_75t_L g927 ( .A1(n_526), .A2(n_904), .B1(n_905), .B2(n_928), .Y(n_927) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g934 ( .A(n_534), .Y(n_934) );
INVx2_ASAP7_75t_L g1349 ( .A(n_534), .Y(n_1349) );
BUFx4f_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
BUFx2_ASAP7_75t_L g866 ( .A(n_538), .Y(n_866) );
INVx1_ASAP7_75t_L g1114 ( .A(n_538), .Y(n_1114) );
INVx1_ASAP7_75t_L g705 ( .A(n_540), .Y(n_705) );
AOI33xp33_ASAP7_75t_L g712 ( .A1(n_540), .A2(n_713), .A3(n_715), .B1(n_717), .B2(n_719), .B3(n_723), .Y(n_712) );
AOI33xp33_ASAP7_75t_L g796 ( .A1(n_540), .A2(n_696), .A3(n_797), .B1(n_799), .B2(n_801), .B3(n_802), .Y(n_796) );
NAND3xp33_ASAP7_75t_L g1263 ( .A(n_540), .B(n_1264), .C(n_1265), .Y(n_1263) );
NAND3xp33_ASAP7_75t_L g1295 ( .A(n_540), .B(n_1296), .C(n_1298), .Y(n_1295) );
NAND3xp33_ASAP7_75t_SL g926 ( .A(n_541), .B(n_927), .C(n_929), .Y(n_926) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
INVx1_ASAP7_75t_L g771 ( .A(n_545), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_545), .B(n_924), .Y(n_923) );
NAND2xp5_ASAP7_75t_L g1078 ( .A(n_545), .B(n_1079), .Y(n_1078) );
NAND2xp5_ASAP7_75t_L g1118 ( .A(n_545), .B(n_1119), .Y(n_1118) );
INVx1_ASAP7_75t_L g1173 ( .A(n_547), .Y(n_1173) );
AND2x2_ASAP7_75t_L g565 ( .A(n_548), .B(n_566), .Y(n_565) );
OAI31xp33_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_569), .A3(n_587), .B(n_590), .Y(n_549) );
BUFx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g1153 ( .A(n_556), .Y(n_1153) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g779 ( .A(n_559), .Y(n_779) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g897 ( .A(n_562), .Y(n_897) );
INVx2_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_565), .A2(n_567), .B1(n_904), .B2(n_905), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_565), .A2(n_567), .B1(n_1105), .B2(n_1106), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g1156 ( .A1(n_565), .A2(n_567), .B1(n_1157), .B2(n_1158), .Y(n_1156) );
AOI22xp5_ASAP7_75t_L g1191 ( .A1(n_565), .A2(n_567), .B1(n_1192), .B2(n_1193), .Y(n_1191) );
AND2x4_ASAP7_75t_L g1734 ( .A(n_566), .B(n_1017), .Y(n_1734) );
CKINVDCx11_ASAP7_75t_R g567 ( .A(n_568), .Y(n_567) );
OAI221xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_573), .B1(n_574), .B2(n_577), .C(n_578), .Y(n_570) );
OAI22xp33_ASAP7_75t_L g1369 ( .A1(n_571), .A2(n_1370), .B1(n_1372), .B2(n_1373), .Y(n_1369) );
OAI22xp33_ASAP7_75t_L g1383 ( .A1(n_571), .A2(n_1092), .B1(n_1384), .B2(n_1385), .Y(n_1383) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g1145 ( .A(n_572), .Y(n_1145) );
OAI221xp5_ASAP7_75t_L g892 ( .A1(n_574), .A2(n_893), .B1(n_895), .B2(n_896), .C(n_897), .Y(n_892) );
OAI221xp5_ASAP7_75t_L g1144 ( .A1(n_574), .A2(n_578), .B1(n_1123), .B2(n_1124), .C(n_1145), .Y(n_1144) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g921 ( .A(n_576), .Y(n_921) );
BUFx2_ASAP7_75t_L g1092 ( .A(n_576), .Y(n_1092) );
OAI221xp5_ASAP7_75t_L g916 ( .A1(n_578), .A2(n_917), .B1(n_919), .B2(n_920), .C(n_922), .Y(n_916) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g645 ( .A(n_585), .Y(n_645) );
AOI31xp33_ASAP7_75t_L g1388 ( .A1(n_590), .A2(n_1389), .A3(n_1398), .B(n_1405), .Y(n_1388) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
CKINVDCx8_ASAP7_75t_R g591 ( .A(n_592), .Y(n_591) );
OAI31xp33_ASAP7_75t_SL g1080 ( .A1(n_592), .A2(n_1081), .A3(n_1082), .B(n_1093), .Y(n_1080) );
AOI221x1_ASAP7_75t_SL g1169 ( .A1(n_592), .A2(n_634), .B1(n_1170), .B2(n_1199), .C(n_1209), .Y(n_1169) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
HB1xp67_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
OAI22x1_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B1(n_707), .B2(n_708), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g706 ( .A(n_601), .Y(n_706) );
AOI221x1_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_634), .B1(n_638), .B2(n_669), .C(n_671), .Y(n_601) );
NAND3xp33_ASAP7_75t_L g602 ( .A(n_603), .B(n_619), .C(n_628), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_604), .B(n_608), .Y(n_603) );
INVx5_ASAP7_75t_L g818 ( .A(n_604), .Y(n_818) );
AOI211xp5_ASAP7_75t_L g1273 ( .A1(n_604), .A2(n_1274), .B(n_1275), .C(n_1276), .Y(n_1273) );
CKINVDCx8_ASAP7_75t_R g1663 ( .A(n_604), .Y(n_1663) );
OAI21xp33_ASAP7_75t_L g1233 ( .A1(n_605), .A2(n_859), .B(n_1234), .Y(n_1233) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g1669 ( .A(n_606), .Y(n_1669) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g1232 ( .A(n_610), .Y(n_1232) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx1_ASAP7_75t_SL g622 ( .A(n_611), .Y(n_622) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g829 ( .A(n_613), .Y(n_829) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
HB1xp67_ASAP7_75t_L g1722 ( .A(n_616), .Y(n_1722) );
INVx3_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AOI222xp33_ASAP7_75t_L g822 ( .A1(n_618), .A2(n_823), .B1(n_824), .B2(n_826), .C1(n_827), .C2(n_830), .Y(n_822) );
AOI222xp33_ASAP7_75t_L g1205 ( .A1(n_618), .A2(n_827), .B1(n_1192), .B2(n_1193), .C1(n_1197), .C2(n_1206), .Y(n_1205) );
AOI222xp33_ASAP7_75t_L g1322 ( .A1(n_618), .A2(n_718), .B1(n_1323), .B2(n_1324), .C1(n_1325), .C2(n_1326), .Y(n_1322) );
AOI22xp33_ASAP7_75t_L g1660 ( .A1(n_618), .A2(n_828), .B1(n_1661), .B2(n_1662), .Y(n_1660) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_621), .B1(n_624), .B2(n_625), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_621), .A2(n_630), .B1(n_832), .B2(n_833), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g1200 ( .A1(n_621), .A2(n_630), .B1(n_1201), .B2(n_1202), .Y(n_1200) );
AOI22xp33_ASAP7_75t_L g1225 ( .A1(n_621), .A2(n_632), .B1(n_1226), .B2(n_1227), .Y(n_1225) );
AOI22xp33_ASAP7_75t_L g1278 ( .A1(n_621), .A2(n_625), .B1(n_1279), .B2(n_1280), .Y(n_1278) );
AOI22xp33_ASAP7_75t_L g1316 ( .A1(n_621), .A2(n_630), .B1(n_1317), .B2(n_1318), .Y(n_1316) );
AND2x4_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
AND2x6_ASAP7_75t_L g632 ( .A(n_622), .B(n_633), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_624), .A2(n_662), .B1(n_663), .B2(n_664), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_625), .A2(n_632), .B1(n_820), .B2(n_821), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g1203 ( .A1(n_625), .A2(n_632), .B1(n_1172), .B2(n_1204), .Y(n_1203) );
AOI221xp5_ASAP7_75t_L g1228 ( .A1(n_625), .A2(n_630), .B1(n_1229), .B2(n_1230), .C(n_1231), .Y(n_1228) );
AOI22xp33_ASAP7_75t_L g1319 ( .A1(n_625), .A2(n_632), .B1(n_1320), .B2(n_1321), .Y(n_1319) );
INVx4_ASAP7_75t_L g1670 ( .A(n_625), .Y(n_1670) );
AND2x4_ASAP7_75t_L g828 ( .A(n_626), .B(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_630), .B1(n_631), .B2(n_632), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g1281 ( .A1(n_630), .A2(n_632), .B1(n_1282), .B2(n_1283), .Y(n_1281) );
CKINVDCx6p67_ASAP7_75t_R g1665 ( .A(n_630), .Y(n_1665) );
INVx4_ASAP7_75t_L g1666 ( .A(n_632), .Y(n_1666) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_633), .Y(n_724) );
INVx2_ASAP7_75t_L g1137 ( .A(n_633), .Y(n_1137) );
BUFx6f_ASAP7_75t_L g1725 ( .A(n_633), .Y(n_1725) );
AOI221x1_ASAP7_75t_L g1223 ( .A1(n_634), .A2(n_669), .B1(n_1224), .B2(n_1235), .C(n_1249), .Y(n_1223) );
AOI211x1_ASAP7_75t_L g1314 ( .A1(n_634), .A2(n_1315), .B(n_1327), .C(n_1336), .Y(n_1314) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AOI211x1_ASAP7_75t_SL g816 ( .A1(n_635), .A2(n_817), .B(n_834), .C(n_867), .Y(n_816) );
AO211x2_ASAP7_75t_L g1271 ( .A1(n_635), .A2(n_1272), .B(n_1284), .C(n_1299), .Y(n_1271) );
AND2x4_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
AND2x4_ASAP7_75t_L g1671 ( .A(n_636), .B(n_637), .Y(n_1671) );
INVx2_ASAP7_75t_L g758 ( .A(n_637), .Y(n_758) );
BUFx2_ASAP7_75t_L g1731 ( .A(n_637), .Y(n_1731) );
NAND4xp25_ASAP7_75t_SL g638 ( .A(n_639), .B(n_646), .C(n_661), .D(n_666), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_641), .B1(n_643), .B2(n_644), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_641), .A2(n_874), .B1(n_875), .B2(n_876), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g1236 ( .A1(n_641), .A2(n_644), .B1(n_1237), .B2(n_1238), .Y(n_1236) );
AOI22xp33_ASAP7_75t_SL g1304 ( .A1(n_641), .A2(n_875), .B1(n_1305), .B2(n_1306), .Y(n_1304) );
AOI22xp33_ASAP7_75t_L g1331 ( .A1(n_641), .A2(n_644), .B1(n_1332), .B2(n_1333), .Y(n_1331) );
AOI22xp5_ASAP7_75t_L g1677 ( .A1(n_641), .A2(n_875), .B1(n_1678), .B2(n_1679), .Y(n_1677) );
AND2x4_ASAP7_75t_L g644 ( .A(n_642), .B(n_645), .Y(n_644) );
AND2x4_ASAP7_75t_L g875 ( .A(n_642), .B(n_645), .Y(n_875) );
AOI222xp33_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_648), .B1(n_651), .B2(n_652), .C1(n_655), .C2(n_656), .Y(n_646) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx2_ASAP7_75t_SL g840 ( .A(n_649), .Y(n_840) );
INVx2_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
BUFx6f_ASAP7_75t_L g1103 ( .A(n_650), .Y(n_1103) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g871 ( .A(n_654), .Y(n_871) );
AOI222xp33_ASAP7_75t_L g1239 ( .A1(n_654), .A2(n_656), .B1(n_1240), .B2(n_1241), .C1(n_1242), .C2(n_1243), .Y(n_1239) );
INVx2_ASAP7_75t_L g1675 ( .A(n_654), .Y(n_1675) );
AND2x4_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_657), .A2(n_727), .B1(n_728), .B2(n_755), .Y(n_754) );
AND2x4_ASAP7_75t_L g1736 ( .A(n_657), .B(n_1017), .Y(n_1736) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVxp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g668 ( .A(n_660), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_663), .A2(n_664), .B1(n_820), .B2(n_878), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g1246 ( .A1(n_663), .A2(n_1229), .B1(n_1247), .B2(n_1248), .Y(n_1246) );
AOI22xp33_ASAP7_75t_SL g1307 ( .A1(n_663), .A2(n_664), .B1(n_1280), .B2(n_1308), .Y(n_1307) );
AOI22xp33_ASAP7_75t_L g1334 ( .A1(n_663), .A2(n_1248), .B1(n_1320), .B2(n_1335), .Y(n_1334) );
INVx5_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx4_ASAP7_75t_L g1248 ( .A(n_665), .Y(n_1248) );
NAND4xp25_ASAP7_75t_SL g1235 ( .A(n_666), .B(n_1236), .C(n_1239), .D(n_1246), .Y(n_1235) );
CKINVDCx11_ASAP7_75t_R g666 ( .A(n_667), .Y(n_666) );
AOI211xp5_ASAP7_75t_L g868 ( .A1(n_667), .A2(n_779), .B(n_869), .C(n_870), .Y(n_868) );
AOI211xp5_ASAP7_75t_L g1300 ( .A1(n_667), .A2(n_840), .B(n_1301), .C(n_1302), .Y(n_1300) );
AOI211xp5_ASAP7_75t_L g1328 ( .A1(n_667), .A2(n_1254), .B(n_1329), .C(n_1330), .Y(n_1328) );
NOR3xp33_ASAP7_75t_L g1673 ( .A(n_667), .B(n_1674), .C(n_1676), .Y(n_1673) );
CKINVDCx16_ASAP7_75t_R g669 ( .A(n_670), .Y(n_669) );
AOI31xp33_ASAP7_75t_L g1299 ( .A1(n_670), .A2(n_1300), .A3(n_1304), .B(n_1307), .Y(n_1299) );
AOI31xp33_ASAP7_75t_L g1327 ( .A1(n_670), .A2(n_1328), .A3(n_1331), .B(n_1334), .Y(n_1327) );
AO21x1_ASAP7_75t_SL g1672 ( .A1(n_670), .A2(n_1673), .B(n_1677), .Y(n_1672) );
NAND4xp25_ASAP7_75t_L g671 ( .A(n_672), .B(n_683), .C(n_691), .D(n_699), .Y(n_671) );
NAND3xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_676), .C(n_681), .Y(n_672) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx2_ASAP7_75t_SL g1255 ( .A(n_675), .Y(n_1255) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
CKINVDCx8_ASAP7_75t_R g1045 ( .A(n_681), .Y(n_1045) );
NAND3xp33_ASAP7_75t_L g1256 ( .A(n_681), .B(n_1257), .C(n_1259), .Y(n_1256) );
NAND3xp33_ASAP7_75t_L g1288 ( .A(n_681), .B(n_1289), .C(n_1291), .Y(n_1288) );
INVx5_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx6_ASAP7_75t_L g851 ( .A(n_682), .Y(n_851) );
NAND3xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_689), .C(n_690), .Y(n_683) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AND2x4_ASAP7_75t_L g1003 ( .A(n_688), .B(n_1004), .Y(n_1003) );
INVx1_ASAP7_75t_L g1189 ( .A(n_688), .Y(n_1189) );
NAND3xp33_ASAP7_75t_L g1250 ( .A(n_690), .B(n_1251), .C(n_1253), .Y(n_1250) );
AOI33xp33_ASAP7_75t_L g1680 ( .A1(n_690), .A2(n_851), .A3(n_1681), .B1(n_1682), .B2(n_1683), .B3(n_1684), .Y(n_1680) );
AOI222xp33_ASAP7_75t_L g1748 ( .A1(n_690), .A2(n_851), .B1(n_1749), .B2(n_1750), .C1(n_1751), .C2(n_1756), .Y(n_1748) );
NAND3xp33_ASAP7_75t_L g691 ( .A(n_692), .B(n_695), .C(n_696), .Y(n_691) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
NAND3xp33_ASAP7_75t_L g1260 ( .A(n_696), .B(n_1261), .C(n_1262), .Y(n_1260) );
NAND3xp33_ASAP7_75t_L g1285 ( .A(n_696), .B(n_1286), .C(n_1287), .Y(n_1285) );
INVx3_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NAND3xp33_ASAP7_75t_L g699 ( .A(n_700), .B(n_702), .C(n_704), .Y(n_699) );
INVx1_ASAP7_75t_L g1723 ( .A(n_703), .Y(n_1723) );
AOI33xp33_ASAP7_75t_L g929 ( .A1(n_704), .A2(n_930), .A3(n_931), .B1(n_933), .B2(n_935), .B3(n_936), .Y(n_929) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx2_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
NAND4xp75_ASAP7_75t_L g710 ( .A(n_711), .B(n_732), .C(n_759), .D(n_761), .Y(n_710) );
AND2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_725), .Y(n_711) );
INVx1_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
BUFx2_ASAP7_75t_L g1050 ( .A(n_729), .Y(n_1050) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g950 ( .A(n_731), .Y(n_950) );
OAI21xp5_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_744), .B(n_757), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_737), .Y(n_733) );
INVx4_ASAP7_75t_L g844 ( .A(n_740), .Y(n_844) );
BUFx3_ASAP7_75t_L g849 ( .A(n_740), .Y(n_849) );
INVx2_ASAP7_75t_SL g901 ( .A(n_740), .Y(n_901) );
AND2x6_ASAP7_75t_L g1006 ( .A(n_742), .B(n_1004), .Y(n_1006) );
NAND2x1p5_ASAP7_75t_L g1021 ( .A(n_742), .B(n_1017), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_754), .Y(n_751) );
INVx2_ASAP7_75t_L g894 ( .A(n_752), .Y(n_894) );
BUFx3_ASAP7_75t_L g1044 ( .A(n_752), .Y(n_1044) );
BUFx3_ASAP7_75t_L g1183 ( .A(n_752), .Y(n_1183) );
OAI22xp5_ASAP7_75t_L g1752 ( .A1(n_752), .A2(n_1753), .B1(n_1754), .B2(n_1755), .Y(n_1752) );
BUFx6f_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
NAND2x1p5_ASAP7_75t_L g782 ( .A(n_755), .B(n_783), .Y(n_782) );
NAND2x1_ASAP7_75t_SL g1016 ( .A(n_755), .B(n_1017), .Y(n_1016) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
BUFx8_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g946 ( .A(n_758), .Y(n_946) );
OA22x2_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_883), .B1(n_884), .B2(n_1162), .Y(n_764) );
INVx1_ASAP7_75t_L g1162 ( .A(n_765), .Y(n_1162) );
INVx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
AOI21x1_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_814), .B(n_882), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
AND2x2_ASAP7_75t_L g882 ( .A(n_768), .B(n_815), .Y(n_882) );
XOR2x2_ASAP7_75t_L g768 ( .A(n_769), .B(n_813), .Y(n_768) );
NOR3xp33_ASAP7_75t_L g769 ( .A(n_770), .B(n_772), .C(n_795), .Y(n_769) );
AOI31xp33_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_784), .A3(n_787), .B(n_794), .Y(n_772) );
INVx1_ASAP7_75t_L g1099 ( .A(n_791), .Y(n_1099) );
NOR3xp33_ASAP7_75t_L g1179 ( .A(n_792), .B(n_1180), .C(n_1194), .Y(n_1179) );
INVx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
NAND4xp25_ASAP7_75t_L g795 ( .A(n_796), .B(n_804), .C(n_807), .D(n_810), .Y(n_795) );
BUFx6f_ASAP7_75t_L g862 ( .A(n_803), .Y(n_862) );
BUFx3_ASAP7_75t_L g977 ( .A(n_803), .Y(n_977) );
INVx1_ASAP7_75t_L g1063 ( .A(n_803), .Y(n_1063) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g881 ( .A(n_816), .Y(n_881) );
NAND4xp25_ASAP7_75t_L g817 ( .A(n_818), .B(n_819), .C(n_822), .D(n_831), .Y(n_817) );
BUFx2_ASAP7_75t_L g1208 ( .A(n_818), .Y(n_1208) );
NAND4xp25_ASAP7_75t_SL g1315 ( .A(n_818), .B(n_1316), .C(n_1319), .D(n_1322), .Y(n_1315) );
HB1xp67_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
HB1xp67_ASAP7_75t_L g1275 ( .A(n_825), .Y(n_1275) );
BUFx4f_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g1277 ( .A(n_828), .Y(n_1277) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_835), .B(n_852), .Y(n_834) );
AOI33xp33_ASAP7_75t_L g835 ( .A1(n_836), .A2(n_838), .A3(n_841), .B1(n_845), .B2(n_850), .B3(n_851), .Y(n_835) );
AOI33xp33_ASAP7_75t_L g1337 ( .A1(n_836), .A2(n_851), .A3(n_1338), .B1(n_1339), .B2(n_1340), .B3(n_1341), .Y(n_1337) );
BUFx3_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
NAND3xp33_ASAP7_75t_L g1292 ( .A(n_837), .B(n_1293), .C(n_1294), .Y(n_1292) );
INVx2_ASAP7_75t_SL g843 ( .A(n_844), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g1039 ( .A1(n_844), .A2(n_960), .B1(n_989), .B2(n_1033), .Y(n_1039) );
INVx2_ASAP7_75t_L g1195 ( .A(n_844), .Y(n_1195) );
INVx3_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx2_ASAP7_75t_SL g847 ( .A(n_848), .Y(n_847) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_848), .B(n_1004), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1365 ( .A(n_848), .B(n_1004), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1741 ( .A(n_848), .B(n_1004), .Y(n_1741) );
INVx1_ASAP7_75t_L g1381 ( .A(n_849), .Y(n_1381) );
AOI33xp33_ASAP7_75t_L g1344 ( .A1(n_853), .A2(n_1345), .A3(n_1348), .B1(n_1350), .B2(n_1351), .B3(n_1352), .Y(n_1344) );
BUFx3_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
HB1xp67_ASAP7_75t_L g1691 ( .A(n_856), .Y(n_1691) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g972 ( .A(n_859), .Y(n_972) );
AND2x4_ASAP7_75t_L g981 ( .A(n_859), .B(n_982), .Y(n_981) );
INVx1_ASAP7_75t_L g1401 ( .A(n_859), .Y(n_1401) );
BUFx6f_ASAP7_75t_L g1692 ( .A(n_859), .Y(n_1692) );
AOI31xp33_ASAP7_75t_L g867 ( .A1(n_868), .A2(n_873), .A3(n_877), .B(n_879), .Y(n_867) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
XNOR2xp5_ASAP7_75t_L g884 ( .A(n_885), .B(n_1046), .Y(n_884) );
AOI22x1_ASAP7_75t_L g885 ( .A1(n_886), .A2(n_887), .B1(n_941), .B2(n_942), .Y(n_885) );
INVx2_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
NAND3xp33_ASAP7_75t_L g888 ( .A(n_889), .B(n_923), .C(n_925), .Y(n_888) );
INVx2_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g1030 ( .A(n_894), .Y(n_1030) );
OAI22xp5_ASAP7_75t_L g898 ( .A1(n_899), .A2(n_900), .B1(n_901), .B2(n_902), .Y(n_898) );
OAI22xp5_ASAP7_75t_L g1032 ( .A1(n_901), .A2(n_1033), .B1(n_1037), .B2(n_1038), .Y(n_1032) );
OAI22xp5_ASAP7_75t_L g907 ( .A1(n_908), .A2(n_911), .B1(n_912), .B2(n_915), .Y(n_907) );
BUFx2_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
INVx2_ASAP7_75t_L g1085 ( .A(n_909), .Y(n_1085) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
BUFx3_ASAP7_75t_L g1036 ( .A(n_910), .Y(n_1036) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
INVx2_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx2_ASAP7_75t_L g1258 ( .A(n_914), .Y(n_1258) );
INVx2_ASAP7_75t_SL g1378 ( .A(n_914), .Y(n_1378) );
INVx1_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
NOR2xp33_ASAP7_75t_SL g925 ( .A(n_926), .B(n_938), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_939), .B(n_940), .Y(n_938) );
INVx2_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
XNOR2x1_ASAP7_75t_L g942 ( .A(n_943), .B(n_944), .Y(n_942) );
AND2x2_ASAP7_75t_L g944 ( .A(n_945), .B(n_998), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_946), .A2(n_947), .B1(n_992), .B2(n_993), .Y(n_945) );
NAND3xp33_ASAP7_75t_L g947 ( .A(n_948), .B(n_967), .C(n_984), .Y(n_947) );
AOI221xp5_ASAP7_75t_L g948 ( .A1(n_949), .A2(n_954), .B1(n_958), .B2(n_960), .C(n_961), .Y(n_948) );
BUFx2_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
HB1xp67_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
AOI21xp5_ASAP7_75t_L g1389 ( .A1(n_958), .A2(n_1380), .B(n_1390), .Y(n_1389) );
AOI221xp5_ASAP7_75t_L g1719 ( .A1(n_959), .A2(n_986), .B1(n_1720), .B2(n_1721), .C(n_1726), .Y(n_1719) );
INVx2_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
INVx2_ASAP7_75t_SL g965 ( .A(n_966), .Y(n_965) );
AOI221xp5_ASAP7_75t_L g967 ( .A1(n_968), .A2(n_976), .B1(n_978), .B2(n_980), .C(n_981), .Y(n_967) );
BUFx2_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
INVx1_ASAP7_75t_L g1075 ( .A(n_970), .Y(n_1075) );
BUFx3_ASAP7_75t_L g1346 ( .A(n_970), .Y(n_1346) );
INVx1_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
INVx1_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
INVx1_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
AOI221xp5_ASAP7_75t_L g1398 ( .A1(n_978), .A2(n_981), .B1(n_1385), .B2(n_1399), .C(n_1404), .Y(n_1398) );
BUFx6f_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
OAI22xp33_ASAP7_75t_L g1040 ( .A1(n_980), .A2(n_985), .B1(n_1041), .B2(n_1044), .Y(n_1040) );
INVx1_ASAP7_75t_SL g982 ( .A(n_983), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_985), .A2(n_986), .B1(n_989), .B2(n_990), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g1405 ( .A1(n_986), .A2(n_990), .B1(n_1382), .B2(n_1384), .Y(n_1405) );
INVx6_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
INVx1_ASAP7_75t_L g1055 ( .A(n_988), .Y(n_1055) );
INVx2_ASAP7_75t_L g1067 ( .A(n_988), .Y(n_1067) );
OR2x2_ASAP7_75t_L g1668 ( .A(n_988), .B(n_1669), .Y(n_1668) );
INVx4_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
AOI21xp33_ASAP7_75t_L g1386 ( .A1(n_993), .A2(n_1387), .B(n_1388), .Y(n_1386) );
INVx5_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
AND2x4_ASAP7_75t_L g994 ( .A(n_995), .B(n_997), .Y(n_994) );
INVx2_ASAP7_75t_L g1747 ( .A(n_995), .Y(n_1747) );
INVx3_ASAP7_75t_L g1017 ( .A(n_996), .Y(n_1017) );
NOR3xp33_ASAP7_75t_SL g998 ( .A(n_999), .B(n_1013), .C(n_1022), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1007), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_1001), .A2(n_1002), .B1(n_1005), .B2(n_1006), .Y(n_1000) );
BUFx2_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
BUFx2_ASAP7_75t_L g1360 ( .A(n_1003), .Y(n_1360) );
BUFx2_ASAP7_75t_L g1745 ( .A(n_1003), .Y(n_1745) );
AND2x4_ASAP7_75t_L g1009 ( .A(n_1004), .B(n_1010), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g1358 ( .A1(n_1006), .A2(n_1359), .B1(n_1360), .B2(n_1361), .Y(n_1358) );
AOI22xp5_ASAP7_75t_L g1739 ( .A1(n_1006), .A2(n_1740), .B1(n_1741), .B2(n_1742), .Y(n_1739) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_1008), .A2(n_1009), .B1(n_1011), .B2(n_1012), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1362 ( .A1(n_1009), .A2(n_1363), .B1(n_1364), .B2(n_1365), .Y(n_1362) );
INVx2_ASAP7_75t_SL g1014 ( .A(n_1015), .Y(n_1014) );
INVx2_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
AND2x4_ASAP7_75t_L g1738 ( .A(n_1017), .B(n_1245), .Y(n_1738) );
BUFx4f_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
BUFx2_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
BUFx2_ASAP7_75t_L g1367 ( .A(n_1021), .Y(n_1367) );
OAI33xp33_ASAP7_75t_L g1022 ( .A1(n_1023), .A2(n_1026), .A3(n_1032), .B1(n_1039), .B2(n_1040), .B3(n_1045), .Y(n_1022) );
OAI33xp33_ASAP7_75t_L g1368 ( .A1(n_1023), .A2(n_1045), .A3(n_1369), .B1(n_1374), .B2(n_1379), .B3(n_1383), .Y(n_1368) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
OAI22xp33_ASAP7_75t_L g1026 ( .A1(n_1027), .A2(n_1029), .B1(n_1030), .B2(n_1031), .Y(n_1026) );
INVx2_ASAP7_75t_L g1027 ( .A(n_1028), .Y(n_1027) );
INVx2_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
INVx2_ASAP7_75t_L g1034 ( .A(n_1035), .Y(n_1034) );
INVx2_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
BUFx2_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
INVx2_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
XOR2x2_ASAP7_75t_L g1046 ( .A(n_1047), .B(n_1115), .Y(n_1046) );
AND4x1_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1078), .C(n_1080), .D(n_1107), .Y(n_1048) );
NOR3xp33_ASAP7_75t_SL g1049 ( .A(n_1050), .B(n_1051), .C(n_1076), .Y(n_1049) );
NOR3xp33_ASAP7_75t_SL g1120 ( .A(n_1050), .B(n_1121), .C(n_1138), .Y(n_1120) );
OAI221xp5_ASAP7_75t_L g1052 ( .A1(n_1053), .A2(n_1056), .B1(n_1057), .B2(n_1058), .C(n_1061), .Y(n_1052) );
OAI221xp5_ASAP7_75t_L g1122 ( .A1(n_1053), .A2(n_1058), .B1(n_1123), .B2(n_1124), .C(n_1125), .Y(n_1122) );
OAI221xp5_ASAP7_75t_L g1210 ( .A1(n_1053), .A2(n_1190), .B1(n_1211), .B2(n_1212), .C(n_1213), .Y(n_1210) );
BUFx2_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
OAI221xp5_ASAP7_75t_L g1216 ( .A1(n_1054), .A2(n_1069), .B1(n_1174), .B2(n_1175), .C(n_1217), .Y(n_1216) );
INVx2_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
BUFx2_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1060), .Y(n_1131) );
INVx2_ASAP7_75t_SL g1394 ( .A(n_1060), .Y(n_1394) );
INVx1_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
OAI221xp5_ASAP7_75t_L g1065 ( .A1(n_1066), .A2(n_1068), .B1(n_1069), .B2(n_1072), .C(n_1073), .Y(n_1065) );
OAI221xp5_ASAP7_75t_L g1129 ( .A1(n_1066), .A2(n_1130), .B1(n_1131), .B2(n_1132), .C(n_1133), .Y(n_1129) );
INVx2_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1067), .Y(n_1112) );
INVx2_ASAP7_75t_L g1069 ( .A(n_1070), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1075), .Y(n_1074) );
OAI22xp5_ASAP7_75t_L g1083 ( .A1(n_1084), .A2(n_1086), .B1(n_1087), .B2(n_1090), .Y(n_1083) );
OAI22xp5_ASAP7_75t_L g1374 ( .A1(n_1084), .A2(n_1375), .B1(n_1376), .B2(n_1377), .Y(n_1374) );
OAI22xp5_ASAP7_75t_L g1379 ( .A1(n_1084), .A2(n_1380), .B1(n_1381), .B2(n_1382), .Y(n_1379) );
INVx2_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
INVx2_ASAP7_75t_L g1095 ( .A(n_1085), .Y(n_1095) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1088), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
OAI221xp5_ASAP7_75t_L g1094 ( .A1(n_1095), .A2(n_1096), .B1(n_1097), .B2(n_1100), .C(n_1101), .Y(n_1094) );
OAI221xp5_ASAP7_75t_L g1150 ( .A1(n_1095), .A2(n_1151), .B1(n_1152), .B2(n_1154), .C(n_1155), .Y(n_1150) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
NOR2xp33_ASAP7_75t_L g1107 ( .A(n_1108), .B(n_1110), .Y(n_1107) );
XNOR2xp5_ASAP7_75t_L g1115 ( .A(n_1116), .B(n_1117), .Y(n_1115) );
AND4x1_ASAP7_75t_L g1117 ( .A(n_1118), .B(n_1120), .C(n_1141), .D(n_1159), .Y(n_1117) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1126), .Y(n_1212) );
CKINVDCx5p33_ASAP7_75t_R g1127 ( .A(n_1128), .Y(n_1127) );
BUFx3_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1137), .Y(n_1136) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1137), .Y(n_1347) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
NOR2xp33_ASAP7_75t_L g1159 ( .A(n_1160), .B(n_1161), .Y(n_1159) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
XNOR2xp5_ASAP7_75t_L g1164 ( .A(n_1165), .B(n_1311), .Y(n_1164) );
AOI22xp5_ASAP7_75t_L g1165 ( .A1(n_1166), .A2(n_1269), .B1(n_1309), .B2(n_1310), .Y(n_1165) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1166), .Y(n_1309) );
AOI22xp5_ASAP7_75t_L g1166 ( .A1(n_1167), .A2(n_1168), .B1(n_1221), .B2(n_1268), .Y(n_1166) );
INVx2_ASAP7_75t_SL g1167 ( .A(n_1168), .Y(n_1167) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1169), .Y(n_1220) );
NAND3xp33_ASAP7_75t_L g1170 ( .A(n_1171), .B(n_1176), .C(n_1179), .Y(n_1170) );
OAI21xp5_ASAP7_75t_SL g1180 ( .A1(n_1181), .A2(n_1185), .B(n_1191), .Y(n_1180) );
OAI21xp5_ASAP7_75t_L g1181 ( .A1(n_1182), .A2(n_1183), .B(n_1184), .Y(n_1181) );
OAI22xp5_ASAP7_75t_L g1185 ( .A1(n_1186), .A2(n_1188), .B1(n_1189), .B2(n_1190), .Y(n_1185) );
BUFx2_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
NAND4xp25_ASAP7_75t_SL g1199 ( .A(n_1200), .B(n_1203), .C(n_1205), .D(n_1208), .Y(n_1199) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1207), .Y(n_1206) );
HB1xp67_ASAP7_75t_L g1221 ( .A(n_1222), .Y(n_1221) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1222), .Y(n_1268) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1223), .Y(n_1267) );
NAND2xp5_ASAP7_75t_L g1224 ( .A(n_1225), .B(n_1228), .Y(n_1224) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1244), .Y(n_1243) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1245), .Y(n_1244) );
NAND4xp25_ASAP7_75t_L g1249 ( .A(n_1250), .B(n_1256), .C(n_1260), .D(n_1263), .Y(n_1249) );
INVx2_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1269), .Y(n_1310) );
HB1xp67_ASAP7_75t_L g1269 ( .A(n_1270), .Y(n_1269) );
NAND3xp33_ASAP7_75t_L g1272 ( .A(n_1273), .B(n_1278), .C(n_1281), .Y(n_1272) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1277), .Y(n_1325) );
NAND4xp25_ASAP7_75t_L g1284 ( .A(n_1285), .B(n_1288), .C(n_1292), .D(n_1295), .Y(n_1284) );
HB1xp67_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
XNOR2xp5_ASAP7_75t_L g1312 ( .A(n_1313), .B(n_1353), .Y(n_1312) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_1337), .B(n_1344), .Y(n_1336) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1343), .Y(n_1342) );
NAND2xp5_ASAP7_75t_L g1658 ( .A(n_1349), .B(n_1659), .Y(n_1658) );
XNOR2x1_ASAP7_75t_L g1353 ( .A(n_1354), .B(n_1355), .Y(n_1353) );
AND2x2_ASAP7_75t_L g1355 ( .A(n_1356), .B(n_1386), .Y(n_1355) );
NOR3xp33_ASAP7_75t_SL g1356 ( .A(n_1357), .B(n_1366), .C(n_1368), .Y(n_1356) );
NAND2xp5_ASAP7_75t_L g1357 ( .A(n_1358), .B(n_1362), .Y(n_1357) );
OAI211xp5_ASAP7_75t_L g1393 ( .A1(n_1361), .A2(n_1394), .B(n_1395), .C(n_1396), .Y(n_1393) );
INVx3_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
INVx1_ASAP7_75t_SL g1391 ( .A(n_1392), .Y(n_1391) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1401), .Y(n_1400) );
INVx1_ASAP7_75t_L g1402 ( .A(n_1403), .Y(n_1402) );
OAI221xp5_ASAP7_75t_L g1406 ( .A1(n_1407), .A2(n_1648), .B1(n_1652), .B2(n_1695), .C(n_1700), .Y(n_1406) );
AOI21xp5_ASAP7_75t_L g1407 ( .A1(n_1408), .A2(n_1553), .B(n_1597), .Y(n_1407) );
NAND5xp2_ASAP7_75t_SL g1408 ( .A(n_1409), .B(n_1492), .C(n_1521), .D(n_1544), .E(n_1548), .Y(n_1408) );
AOI21xp5_ASAP7_75t_L g1409 ( .A1(n_1410), .A2(n_1448), .B(n_1470), .Y(n_1409) );
AND2x2_ASAP7_75t_L g1410 ( .A(n_1411), .B(n_1431), .Y(n_1410) );
AND2x2_ASAP7_75t_L g1509 ( .A(n_1411), .B(n_1458), .Y(n_1509) );
AND2x2_ASAP7_75t_L g1546 ( .A(n_1411), .B(n_1547), .Y(n_1546) );
NAND2xp5_ASAP7_75t_L g1571 ( .A(n_1411), .B(n_1481), .Y(n_1571) );
NOR2xp33_ASAP7_75t_L g1582 ( .A(n_1411), .B(n_1458), .Y(n_1582) );
INVx2_ASAP7_75t_L g1411 ( .A(n_1412), .Y(n_1411) );
AND2x2_ASAP7_75t_L g1478 ( .A(n_1412), .B(n_1479), .Y(n_1478) );
NAND2xp5_ASAP7_75t_L g1491 ( .A(n_1412), .B(n_1458), .Y(n_1491) );
BUFx2_ASAP7_75t_L g1498 ( .A(n_1412), .Y(n_1498) );
INVx2_ASAP7_75t_L g1505 ( .A(n_1412), .Y(n_1505) );
NAND2xp5_ASAP7_75t_L g1556 ( .A(n_1412), .B(n_1431), .Y(n_1556) );
OR2x2_ASAP7_75t_L g1580 ( .A(n_1412), .B(n_1489), .Y(n_1580) );
NAND2xp5_ASAP7_75t_L g1613 ( .A(n_1412), .B(n_1481), .Y(n_1613) );
AND2x2_ASAP7_75t_L g1412 ( .A(n_1413), .B(n_1425), .Y(n_1412) );
AND2x4_ASAP7_75t_L g1414 ( .A(n_1415), .B(n_1420), .Y(n_1414) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1416), .Y(n_1415) );
OR2x2_ASAP7_75t_L g1445 ( .A(n_1416), .B(n_1421), .Y(n_1445) );
NAND2xp5_ASAP7_75t_L g1416 ( .A(n_1417), .B(n_1419), .Y(n_1416) );
HB1xp67_ASAP7_75t_L g1766 ( .A(n_1417), .Y(n_1766) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
INVx1_ASAP7_75t_L g1428 ( .A(n_1419), .Y(n_1428) );
AND2x4_ASAP7_75t_L g1422 ( .A(n_1420), .B(n_1423), .Y(n_1422) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1421), .Y(n_1420) );
OR2x2_ASAP7_75t_L g1447 ( .A(n_1421), .B(n_1424), .Y(n_1447) );
BUFx2_ASAP7_75t_L g1453 ( .A(n_1422), .Y(n_1453) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1424), .Y(n_1423) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1426), .Y(n_1467) );
BUFx3_ASAP7_75t_L g1513 ( .A(n_1426), .Y(n_1513) );
AND2x4_ASAP7_75t_L g1426 ( .A(n_1427), .B(n_1429), .Y(n_1426) );
AND2x2_ASAP7_75t_L g1436 ( .A(n_1427), .B(n_1429), .Y(n_1436) );
HB1xp67_ASAP7_75t_L g1764 ( .A(n_1427), .Y(n_1764) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
AND2x4_ASAP7_75t_L g1430 ( .A(n_1428), .B(n_1429), .Y(n_1430) );
INVx2_ASAP7_75t_L g1456 ( .A(n_1430), .Y(n_1456) );
AND2x2_ASAP7_75t_L g1431 ( .A(n_1432), .B(n_1437), .Y(n_1431) );
NAND2xp5_ASAP7_75t_L g1484 ( .A(n_1432), .B(n_1485), .Y(n_1484) );
AND2x2_ASAP7_75t_L g1541 ( .A(n_1432), .B(n_1476), .Y(n_1541) );
A2O1A1Ixp33_ASAP7_75t_L g1614 ( .A1(n_1432), .A2(n_1615), .B(n_1618), .C(n_1619), .Y(n_1614) );
INVxp67_ASAP7_75t_L g1432 ( .A(n_1433), .Y(n_1432) );
BUFx2_ASAP7_75t_L g1479 ( .A(n_1433), .Y(n_1479) );
BUFx3_ASAP7_75t_L g1489 ( .A(n_1433), .Y(n_1489) );
AND2x2_ASAP7_75t_L g1552 ( .A(n_1433), .B(n_1476), .Y(n_1552) );
AND2x2_ASAP7_75t_L g1433 ( .A(n_1434), .B(n_1435), .Y(n_1433) );
AND2x2_ASAP7_75t_L g1510 ( .A(n_1437), .B(n_1479), .Y(n_1510) );
INVx1_ASAP7_75t_L g1617 ( .A(n_1437), .Y(n_1617) );
AND2x2_ASAP7_75t_L g1437 ( .A(n_1438), .B(n_1442), .Y(n_1437) );
NAND2xp5_ASAP7_75t_L g1494 ( .A(n_1438), .B(n_1489), .Y(n_1494) );
NOR2xp33_ASAP7_75t_L g1560 ( .A(n_1438), .B(n_1479), .Y(n_1560) );
INVx2_ASAP7_75t_L g1438 ( .A(n_1439), .Y(n_1438) );
OR2x2_ASAP7_75t_L g1477 ( .A(n_1439), .B(n_1442), .Y(n_1477) );
AND2x2_ASAP7_75t_L g1485 ( .A(n_1439), .B(n_1486), .Y(n_1485) );
AND2x2_ASAP7_75t_L g1488 ( .A(n_1439), .B(n_1489), .Y(n_1488) );
AND2x2_ASAP7_75t_L g1525 ( .A(n_1439), .B(n_1442), .Y(n_1525) );
NOR2xp33_ASAP7_75t_L g1532 ( .A(n_1439), .B(n_1489), .Y(n_1532) );
AND2x2_ASAP7_75t_L g1439 ( .A(n_1440), .B(n_1441), .Y(n_1439) );
INVx2_ASAP7_75t_SL g1486 ( .A(n_1442), .Y(n_1486) );
AND2x2_ASAP7_75t_L g1506 ( .A(n_1442), .B(n_1489), .Y(n_1506) );
OAI22xp5_ASAP7_75t_L g1443 ( .A1(n_1444), .A2(n_1445), .B1(n_1446), .B2(n_1447), .Y(n_1443) );
BUFx6f_ASAP7_75t_L g1461 ( .A(n_1445), .Y(n_1461) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1447), .Y(n_1464) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1448), .Y(n_1566) );
AND2x2_ASAP7_75t_L g1448 ( .A(n_1449), .B(n_1457), .Y(n_1448) );
NAND2xp5_ASAP7_75t_L g1519 ( .A(n_1449), .B(n_1520), .Y(n_1519) );
INVx2_ASAP7_75t_L g1536 ( .A(n_1449), .Y(n_1536) );
AND2x2_ASAP7_75t_L g1550 ( .A(n_1449), .B(n_1551), .Y(n_1550) );
NAND2xp5_ASAP7_75t_L g1586 ( .A(n_1449), .B(n_1458), .Y(n_1586) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1450), .Y(n_1449) );
INVx1_ASAP7_75t_L g1600 ( .A(n_1450), .Y(n_1600) );
AND2x2_ASAP7_75t_L g1634 ( .A(n_1450), .B(n_1471), .Y(n_1634) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1451), .Y(n_1450) );
OR2x2_ASAP7_75t_L g1527 ( .A(n_1451), .B(n_1471), .Y(n_1527) );
AND2x2_ASAP7_75t_L g1529 ( .A(n_1451), .B(n_1482), .Y(n_1529) );
INVx1_ASAP7_75t_L g1609 ( .A(n_1451), .Y(n_1609) );
AND2x2_ASAP7_75t_L g1451 ( .A(n_1452), .B(n_1454), .Y(n_1451) );
INVx2_ASAP7_75t_L g1455 ( .A(n_1456), .Y(n_1455) );
OAI22xp5_ASAP7_75t_L g1466 ( .A1(n_1456), .A2(n_1467), .B1(n_1468), .B2(n_1469), .Y(n_1466) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1456), .Y(n_1651) );
NAND2xp5_ASAP7_75t_L g1528 ( .A(n_1457), .B(n_1529), .Y(n_1528) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1457), .Y(n_1596) );
INVx1_ASAP7_75t_L g1457 ( .A(n_1458), .Y(n_1457) );
AND2x2_ASAP7_75t_L g1499 ( .A(n_1458), .B(n_1471), .Y(n_1499) );
INVx2_ASAP7_75t_SL g1535 ( .A(n_1458), .Y(n_1535) );
AND2x4_ASAP7_75t_L g1551 ( .A(n_1458), .B(n_1482), .Y(n_1551) );
HB1xp67_ASAP7_75t_L g1588 ( .A(n_1458), .Y(n_1588) );
CKINVDCx5p33_ASAP7_75t_R g1458 ( .A(n_1459), .Y(n_1458) );
AND2x2_ASAP7_75t_L g1481 ( .A(n_1459), .B(n_1482), .Y(n_1481) );
AND2x2_ASAP7_75t_L g1543 ( .A(n_1459), .B(n_1471), .Y(n_1543) );
OR2x2_ASAP7_75t_L g1459 ( .A(n_1460), .B(n_1466), .Y(n_1459) );
OAI22xp5_ASAP7_75t_L g1460 ( .A1(n_1461), .A2(n_1462), .B1(n_1463), .B2(n_1465), .Y(n_1460) );
BUFx3_ASAP7_75t_L g1516 ( .A(n_1461), .Y(n_1516) );
HB1xp67_ASAP7_75t_L g1518 ( .A(n_1463), .Y(n_1518) );
INVx1_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
OAI211xp5_ASAP7_75t_SL g1470 ( .A1(n_1471), .A2(n_1474), .B(n_1480), .C(n_1487), .Y(n_1470) );
INVx3_ASAP7_75t_L g1482 ( .A(n_1471), .Y(n_1482) );
INVx1_ASAP7_75t_L g1573 ( .A(n_1471), .Y(n_1573) );
AND2x2_ASAP7_75t_L g1471 ( .A(n_1472), .B(n_1473), .Y(n_1471) );
OAI321xp33_ASAP7_75t_L g1579 ( .A1(n_1474), .A2(n_1494), .A3(n_1525), .B1(n_1573), .B2(n_1580), .C(n_1581), .Y(n_1579) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
AND2x2_ASAP7_75t_L g1601 ( .A(n_1475), .B(n_1535), .Y(n_1601) );
NAND2xp5_ASAP7_75t_L g1625 ( .A(n_1475), .B(n_1626), .Y(n_1625) );
AND2x2_ASAP7_75t_L g1475 ( .A(n_1476), .B(n_1478), .Y(n_1475) );
AND2x2_ASAP7_75t_L g1590 ( .A(n_1476), .B(n_1505), .Y(n_1590) );
INVx1_ASAP7_75t_L g1476 ( .A(n_1477), .Y(n_1476) );
OR2x2_ASAP7_75t_L g1603 ( .A(n_1477), .B(n_1580), .Y(n_1603) );
NAND2xp5_ASAP7_75t_L g1611 ( .A(n_1478), .B(n_1525), .Y(n_1611) );
NOR2x1_ASAP7_75t_L g1578 ( .A(n_1479), .B(n_1486), .Y(n_1578) );
AND2x2_ASAP7_75t_L g1584 ( .A(n_1479), .B(n_1525), .Y(n_1584) );
NAND2xp5_ASAP7_75t_L g1480 ( .A(n_1481), .B(n_1483), .Y(n_1480) );
AOI221xp5_ASAP7_75t_L g1554 ( .A1(n_1481), .A2(n_1555), .B1(n_1557), .B2(n_1563), .C(n_1564), .Y(n_1554) );
NOR2xp33_ASAP7_75t_L g1490 ( .A(n_1482), .B(n_1491), .Y(n_1490) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1482), .Y(n_1502) );
OR2x2_ASAP7_75t_L g1608 ( .A(n_1482), .B(n_1609), .Y(n_1608) );
AOI221xp5_ASAP7_75t_L g1623 ( .A1(n_1482), .A2(n_1526), .B1(n_1624), .B2(n_1627), .C(n_1630), .Y(n_1623) );
O2A1O1Ixp33_ASAP7_75t_L g1567 ( .A1(n_1483), .A2(n_1550), .B(n_1568), .C(n_1570), .Y(n_1567) );
AOI222xp33_ASAP7_75t_L g1604 ( .A1(n_1483), .A2(n_1529), .B1(n_1605), .B2(n_1607), .C1(n_1610), .C2(n_1612), .Y(n_1604) );
INVx2_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
OR2x2_ASAP7_75t_L g1606 ( .A(n_1484), .B(n_1497), .Y(n_1606) );
AND2x2_ASAP7_75t_L g1547 ( .A(n_1485), .B(n_1489), .Y(n_1547) );
NAND2xp5_ASAP7_75t_L g1565 ( .A(n_1485), .B(n_1498), .Y(n_1565) );
INVx1_ASAP7_75t_L g1616 ( .A(n_1485), .Y(n_1616) );
AND2x2_ASAP7_75t_L g1629 ( .A(n_1486), .B(n_1489), .Y(n_1629) );
NAND2xp5_ASAP7_75t_L g1487 ( .A(n_1488), .B(n_1490), .Y(n_1487) );
INVx1_ASAP7_75t_L g1631 ( .A(n_1488), .Y(n_1631) );
AND2x2_ASAP7_75t_L g1645 ( .A(n_1488), .B(n_1505), .Y(n_1645) );
OR2x2_ASAP7_75t_L g1523 ( .A(n_1489), .B(n_1524), .Y(n_1523) );
AND2x2_ASAP7_75t_L g1595 ( .A(n_1489), .B(n_1538), .Y(n_1595) );
AND2x2_ASAP7_75t_L g1618 ( .A(n_1489), .B(n_1590), .Y(n_1618) );
O2A1O1Ixp33_ASAP7_75t_L g1630 ( .A1(n_1491), .A2(n_1631), .B(n_1632), .C(n_1633), .Y(n_1630) );
A2O1A1Ixp33_ASAP7_75t_L g1492 ( .A1(n_1493), .A2(n_1495), .B(n_1500), .C(n_1519), .Y(n_1492) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1494), .Y(n_1493) );
NAND2xp5_ASAP7_75t_L g1522 ( .A(n_1494), .B(n_1523), .Y(n_1522) );
O2A1O1Ixp33_ASAP7_75t_L g1564 ( .A1(n_1494), .A2(n_1498), .B(n_1565), .C(n_1566), .Y(n_1564) );
NOR2xp33_ASAP7_75t_L g1570 ( .A(n_1494), .B(n_1571), .Y(n_1570) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1496), .Y(n_1495) );
NAND2xp5_ASAP7_75t_L g1496 ( .A(n_1497), .B(n_1499), .Y(n_1496) );
NAND2xp5_ASAP7_75t_L g1569 ( .A(n_1497), .B(n_1532), .Y(n_1569) );
NAND2xp5_ASAP7_75t_L g1577 ( .A(n_1497), .B(n_1578), .Y(n_1577) );
INVx2_ASAP7_75t_L g1497 ( .A(n_1498), .Y(n_1497) );
AOI321xp33_ASAP7_75t_L g1521 ( .A1(n_1498), .A2(n_1522), .A3(n_1526), .B1(n_1528), .B2(n_1530), .C(n_1539), .Y(n_1521) );
NAND2xp5_ASAP7_75t_L g1542 ( .A(n_1498), .B(n_1543), .Y(n_1542) );
AND2x2_ASAP7_75t_L g1559 ( .A(n_1498), .B(n_1560), .Y(n_1559) );
NAND2xp5_ASAP7_75t_SL g1594 ( .A(n_1498), .B(n_1532), .Y(n_1594) );
INVx1_ASAP7_75t_L g1562 ( .A(n_1499), .Y(n_1562) );
OAI211xp5_ASAP7_75t_SL g1500 ( .A1(n_1501), .A2(n_1503), .B(n_1507), .C(n_1511), .Y(n_1500) );
OAI22xp5_ASAP7_75t_L g1557 ( .A1(n_1501), .A2(n_1558), .B1(n_1561), .B2(n_1562), .Y(n_1557) );
INVx1_ASAP7_75t_L g1501 ( .A(n_1502), .Y(n_1501) );
A2O1A1Ixp33_ASAP7_75t_L g1592 ( .A1(n_1502), .A2(n_1593), .B(n_1595), .C(n_1596), .Y(n_1592) );
AOI31xp33_ASAP7_75t_L g1643 ( .A1(n_1503), .A2(n_1540), .A3(n_1644), .B(n_1646), .Y(n_1643) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1504), .Y(n_1503) );
AND2x2_ASAP7_75t_L g1504 ( .A(n_1505), .B(n_1506), .Y(n_1504) );
AND2x2_ASAP7_75t_L g1538 ( .A(n_1505), .B(n_1525), .Y(n_1538) );
AND2x2_ASAP7_75t_L g1640 ( .A(n_1505), .B(n_1535), .Y(n_1640) );
INVxp67_ASAP7_75t_L g1561 ( .A(n_1506), .Y(n_1561) );
INVxp67_ASAP7_75t_L g1507 ( .A(n_1508), .Y(n_1507) );
AND2x2_ASAP7_75t_L g1508 ( .A(n_1509), .B(n_1510), .Y(n_1508) );
INVx2_ASAP7_75t_L g1591 ( .A(n_1511), .Y(n_1591) );
INVx3_ASAP7_75t_L g1511 ( .A(n_1512), .Y(n_1511) );
INVx3_ASAP7_75t_L g1520 ( .A(n_1512), .Y(n_1520) );
OAI22xp33_ASAP7_75t_L g1514 ( .A1(n_1515), .A2(n_1516), .B1(n_1517), .B2(n_1518), .Y(n_1514) );
AOI21xp5_ASAP7_75t_L g1539 ( .A1(n_1524), .A2(n_1540), .B(n_1542), .Y(n_1539) );
INVx1_ASAP7_75t_L g1524 ( .A(n_1525), .Y(n_1524) );
AND2x2_ASAP7_75t_L g1545 ( .A(n_1526), .B(n_1546), .Y(n_1545) );
INVx1_ASAP7_75t_L g1526 ( .A(n_1527), .Y(n_1526) );
NOR2xp33_ASAP7_75t_L g1534 ( .A(n_1527), .B(n_1535), .Y(n_1534) );
OAI22xp33_ASAP7_75t_L g1530 ( .A1(n_1531), .A2(n_1533), .B1(n_1536), .B2(n_1537), .Y(n_1530) );
INVxp33_ASAP7_75t_L g1531 ( .A(n_1532), .Y(n_1531) );
INVx1_ASAP7_75t_L g1533 ( .A(n_1534), .Y(n_1533) );
NAND2xp5_ASAP7_75t_L g1575 ( .A(n_1535), .B(n_1576), .Y(n_1575) );
NOR2xp33_ASAP7_75t_L g1602 ( .A(n_1535), .B(n_1603), .Y(n_1602) );
INVx2_ASAP7_75t_L g1626 ( .A(n_1535), .Y(n_1626) );
NAND2xp5_ASAP7_75t_L g1628 ( .A(n_1535), .B(n_1629), .Y(n_1628) );
NOR2xp33_ASAP7_75t_L g1647 ( .A(n_1535), .B(n_1608), .Y(n_1647) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1536), .Y(n_1563) );
A2O1A1Ixp33_ASAP7_75t_L g1572 ( .A1(n_1536), .A2(n_1573), .B(n_1574), .C(n_1579), .Y(n_1572) );
INVx1_ASAP7_75t_L g1537 ( .A(n_1538), .Y(n_1537) );
INVx1_ASAP7_75t_L g1540 ( .A(n_1541), .Y(n_1540) );
NOR2xp33_ASAP7_75t_L g1642 ( .A(n_1541), .B(n_1547), .Y(n_1642) );
AOI221xp5_ASAP7_75t_L g1583 ( .A1(n_1543), .A2(n_1552), .B1(n_1584), .B2(n_1585), .C(n_1587), .Y(n_1583) );
CKINVDCx5p33_ASAP7_75t_R g1622 ( .A(n_1543), .Y(n_1622) );
INVxp67_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
INVxp67_ASAP7_75t_L g1548 ( .A(n_1549), .Y(n_1548) );
AND2x2_ASAP7_75t_L g1549 ( .A(n_1550), .B(n_1552), .Y(n_1549) );
NAND5xp2_ASAP7_75t_L g1553 ( .A(n_1554), .B(n_1567), .C(n_1572), .D(n_1583), .E(n_1592), .Y(n_1553) );
INVx1_ASAP7_75t_L g1555 ( .A(n_1556), .Y(n_1555) );
INVx1_ASAP7_75t_L g1558 ( .A(n_1559), .Y(n_1558) );
AOI22xp5_ASAP7_75t_L g1598 ( .A1(n_1563), .A2(n_1599), .B1(n_1601), .B2(n_1602), .Y(n_1598) );
INVx1_ASAP7_75t_L g1568 ( .A(n_1569), .Y(n_1568) );
INVx1_ASAP7_75t_L g1636 ( .A(n_1571), .Y(n_1636) );
INVxp67_ASAP7_75t_L g1574 ( .A(n_1575), .Y(n_1574) );
INVx1_ASAP7_75t_L g1576 ( .A(n_1577), .Y(n_1576) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1582), .Y(n_1581) );
INVx1_ASAP7_75t_L g1632 ( .A(n_1584), .Y(n_1632) );
INVx1_ASAP7_75t_L g1585 ( .A(n_1586), .Y(n_1585) );
OAI21xp33_ASAP7_75t_L g1587 ( .A1(n_1588), .A2(n_1589), .B(n_1591), .Y(n_1587) );
NOR2xp33_ASAP7_75t_L g1610 ( .A(n_1588), .B(n_1611), .Y(n_1610) );
INVx1_ASAP7_75t_L g1589 ( .A(n_1590), .Y(n_1589) );
INVx1_ASAP7_75t_L g1593 ( .A(n_1594), .Y(n_1593) );
NAND5xp2_ASAP7_75t_L g1597 ( .A(n_1598), .B(n_1604), .C(n_1614), .D(n_1623), .E(n_1635), .Y(n_1597) );
INVx1_ASAP7_75t_L g1599 ( .A(n_1600), .Y(n_1599) );
INVx1_ASAP7_75t_L g1621 ( .A(n_1600), .Y(n_1621) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1600), .Y(n_1639) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1606), .Y(n_1605) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1608), .Y(n_1607) );
INVx1_ASAP7_75t_L g1612 ( .A(n_1613), .Y(n_1612) );
NAND2xp5_ASAP7_75t_L g1615 ( .A(n_1616), .B(n_1617), .Y(n_1615) );
INVx1_ASAP7_75t_L g1619 ( .A(n_1620), .Y(n_1619) );
OR2x2_ASAP7_75t_L g1620 ( .A(n_1621), .B(n_1622), .Y(n_1620) );
INVxp67_ASAP7_75t_SL g1624 ( .A(n_1625), .Y(n_1624) );
INVxp67_ASAP7_75t_SL g1627 ( .A(n_1628), .Y(n_1627) );
INVx1_ASAP7_75t_L g1633 ( .A(n_1634), .Y(n_1633) );
O2A1O1Ixp33_ASAP7_75t_L g1635 ( .A1(n_1636), .A2(n_1637), .B(n_1641), .C(n_1643), .Y(n_1635) );
INVx1_ASAP7_75t_L g1637 ( .A(n_1638), .Y(n_1637) );
NAND2xp5_ASAP7_75t_L g1638 ( .A(n_1639), .B(n_1640), .Y(n_1638) );
INVx1_ASAP7_75t_L g1641 ( .A(n_1642), .Y(n_1641) );
INVx1_ASAP7_75t_L g1644 ( .A(n_1645), .Y(n_1644) );
INVxp67_ASAP7_75t_L g1646 ( .A(n_1647), .Y(n_1646) );
CKINVDCx5p33_ASAP7_75t_R g1648 ( .A(n_1649), .Y(n_1648) );
INVx1_ASAP7_75t_L g1649 ( .A(n_1650), .Y(n_1649) );
INVx1_ASAP7_75t_L g1650 ( .A(n_1651), .Y(n_1650) );
INVx1_ASAP7_75t_L g1694 ( .A(n_1654), .Y(n_1694) );
HB1xp67_ASAP7_75t_L g1654 ( .A(n_1655), .Y(n_1654) );
AND4x1_ASAP7_75t_L g1655 ( .A(n_1656), .B(n_1672), .C(n_1680), .D(n_1685), .Y(n_1655) );
OAI31xp33_ASAP7_75t_L g1656 ( .A1(n_1657), .A2(n_1664), .A3(n_1667), .B(n_1671), .Y(n_1656) );
NAND3xp33_ASAP7_75t_L g1657 ( .A(n_1658), .B(n_1660), .C(n_1663), .Y(n_1657) );
CKINVDCx14_ASAP7_75t_R g1695 ( .A(n_1696), .Y(n_1695) );
INVx2_ASAP7_75t_L g1696 ( .A(n_1697), .Y(n_1696) );
CKINVDCx5p33_ASAP7_75t_R g1697 ( .A(n_1698), .Y(n_1697) );
A2O1A1Ixp33_ASAP7_75t_L g1762 ( .A1(n_1699), .A2(n_1763), .B(n_1765), .C(n_1767), .Y(n_1762) );
BUFx2_ASAP7_75t_L g1701 ( .A(n_1702), .Y(n_1701) );
INVx1_ASAP7_75t_L g1702 ( .A(n_1703), .Y(n_1702) );
INVx1_ASAP7_75t_L g1703 ( .A(n_1704), .Y(n_1703) );
INVx1_ASAP7_75t_L g1705 ( .A(n_1706), .Y(n_1705) );
HB1xp67_ASAP7_75t_L g1706 ( .A(n_1707), .Y(n_1706) );
NOR2x1_ASAP7_75t_L g1708 ( .A(n_1709), .B(n_1732), .Y(n_1708) );
AOI21xp5_ASAP7_75t_L g1709 ( .A1(n_1710), .A2(n_1719), .B(n_1730), .Y(n_1709) );
AOI221xp5_ASAP7_75t_L g1710 ( .A1(n_1711), .A2(n_1712), .B1(n_1713), .B2(n_1715), .C(n_1717), .Y(n_1710) );
INVx2_ASAP7_75t_SL g1724 ( .A(n_1725), .Y(n_1724) );
INVx2_ASAP7_75t_L g1728 ( .A(n_1729), .Y(n_1728) );
INVx2_ASAP7_75t_L g1730 ( .A(n_1731), .Y(n_1730) );
NAND4xp25_ASAP7_75t_L g1732 ( .A(n_1733), .B(n_1739), .C(n_1743), .D(n_1748), .Y(n_1732) );
AOI221xp5_ASAP7_75t_L g1733 ( .A1(n_1734), .A2(n_1735), .B1(n_1736), .B2(n_1737), .C(n_1738), .Y(n_1733) );
AOI22xp5_ASAP7_75t_L g1743 ( .A1(n_1744), .A2(n_1745), .B1(n_1746), .B2(n_1747), .Y(n_1743) );
INVx1_ASAP7_75t_L g1757 ( .A(n_1758), .Y(n_1757) );
HB1xp67_ASAP7_75t_L g1761 ( .A(n_1762), .Y(n_1761) );
INVx1_ASAP7_75t_L g1763 ( .A(n_1764), .Y(n_1763) );
INVx1_ASAP7_75t_L g1765 ( .A(n_1766), .Y(n_1765) );
endmodule