module fake_netlist_6_4188_n_1678 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1678);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1678;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_544;
wire n_250;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_228;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_139),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_75),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_100),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_58),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_50),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_99),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_7),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_97),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_103),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_106),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_68),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_123),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_148),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_76),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_69),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_59),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_64),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_149),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_124),
.Y(n_172)
);

INVx4_ASAP7_75t_R g173 ( 
.A(n_34),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_114),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_25),
.Y(n_175)
);

BUFx10_ASAP7_75t_L g176 ( 
.A(n_47),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_129),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_40),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_50),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_105),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_74),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_115),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_19),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_78),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_30),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_51),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_136),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_85),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_62),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_12),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_138),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_55),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_93),
.Y(n_194)
);

BUFx10_ASAP7_75t_L g195 ( 
.A(n_18),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_26),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_144),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_72),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_33),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_88),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_135),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_11),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_16),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_27),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_134),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_104),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_66),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_48),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g209 ( 
.A(n_145),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_128),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_32),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_26),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_89),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_41),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_6),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_2),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_33),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_107),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_49),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_55),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_80),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_48),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_18),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_109),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_46),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_96),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_29),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_84),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_132),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_120),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_53),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_36),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_112),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_67),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_125),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_73),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_86),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_121),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_52),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_44),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_102),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_8),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_30),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_82),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_117),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_81),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_19),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_79),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_17),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_32),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_146),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_40),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_27),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_1),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_1),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_101),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_150),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_41),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_0),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_141),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_51),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_46),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_45),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_44),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_8),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_133),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_98),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_17),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_147),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_94),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_52),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_22),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_20),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_45),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_130),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_127),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_90),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_95),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_0),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_14),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_143),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_83),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_65),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_63),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_2),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_29),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_9),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_61),
.Y(n_288)
);

BUFx5_ASAP7_75t_L g289 ( 
.A(n_31),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_70),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_111),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_4),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_110),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_23),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_12),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_31),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_71),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_35),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_131),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_11),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_53),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_28),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_92),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_9),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_57),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

NOR2xp67_ASAP7_75t_L g307 ( 
.A(n_212),
.B(n_3),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_268),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_187),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_289),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_157),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_289),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_199),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_165),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_176),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_171),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_260),
.B(n_3),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_191),
.Y(n_318)
);

NOR2xp67_ASAP7_75t_L g319 ( 
.A(n_212),
.B(n_4),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_193),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g321 ( 
.A(n_181),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_235),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_162),
.B(n_5),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_289),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_289),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_289),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_176),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_289),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_289),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_184),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_184),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_196),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_186),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_186),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_219),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_153),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_162),
.B(n_5),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_219),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_190),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_175),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_180),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_192),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_208),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_168),
.B(n_6),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_155),
.Y(n_345)
);

NOR2xp67_ASAP7_75t_L g346 ( 
.A(n_216),
.B(n_7),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_202),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_176),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_209),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_152),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_233),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_203),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_195),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_204),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_214),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_256),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_195),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_240),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_215),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_257),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_185),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_220),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_153),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_167),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_231),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_211),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_217),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_195),
.Y(n_368)
);

INVxp33_ASAP7_75t_L g369 ( 
.A(n_222),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_225),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_188),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_240),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_249),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_197),
.Y(n_374)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_227),
.B(n_247),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_249),
.Y(n_376)
);

INVxp33_ASAP7_75t_L g377 ( 
.A(n_255),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_198),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_201),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_158),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_232),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_310),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_345),
.Y(n_383)
);

AND2x2_ASAP7_75t_SL g384 ( 
.A(n_344),
.B(n_244),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_306),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_310),
.Y(n_386)
);

NOR2x1_ASAP7_75t_L g387 ( 
.A(n_361),
.B(n_167),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_317),
.B(n_307),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_345),
.Y(n_389)
);

NAND2xp33_ASAP7_75t_L g390 ( 
.A(n_375),
.B(n_216),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_306),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_345),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_312),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_336),
.B(n_168),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_312),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_324),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_345),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_311),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_324),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_325),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_363),
.B(n_266),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_325),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_380),
.B(n_305),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_323),
.B(n_266),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_349),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_326),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_326),
.Y(n_407)
);

AND2x6_ASAP7_75t_L g408 ( 
.A(n_328),
.B(n_244),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_319),
.B(n_293),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_328),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_337),
.B(n_281),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_329),
.B(n_281),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_329),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_308),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_349),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_308),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_330),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_380),
.Y(n_418)
);

AND2x6_ASAP7_75t_L g419 ( 
.A(n_330),
.B(n_155),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_364),
.B(n_177),
.Y(n_420)
);

BUFx8_ASAP7_75t_L g421 ( 
.A(n_333),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_331),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_371),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_334),
.B(n_178),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_331),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_335),
.B(n_253),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_358),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_346),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_358),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_372),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_372),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_338),
.B(n_253),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_373),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_373),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_376),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_376),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_340),
.B(n_154),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_341),
.B(n_154),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_343),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_313),
.A2(n_252),
.B1(n_179),
.B2(n_302),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_309),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_366),
.Y(n_442)
);

INVx6_ASAP7_75t_L g443 ( 
.A(n_375),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_367),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_370),
.B(n_156),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_321),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_322),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_309),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_318),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_318),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_320),
.B(n_170),
.Y(n_451)
);

INVx4_ASAP7_75t_L g452 ( 
.A(n_405),
.Y(n_452)
);

OAI22xp33_ASAP7_75t_L g453 ( 
.A1(n_440),
.A2(n_258),
.B1(n_239),
.B2(n_279),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_451),
.B(n_350),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_385),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_385),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_392),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_382),
.Y(n_458)
);

BUFx10_ASAP7_75t_L g459 ( 
.A(n_451),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_404),
.B(n_320),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_404),
.B(n_411),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_391),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_392),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_394),
.B(n_369),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g465 ( 
.A(n_398),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_450),
.B(n_351),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_411),
.B(n_360),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g468 ( 
.A(n_443),
.Y(n_468)
);

AND2x6_ASAP7_75t_L g469 ( 
.A(n_412),
.B(n_155),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_392),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_388),
.B(n_374),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_L g472 ( 
.A1(n_384),
.A2(n_305),
.B1(n_286),
.B2(n_285),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_382),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_394),
.B(n_332),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_382),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_443),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_391),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_394),
.B(n_332),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_395),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_443),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_395),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_443),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_399),
.Y(n_483)
);

OR2x6_ASAP7_75t_L g484 ( 
.A(n_448),
.B(n_285),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_392),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_399),
.Y(n_486)
);

OAI21xp33_ASAP7_75t_SL g487 ( 
.A1(n_384),
.A2(n_264),
.B(n_263),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_443),
.Y(n_488)
);

CKINVDCx11_ASAP7_75t_R g489 ( 
.A(n_398),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_446),
.B(n_347),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_400),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_388),
.B(n_378),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_400),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_443),
.B(n_379),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_382),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_402),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_446),
.B(n_347),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_428),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_450),
.B(n_368),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_402),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_410),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_386),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_384),
.A2(n_286),
.B1(n_271),
.B2(n_294),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_410),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_386),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_413),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_413),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_392),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_439),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_403),
.B(n_355),
.Y(n_510)
);

BUFx10_ASAP7_75t_L g511 ( 
.A(n_450),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_386),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_446),
.B(n_447),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_392),
.Y(n_514)
);

AND3x2_ASAP7_75t_L g515 ( 
.A(n_414),
.B(n_327),
.C(n_315),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_428),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_386),
.Y(n_517)
);

AND2x2_ASAP7_75t_SL g518 ( 
.A(n_384),
.B(n_155),
.Y(n_518)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_405),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_446),
.B(n_352),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_415),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_415),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_450),
.B(n_352),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_393),
.Y(n_524)
);

NAND3xp33_ASAP7_75t_L g525 ( 
.A(n_418),
.B(n_359),
.C(n_354),
.Y(n_525)
);

AND3x2_ASAP7_75t_L g526 ( 
.A(n_414),
.B(n_353),
.C(n_348),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_403),
.Y(n_527)
);

OAI22xp33_ASAP7_75t_L g528 ( 
.A1(n_440),
.A2(n_274),
.B1(n_243),
.B2(n_272),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_393),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_403),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_448),
.A2(n_381),
.B1(n_365),
.B2(n_362),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_393),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_393),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_396),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_447),
.B(n_377),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_447),
.B(n_354),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_396),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_392),
.Y(n_538)
);

OR2x6_ASAP7_75t_L g539 ( 
.A(n_448),
.B(n_273),
.Y(n_539)
);

AND2x6_ASAP7_75t_L g540 ( 
.A(n_412),
.B(n_155),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_396),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_396),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_418),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_420),
.A2(n_447),
.B1(n_390),
.B2(n_412),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_406),
.Y(n_545)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_405),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_406),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_420),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_406),
.Y(n_549)
);

INVx1_ASAP7_75t_SL g550 ( 
.A(n_414),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_406),
.Y(n_551)
);

AND2x6_ASAP7_75t_L g552 ( 
.A(n_412),
.B(n_270),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_423),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_407),
.Y(n_554)
);

AND2x6_ASAP7_75t_L g555 ( 
.A(n_412),
.B(n_270),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_424),
.B(n_183),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_407),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_420),
.B(n_359),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_407),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_405),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_407),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_397),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_425),
.Y(n_563)
);

INVx5_ASAP7_75t_L g564 ( 
.A(n_408),
.Y(n_564)
);

OR2x6_ASAP7_75t_L g565 ( 
.A(n_448),
.B(n_280),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_425),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_420),
.B(n_362),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_439),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_420),
.A2(n_287),
.B1(n_304),
.B2(n_292),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_425),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_424),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_425),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_431),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_424),
.B(n_189),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_442),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g576 ( 
.A(n_401),
.B(n_357),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_387),
.Y(n_577)
);

INVx4_ASAP7_75t_L g578 ( 
.A(n_405),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_442),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_450),
.B(n_293),
.Y(n_580)
);

AND2x6_ASAP7_75t_L g581 ( 
.A(n_387),
.B(n_270),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_431),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_431),
.Y(n_583)
);

NAND3xp33_ASAP7_75t_L g584 ( 
.A(n_390),
.B(n_242),
.C(n_223),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_409),
.B(n_314),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_444),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_424),
.B(n_194),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_431),
.Y(n_588)
);

INVx5_ASAP7_75t_L g589 ( 
.A(n_408),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_424),
.Y(n_590)
);

OR2x6_ASAP7_75t_L g591 ( 
.A(n_409),
.B(n_296),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_SL g592 ( 
.A1(n_441),
.A2(n_356),
.B1(n_342),
.B2(n_339),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_397),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_444),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_397),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_461),
.B(n_401),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_548),
.B(n_518),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_535),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_548),
.B(n_405),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_544),
.B(n_405),
.Y(n_600)
);

OAI221xp5_ASAP7_75t_L g601 ( 
.A1(n_472),
.A2(n_445),
.B1(n_438),
.B2(n_437),
.C(n_200),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_513),
.B(n_437),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_460),
.B(n_441),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_518),
.B(n_438),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_577),
.B(n_449),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_577),
.B(n_449),
.Y(n_606)
);

INVxp67_ASAP7_75t_L g607 ( 
.A(n_510),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_468),
.B(n_445),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_467),
.B(n_416),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_456),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_571),
.B(n_426),
.Y(n_611)
);

OR2x6_ASAP7_75t_L g612 ( 
.A(n_539),
.B(n_426),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_535),
.B(n_416),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_464),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_568),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_568),
.Y(n_616)
);

INVxp33_ASAP7_75t_L g617 ( 
.A(n_510),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_468),
.B(n_417),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_575),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_482),
.B(n_417),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_482),
.B(n_417),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_490),
.B(n_416),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_503),
.A2(n_408),
.B1(n_205),
.B2(n_284),
.Y(n_623)
);

NOR2xp67_ASAP7_75t_L g624 ( 
.A(n_525),
.B(n_423),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_497),
.B(n_316),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_464),
.B(n_426),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_520),
.B(n_536),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_527),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_462),
.Y(n_629)
);

NOR3xp33_ASAP7_75t_L g630 ( 
.A(n_471),
.B(n_432),
.C(n_234),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g631 ( 
.A1(n_567),
.A2(n_218),
.B1(n_206),
.B2(n_210),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_462),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_488),
.B(n_417),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_527),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_488),
.B(n_476),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_476),
.B(n_417),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_571),
.B(n_432),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_530),
.B(n_432),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_575),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_590),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_480),
.B(n_434),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_480),
.B(n_477),
.Y(n_642)
);

INVx8_ASAP7_75t_L g643 ( 
.A(n_539),
.Y(n_643)
);

NAND2xp33_ASAP7_75t_L g644 ( 
.A(n_581),
.B(n_209),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_479),
.B(n_481),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_479),
.B(n_434),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_511),
.B(n_270),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_481),
.B(n_434),
.Y(n_648)
);

NAND3xp33_ASAP7_75t_L g649 ( 
.A(n_474),
.B(n_421),
.C(n_251),
.Y(n_649)
);

INVxp67_ASAP7_75t_SL g650 ( 
.A(n_457),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_511),
.B(n_288),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_483),
.B(n_486),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_579),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_483),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_579),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_486),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_586),
.Y(n_657)
);

NOR2xp67_ASAP7_75t_L g658 ( 
.A(n_492),
.B(n_422),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_SL g659 ( 
.A1(n_585),
.A2(n_259),
.B1(n_160),
.B2(n_302),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_586),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_491),
.B(n_434),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_491),
.B(n_434),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_530),
.B(n_422),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_576),
.B(n_421),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_498),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_509),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_493),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_590),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_493),
.B(n_408),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_478),
.A2(n_558),
.B1(n_565),
.B2(n_539),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_489),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_594),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_506),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_506),
.B(n_408),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_455),
.B(n_408),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_496),
.B(n_408),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_500),
.Y(n_677)
);

OR2x6_ASAP7_75t_L g678 ( 
.A(n_539),
.B(n_565),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_498),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_553),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_501),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_543),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_504),
.Y(n_683)
);

AO221x1_ASAP7_75t_L g684 ( 
.A1(n_453),
.A2(n_291),
.B1(n_288),
.B2(n_207),
.C(n_213),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_507),
.B(n_408),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_458),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_531),
.B(n_421),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_487),
.B(n_567),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_SL g689 ( 
.A1(n_459),
.A2(n_421),
.B1(n_265),
.B2(n_179),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_556),
.B(n_574),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_457),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_473),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_473),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_556),
.A2(n_408),
.B1(n_221),
.B2(n_230),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_556),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_574),
.B(n_288),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_574),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_581),
.B(n_408),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_587),
.B(n_288),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_587),
.B(n_291),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_581),
.B(n_408),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_587),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_484),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_459),
.B(n_156),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_484),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_581),
.B(n_383),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_484),
.Y(n_707)
);

INVxp67_ASAP7_75t_L g708 ( 
.A(n_543),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_484),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_523),
.B(n_291),
.Y(n_710)
);

BUFx12f_ASAP7_75t_SL g711 ( 
.A(n_591),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_581),
.B(n_383),
.Y(n_712)
);

OR2x2_ASAP7_75t_L g713 ( 
.A(n_550),
.B(n_158),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_563),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_581),
.B(n_383),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_475),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_565),
.B(n_383),
.Y(n_717)
);

NAND2xp33_ASAP7_75t_L g718 ( 
.A(n_469),
.B(n_209),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_459),
.B(n_159),
.Y(n_719)
);

INVxp67_ASAP7_75t_SL g720 ( 
.A(n_457),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_494),
.B(n_291),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_565),
.B(n_383),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_563),
.Y(n_723)
);

NAND2xp33_ASAP7_75t_L g724 ( 
.A(n_469),
.B(n_209),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_454),
.B(n_159),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_516),
.B(n_161),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_463),
.B(n_389),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_463),
.B(n_485),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_466),
.B(n_161),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_463),
.B(n_389),
.Y(n_730)
);

OAI21xp5_ASAP7_75t_L g731 ( 
.A1(n_524),
.A2(n_245),
.B(n_282),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_485),
.B(n_389),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_566),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_495),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_499),
.B(n_163),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_485),
.B(n_508),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_508),
.B(n_514),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_591),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_580),
.B(n_209),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_584),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_591),
.Y(n_741)
);

AOI221xp5_ASAP7_75t_L g742 ( 
.A1(n_528),
.A2(n_254),
.B1(n_223),
.B2(n_301),
.C(n_300),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_495),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_569),
.A2(n_283),
.B1(n_241),
.B2(n_303),
.Y(n_744)
);

O2A1O1Ixp33_ASAP7_75t_L g745 ( 
.A1(n_524),
.A2(n_436),
.B(n_430),
.C(n_429),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_SL g746 ( 
.A(n_465),
.B(n_163),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_529),
.B(n_427),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_533),
.B(n_209),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_591),
.B(n_164),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_529),
.B(n_427),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_604),
.B(n_452),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_600),
.A2(n_519),
.B(n_452),
.Y(n_752)
);

OAI21xp33_ASAP7_75t_L g753 ( 
.A1(n_603),
.A2(n_250),
.B(n_160),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_SL g754 ( 
.A(n_711),
.B(n_553),
.Y(n_754)
);

NOR3xp33_ASAP7_75t_L g755 ( 
.A(n_609),
.B(n_592),
.C(n_489),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_611),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_635),
.A2(n_519),
.B(n_452),
.Y(n_757)
);

O2A1O1Ixp33_ASAP7_75t_L g758 ( 
.A1(n_596),
.A2(n_549),
.B(n_532),
.C(n_542),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_613),
.B(n_515),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_611),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_599),
.A2(n_546),
.B(n_519),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_690),
.A2(n_560),
.B(n_546),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_614),
.B(n_164),
.Y(n_763)
);

OAI21xp5_ASAP7_75t_L g764 ( 
.A1(n_597),
.A2(n_542),
.B(n_532),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_627),
.B(n_545),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_614),
.Y(n_766)
);

NOR3xp33_ASAP7_75t_L g767 ( 
.A(n_625),
.B(n_297),
.C(n_267),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_690),
.A2(n_546),
.B(n_560),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_598),
.B(n_602),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_598),
.B(n_545),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_608),
.B(n_547),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_638),
.B(n_526),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_650),
.A2(n_578),
.B(n_560),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_617),
.B(n_547),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_611),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_640),
.B(n_578),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_720),
.A2(n_578),
.B(n_593),
.Y(n_777)
);

OAI21xp5_ASAP7_75t_L g778 ( 
.A1(n_597),
.A2(n_549),
.B(n_557),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_642),
.A2(n_595),
.B(n_593),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_658),
.B(n_554),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_622),
.B(n_554),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_688),
.A2(n_557),
.B1(n_172),
.B2(n_169),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_680),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_636),
.A2(n_595),
.B(n_593),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_637),
.B(n_429),
.Y(n_785)
);

NAND2x1_ASAP7_75t_L g786 ( 
.A(n_691),
.B(n_457),
.Y(n_786)
);

INVx3_ASAP7_75t_L g787 ( 
.A(n_640),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_637),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_637),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_617),
.B(n_533),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_607),
.B(n_534),
.Y(n_791)
);

NAND2xp33_ASAP7_75t_L g792 ( 
.A(n_640),
.B(n_469),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_626),
.B(n_534),
.Y(n_793)
);

NAND3xp33_ASAP7_75t_L g794 ( 
.A(n_742),
.B(n_725),
.C(n_719),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_610),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_SL g796 ( 
.A1(n_659),
.A2(n_250),
.B1(n_254),
.B2(n_259),
.Y(n_796)
);

NAND3xp33_ASAP7_75t_L g797 ( 
.A(n_704),
.B(n_248),
.C(n_246),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_615),
.B(n_537),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_688),
.A2(n_248),
.B1(n_169),
.B2(n_166),
.Y(n_799)
);

AND2x4_ASAP7_75t_SL g800 ( 
.A(n_680),
.B(n_457),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_616),
.B(n_537),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_610),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_682),
.B(n_541),
.Y(n_803)
);

A2O1A1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_601),
.A2(n_561),
.B(n_541),
.C(n_551),
.Y(n_804)
);

OR2x6_ASAP7_75t_L g805 ( 
.A(n_643),
.B(n_430),
.Y(n_805)
);

AOI21x1_ASAP7_75t_L g806 ( 
.A1(n_647),
.A2(n_551),
.B(n_559),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_619),
.B(n_559),
.Y(n_807)
);

CKINVDCx20_ASAP7_75t_R g808 ( 
.A(n_671),
.Y(n_808)
);

AOI22xp5_ASAP7_75t_L g809 ( 
.A1(n_670),
.A2(n_552),
.B1(n_540),
.B2(n_469),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_641),
.A2(n_595),
.B(n_593),
.Y(n_810)
);

A2O1A1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_735),
.A2(n_729),
.B(n_749),
.C(n_664),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_618),
.A2(n_595),
.B(n_593),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_663),
.B(n_436),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_640),
.B(n_166),
.Y(n_814)
);

OAI21xp33_ASAP7_75t_L g815 ( 
.A1(n_726),
.A2(n_262),
.B(n_300),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_620),
.A2(n_595),
.B(n_470),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_629),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_621),
.A2(n_470),
.B(n_538),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_633),
.A2(n_470),
.B(n_538),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_668),
.A2(n_687),
.B1(n_697),
.B2(n_695),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_740),
.A2(n_630),
.B1(n_702),
.B2(n_668),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_632),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_L g823 ( 
.A1(n_668),
.A2(n_174),
.B1(n_182),
.B2(n_172),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_639),
.B(n_502),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_653),
.B(n_655),
.Y(n_825)
);

OR2x2_ASAP7_75t_SL g826 ( 
.A(n_713),
.B(n_649),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_657),
.B(n_502),
.Y(n_827)
);

O2A1O1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_645),
.A2(n_652),
.B(n_606),
.C(n_605),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_728),
.A2(n_470),
.B(n_538),
.Y(n_829)
);

OAI21x1_ASAP7_75t_L g830 ( 
.A1(n_736),
.A2(n_517),
.B(n_512),
.Y(n_830)
);

NOR3xp33_ASAP7_75t_L g831 ( 
.A(n_605),
.B(n_297),
.C(n_182),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_660),
.B(n_505),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_691),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_737),
.A2(n_538),
.B(n_470),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_L g835 ( 
.A1(n_646),
.A2(n_661),
.B(n_648),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_654),
.B(n_521),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_691),
.Y(n_837)
);

NOR3xp33_ASAP7_75t_L g838 ( 
.A(n_606),
.B(n_299),
.C(n_174),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_647),
.A2(n_562),
.B(n_538),
.Y(n_839)
);

AND2x2_ASAP7_75t_SL g840 ( 
.A(n_644),
.B(n_570),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_651),
.A2(n_562),
.B(n_589),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_654),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_656),
.B(n_667),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_628),
.B(n_261),
.Y(n_844)
);

NOR2x1_ASAP7_75t_R g845 ( 
.A(n_671),
.B(n_261),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_651),
.A2(n_562),
.B(n_589),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_708),
.B(n_262),
.Y(n_847)
);

OAI21xp33_ASAP7_75t_L g848 ( 
.A1(n_746),
.A2(n_298),
.B(n_295),
.Y(n_848)
);

O2A1O1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_710),
.A2(n_572),
.B(n_588),
.C(n_583),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_691),
.A2(n_730),
.B(n_727),
.Y(n_850)
);

AOI21x1_ASAP7_75t_L g851 ( 
.A1(n_706),
.A2(n_715),
.B(n_712),
.Y(n_851)
);

INVxp67_ASAP7_75t_L g852 ( 
.A(n_665),
.Y(n_852)
);

AOI33xp33_ASAP7_75t_L g853 ( 
.A1(n_679),
.A2(n_265),
.A3(n_295),
.B1(n_298),
.B2(n_301),
.B3(n_433),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_673),
.B(n_564),
.Y(n_854)
);

A2O1A1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_673),
.A2(n_573),
.B(n_588),
.C(n_583),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_677),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_681),
.B(n_522),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_683),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_732),
.A2(n_589),
.B(n_564),
.Y(n_859)
);

AOI21xp33_ASAP7_75t_L g860 ( 
.A1(n_634),
.A2(n_246),
.B(n_251),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_684),
.A2(n_623),
.B1(n_721),
.B2(n_644),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_SL g862 ( 
.A(n_711),
.B(n_267),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_666),
.Y(n_863)
);

BUFx12f_ASAP7_75t_L g864 ( 
.A(n_612),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_672),
.B(n_433),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_631),
.B(n_299),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_686),
.Y(n_867)
);

OAI321xp33_ASAP7_75t_L g868 ( 
.A1(n_744),
.A2(n_173),
.A3(n_435),
.B1(n_433),
.B2(n_572),
.C(n_582),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_SL g869 ( 
.A(n_624),
.B(n_224),
.Y(n_869)
);

A2O1A1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_703),
.A2(n_582),
.B(n_277),
.C(n_276),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_662),
.B(n_555),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_686),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_705),
.B(n_555),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_675),
.B(n_209),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_741),
.B(n_226),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_L g876 ( 
.A1(n_678),
.A2(n_278),
.B1(n_228),
.B2(n_229),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_707),
.B(n_555),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_738),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_643),
.Y(n_879)
);

A2O1A1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_709),
.A2(n_290),
.B(n_236),
.C(n_237),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_717),
.A2(n_397),
.B(n_435),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_678),
.A2(n_238),
.B1(n_269),
.B2(n_275),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_738),
.Y(n_883)
);

INVx2_ASAP7_75t_SL g884 ( 
.A(n_739),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_722),
.A2(n_435),
.B(n_427),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_689),
.B(n_209),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_676),
.B(n_427),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_SL g888 ( 
.A(n_643),
.B(n_555),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_692),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_612),
.B(n_427),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_692),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_693),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_R g893 ( 
.A(n_643),
.B(n_118),
.Y(n_893)
);

OR2x2_ASAP7_75t_SL g894 ( 
.A(n_685),
.B(n_10),
.Y(n_894)
);

INVx3_ASAP7_75t_L g895 ( 
.A(n_693),
.Y(n_895)
);

AOI21x1_ASAP7_75t_L g896 ( 
.A1(n_669),
.A2(n_674),
.B(n_710),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_612),
.B(n_10),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_612),
.Y(n_898)
);

OAI22xp5_ASAP7_75t_L g899 ( 
.A1(n_678),
.A2(n_427),
.B1(n_469),
.B2(n_142),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_716),
.A2(n_419),
.B(n_140),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_678),
.B(n_13),
.Y(n_901)
);

A2O1A1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_745),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_731),
.A2(n_419),
.B(n_137),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_696),
.A2(n_419),
.B(n_126),
.Y(n_904)
);

NOR2x1p5_ASAP7_75t_L g905 ( 
.A(n_698),
.B(n_15),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_SL g906 ( 
.A(n_701),
.B(n_419),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_696),
.A2(n_16),
.B(n_20),
.C(n_21),
.Y(n_907)
);

OR2x2_ASAP7_75t_SL g908 ( 
.A(n_716),
.B(n_21),
.Y(n_908)
);

A2O1A1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_699),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_734),
.A2(n_419),
.B(n_122),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_739),
.A2(n_419),
.B1(n_119),
.B2(n_113),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_699),
.A2(n_419),
.B(n_91),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_743),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_714),
.B(n_24),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_811),
.A2(n_700),
.B1(n_694),
.B2(n_733),
.Y(n_915)
);

AOI221x1_ASAP7_75t_L g916 ( 
.A1(n_767),
.A2(n_820),
.B1(n_838),
.B2(n_831),
.C(n_755),
.Y(n_916)
);

O2A1O1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_767),
.A2(n_700),
.B(n_748),
.C(n_718),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_844),
.B(n_748),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_828),
.A2(n_723),
.B(n_724),
.C(n_718),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_769),
.B(n_750),
.Y(n_920)
);

OR2x6_ASAP7_75t_SL g921 ( 
.A(n_878),
.B(n_747),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_756),
.B(n_87),
.Y(n_922)
);

OR2x6_ASAP7_75t_L g923 ( 
.A(n_898),
.B(n_724),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_765),
.B(n_419),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_821),
.B(n_77),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_879),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_751),
.A2(n_60),
.B(n_419),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_852),
.B(n_25),
.Y(n_928)
);

AND2x6_ASAP7_75t_SL g929 ( 
.A(n_847),
.B(n_34),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_833),
.Y(n_930)
);

OA22x2_ASAP7_75t_L g931 ( 
.A1(n_753),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_817),
.Y(n_932)
);

O2A1O1Ixp5_ASAP7_75t_SL g933 ( 
.A1(n_886),
.A2(n_37),
.B(n_38),
.C(n_39),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_760),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_752),
.A2(n_57),
.B(n_43),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_822),
.Y(n_936)
);

AOI21xp33_ASAP7_75t_L g937 ( 
.A1(n_790),
.A2(n_42),
.B(n_43),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_902),
.A2(n_47),
.B(n_49),
.C(n_54),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_SL g939 ( 
.A1(n_808),
.A2(n_54),
.B1(n_56),
.B2(n_783),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_766),
.B(n_56),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_835),
.A2(n_804),
.B(n_840),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_813),
.B(n_774),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_831),
.A2(n_838),
.B(n_884),
.C(n_825),
.Y(n_943)
);

AOI21x1_ASAP7_75t_L g944 ( 
.A1(n_776),
.A2(n_806),
.B(n_843),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_777),
.A2(n_768),
.B(n_762),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_759),
.B(n_772),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_898),
.B(n_775),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_766),
.B(n_862),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_R g949 ( 
.A(n_883),
.B(n_754),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_861),
.A2(n_781),
.B1(n_840),
.B2(n_796),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_774),
.B(n_790),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_847),
.B(n_800),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_898),
.B(n_788),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_793),
.B(n_771),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_795),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_785),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_776),
.A2(n_757),
.B(n_761),
.Y(n_957)
);

AND2x2_ASAP7_75t_SL g958 ( 
.A(n_755),
.B(n_897),
.Y(n_958)
);

O2A1O1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_860),
.A2(n_866),
.B(n_909),
.C(n_907),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_779),
.A2(n_829),
.B(n_834),
.Y(n_960)
);

AND2x2_ASAP7_75t_SL g961 ( 
.A(n_897),
.B(n_901),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_864),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_879),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_799),
.A2(n_763),
.B(n_880),
.C(n_815),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_784),
.A2(n_810),
.B(n_850),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_802),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_826),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_842),
.B(n_791),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_R g969 ( 
.A(n_879),
.B(n_787),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_R g970 ( 
.A(n_879),
.B(n_787),
.Y(n_970)
);

NAND3xp33_ASAP7_75t_L g971 ( 
.A(n_796),
.B(n_875),
.C(n_797),
.Y(n_971)
);

BUFx12f_ASAP7_75t_L g972 ( 
.A(n_908),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_861),
.A2(n_863),
.B1(n_856),
.B2(n_858),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_791),
.B(n_770),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_870),
.A2(n_814),
.B(n_914),
.C(n_875),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_812),
.A2(n_816),
.B(n_818),
.Y(n_976)
);

NOR3xp33_ASAP7_75t_SL g977 ( 
.A(n_848),
.B(n_901),
.C(n_876),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_898),
.B(n_789),
.Y(n_978)
);

OR2x2_ASAP7_75t_L g979 ( 
.A(n_785),
.B(n_803),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_803),
.A2(n_914),
.B(n_865),
.C(n_868),
.Y(n_980)
);

OR2x6_ASAP7_75t_SL g981 ( 
.A(n_882),
.B(n_823),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_869),
.B(n_845),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_894),
.A2(n_805),
.B1(n_809),
.B2(n_899),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_865),
.B(n_780),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_867),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_758),
.A2(n_764),
.B(n_778),
.C(n_890),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_872),
.B(n_891),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_853),
.B(n_905),
.Y(n_988)
);

INVx5_ASAP7_75t_L g989 ( 
.A(n_833),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_893),
.B(n_833),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_892),
.B(n_913),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_805),
.A2(n_873),
.B1(n_877),
.B2(n_782),
.Y(n_992)
);

INVx1_ASAP7_75t_SL g993 ( 
.A(n_893),
.Y(n_993)
);

NOR3xp33_ASAP7_75t_SL g994 ( 
.A(n_874),
.B(n_854),
.C(n_904),
.Y(n_994)
);

AOI22xp5_ASAP7_75t_L g995 ( 
.A1(n_805),
.A2(n_874),
.B1(n_888),
.B2(n_854),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_819),
.A2(n_792),
.B(n_871),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_895),
.B(n_857),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_895),
.B(n_798),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_833),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_801),
.B(n_807),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_824),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_827),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_SL g1003 ( 
.A1(n_855),
.A2(n_887),
.B(n_910),
.C(n_900),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_832),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_836),
.A2(n_786),
.B(n_839),
.Y(n_1005)
);

OR2x6_ASAP7_75t_L g1006 ( 
.A(n_837),
.B(n_851),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_837),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_881),
.A2(n_849),
.B(n_885),
.C(n_903),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_896),
.Y(n_1009)
);

AND3x1_ASAP7_75t_SL g1010 ( 
.A(n_911),
.B(n_912),
.C(n_906),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_887),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_830),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_841),
.Y(n_1013)
);

OAI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_846),
.A2(n_604),
.B(n_518),
.Y(n_1014)
);

OAI22x1_ASAP7_75t_L g1015 ( 
.A1(n_859),
.A2(n_794),
.B1(n_603),
.B2(n_609),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_879),
.Y(n_1016)
);

A2O1A1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_794),
.A2(n_461),
.B(n_811),
.C(n_627),
.Y(n_1017)
);

INVx4_ASAP7_75t_L g1018 ( 
.A(n_879),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_769),
.B(n_596),
.Y(n_1019)
);

OR2x2_ASAP7_75t_L g1020 ( 
.A(n_783),
.B(n_510),
.Y(n_1020)
);

A2O1A1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_794),
.A2(n_461),
.B(n_811),
.C(n_627),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_879),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_794),
.A2(n_461),
.B1(n_596),
.B2(n_811),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_773),
.A2(n_600),
.B(n_548),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_844),
.B(n_613),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_773),
.A2(n_600),
.B(n_548),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_769),
.B(n_596),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_794),
.A2(n_461),
.B1(n_596),
.B2(n_811),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_844),
.B(n_613),
.Y(n_1029)
);

OAI21xp33_ASAP7_75t_L g1030 ( 
.A1(n_753),
.A2(n_461),
.B(n_603),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_794),
.B(n_603),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_833),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_773),
.A2(n_600),
.B(n_548),
.Y(n_1033)
);

HB1xp67_ASAP7_75t_L g1034 ( 
.A(n_852),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_794),
.A2(n_461),
.B1(n_601),
.B2(n_384),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_794),
.A2(n_461),
.B1(n_596),
.B2(n_811),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_769),
.B(n_596),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_769),
.B(n_596),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_773),
.A2(n_600),
.B(n_548),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_889),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_769),
.B(n_627),
.Y(n_1041)
);

OA22x2_ASAP7_75t_L g1042 ( 
.A1(n_753),
.A2(n_440),
.B1(n_607),
.B2(n_530),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_783),
.Y(n_1043)
);

O2A1O1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_811),
.A2(n_794),
.B(n_461),
.C(n_603),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_794),
.A2(n_461),
.B1(n_596),
.B2(n_811),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_844),
.B(n_613),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_1044),
.A2(n_1031),
.B(n_1030),
.C(n_1021),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_945),
.A2(n_957),
.B(n_1024),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_1026),
.A2(n_1039),
.B(n_1033),
.Y(n_1049)
);

INVx1_ASAP7_75t_SL g1050 ( 
.A(n_1020),
.Y(n_1050)
);

OAI22x1_ASAP7_75t_L g1051 ( 
.A1(n_971),
.A2(n_967),
.B1(n_948),
.B2(n_940),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_985),
.Y(n_1052)
);

OR2x2_ASAP7_75t_L g1053 ( 
.A(n_1025),
.B(n_1029),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_926),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_952),
.B(n_979),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_932),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_936),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_1019),
.B(n_1027),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_1041),
.B(n_1037),
.Y(n_1059)
);

HB1xp67_ASAP7_75t_L g1060 ( 
.A(n_1034),
.Y(n_1060)
);

AO31x2_ASAP7_75t_L g1061 ( 
.A1(n_1008),
.A2(n_1012),
.A3(n_986),
.B(n_950),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_996),
.A2(n_960),
.B(n_976),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_965),
.A2(n_1005),
.B(n_944),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_1041),
.B(n_1038),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_1017),
.A2(n_975),
.B(n_964),
.C(n_1035),
.Y(n_1065)
);

HB1xp67_ASAP7_75t_L g1066 ( 
.A(n_956),
.Y(n_1066)
);

OA21x2_ASAP7_75t_L g1067 ( 
.A1(n_941),
.A2(n_1014),
.B(n_919),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_1023),
.A2(n_1028),
.B1(n_1045),
.B2(n_1036),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_961),
.B(n_1046),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_941),
.A2(n_954),
.B(n_1003),
.Y(n_1070)
);

AOI221x1_ASAP7_75t_L g1071 ( 
.A1(n_1023),
.A2(n_1036),
.B1(n_1045),
.B2(n_1028),
.C(n_950),
.Y(n_1071)
);

OA21x2_ASAP7_75t_L g1072 ( 
.A1(n_1014),
.A2(n_1009),
.B(n_980),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_959),
.A2(n_977),
.B(n_943),
.C(n_917),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_954),
.A2(n_920),
.B(n_974),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_974),
.A2(n_915),
.B(n_1000),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_915),
.A2(n_942),
.B(n_951),
.Y(n_1076)
);

BUFx3_ASAP7_75t_L g1077 ( 
.A(n_1043),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_984),
.A2(n_997),
.B(n_998),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_946),
.B(n_958),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_992),
.A2(n_918),
.B(n_938),
.C(n_925),
.Y(n_1080)
);

BUFx10_ASAP7_75t_L g1081 ( 
.A(n_982),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_988),
.B(n_993),
.Y(n_1082)
);

OAI21xp5_ASAP7_75t_SL g1083 ( 
.A1(n_934),
.A2(n_916),
.B(n_937),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_927),
.A2(n_987),
.B(n_991),
.Y(n_1084)
);

AO31x2_ASAP7_75t_L g1085 ( 
.A1(n_1015),
.A2(n_983),
.A3(n_973),
.B(n_935),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_995),
.A2(n_947),
.B(n_978),
.Y(n_1086)
);

OAI21xp33_ASAP7_75t_SL g1087 ( 
.A1(n_1001),
.A2(n_1002),
.B(n_1004),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_968),
.A2(n_990),
.B(n_924),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_953),
.A2(n_973),
.B(n_983),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_993),
.B(n_949),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1011),
.B(n_955),
.Y(n_1091)
);

INVxp67_ASAP7_75t_L g1092 ( 
.A(n_928),
.Y(n_1092)
);

OA21x2_ASAP7_75t_L g1093 ( 
.A1(n_994),
.A2(n_966),
.B(n_937),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_923),
.A2(n_989),
.B(n_1006),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_923),
.A2(n_989),
.B(n_1006),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_962),
.Y(n_1096)
);

BUFx2_ASAP7_75t_L g1097 ( 
.A(n_972),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_981),
.A2(n_1042),
.B1(n_923),
.B2(n_931),
.Y(n_1098)
);

NAND2xp33_ASAP7_75t_SL g1099 ( 
.A(n_969),
.B(n_970),
.Y(n_1099)
);

NAND3xp33_ASAP7_75t_L g1100 ( 
.A(n_933),
.B(n_939),
.C(n_922),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_989),
.A2(n_1006),
.B(n_1013),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1040),
.Y(n_1102)
);

BUFx2_ASAP7_75t_L g1103 ( 
.A(n_921),
.Y(n_1103)
);

OAI21xp33_ASAP7_75t_L g1104 ( 
.A1(n_1042),
.A2(n_931),
.B(n_922),
.Y(n_1104)
);

AOI21xp33_ASAP7_75t_L g1105 ( 
.A1(n_1013),
.A2(n_999),
.B(n_1018),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_930),
.A2(n_1032),
.B(n_1013),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_926),
.A2(n_1016),
.B1(n_963),
.B2(n_1022),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1032),
.B(n_1007),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_926),
.A2(n_963),
.B1(n_1016),
.B2(n_1022),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_989),
.A2(n_1018),
.B(n_1010),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_963),
.A2(n_1016),
.B(n_1022),
.C(n_929),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_949),
.Y(n_1112)
);

OR2x2_ASAP7_75t_L g1113 ( 
.A(n_1020),
.B(n_465),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_1031),
.A2(n_811),
.B(n_1044),
.C(n_1021),
.Y(n_1114)
);

CKINVDCx20_ASAP7_75t_R g1115 ( 
.A(n_949),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1017),
.A2(n_1021),
.B(n_1044),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_945),
.A2(n_957),
.B(n_1024),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1019),
.B(n_1027),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_1044),
.A2(n_1031),
.B(n_794),
.C(n_811),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1017),
.A2(n_1021),
.B(n_1044),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_1044),
.A2(n_1031),
.B(n_794),
.C(n_811),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_949),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_996),
.A2(n_830),
.B(n_957),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_1031),
.B(n_311),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_945),
.A2(n_957),
.B(n_1024),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1031),
.A2(n_794),
.B1(n_625),
.B2(n_311),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1019),
.B(n_1027),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1019),
.B(n_1027),
.Y(n_1128)
);

NAND3xp33_ASAP7_75t_L g1129 ( 
.A(n_1031),
.B(n_794),
.C(n_1044),
.Y(n_1129)
);

AO32x2_ASAP7_75t_L g1130 ( 
.A1(n_1023),
.A2(n_1045),
.A3(n_1036),
.B1(n_1028),
.B2(n_950),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_996),
.A2(n_830),
.B(n_957),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1019),
.B(n_1027),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1019),
.B(n_1027),
.Y(n_1133)
);

A2O1A1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_1044),
.A2(n_1031),
.B(n_794),
.C(n_811),
.Y(n_1134)
);

NAND3xp33_ASAP7_75t_L g1135 ( 
.A(n_1031),
.B(n_794),
.C(n_1044),
.Y(n_1135)
);

O2A1O1Ixp5_ASAP7_75t_L g1136 ( 
.A1(n_1031),
.A2(n_811),
.B(n_1028),
.C(n_1023),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_1044),
.A2(n_1031),
.B(n_794),
.C(n_811),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_SL g1138 ( 
.A1(n_1031),
.A2(n_461),
.B(n_609),
.C(n_603),
.Y(n_1138)
);

NAND2x1p5_ASAP7_75t_L g1139 ( 
.A(n_989),
.B(n_1018),
.Y(n_1139)
);

NAND3xp33_ASAP7_75t_SL g1140 ( 
.A(n_1031),
.B(n_811),
.C(n_423),
.Y(n_1140)
);

AO31x2_ASAP7_75t_L g1141 ( 
.A1(n_1008),
.A2(n_1012),
.A3(n_986),
.B(n_950),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_945),
.A2(n_957),
.B(n_1024),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1019),
.B(n_1027),
.Y(n_1143)
);

BUFx2_ASAP7_75t_L g1144 ( 
.A(n_1034),
.Y(n_1144)
);

NOR2xp67_ASAP7_75t_L g1145 ( 
.A(n_1034),
.B(n_577),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1019),
.B(n_1027),
.Y(n_1146)
);

OAI21xp33_ASAP7_75t_L g1147 ( 
.A1(n_1031),
.A2(n_461),
.B(n_609),
.Y(n_1147)
);

INVx6_ASAP7_75t_L g1148 ( 
.A(n_962),
.Y(n_1148)
);

INVx3_ASAP7_75t_L g1149 ( 
.A(n_926),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1019),
.B(n_1027),
.Y(n_1150)
);

INVx3_ASAP7_75t_SL g1151 ( 
.A(n_1020),
.Y(n_1151)
);

OR2x2_ASAP7_75t_L g1152 ( 
.A(n_1020),
.B(n_465),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1019),
.B(n_1027),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_1031),
.B(n_311),
.Y(n_1154)
);

AO31x2_ASAP7_75t_L g1155 ( 
.A1(n_1008),
.A2(n_1012),
.A3(n_986),
.B(n_950),
.Y(n_1155)
);

OR2x2_ASAP7_75t_L g1156 ( 
.A(n_1020),
.B(n_465),
.Y(n_1156)
);

NOR2xp67_ASAP7_75t_SL g1157 ( 
.A(n_989),
.B(n_879),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_1034),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1017),
.A2(n_1021),
.B(n_1044),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_952),
.B(n_979),
.Y(n_1160)
);

AOI211xp5_ASAP7_75t_L g1161 ( 
.A1(n_1031),
.A2(n_794),
.B(n_603),
.C(n_609),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1031),
.B(n_311),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1031),
.A2(n_794),
.B1(n_971),
.B2(n_961),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1019),
.B(n_1027),
.Y(n_1164)
);

AO31x2_ASAP7_75t_L g1165 ( 
.A1(n_1008),
.A2(n_1012),
.A3(n_986),
.B(n_950),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1019),
.B(n_1027),
.Y(n_1166)
);

BUFx3_ASAP7_75t_L g1167 ( 
.A(n_1043),
.Y(n_1167)
);

INVx4_ASAP7_75t_SL g1168 ( 
.A(n_926),
.Y(n_1168)
);

AOI221x1_ASAP7_75t_L g1169 ( 
.A1(n_1023),
.A2(n_1036),
.B1(n_1045),
.B2(n_1028),
.C(n_811),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1017),
.A2(n_1021),
.B(n_1044),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_945),
.A2(n_957),
.B(n_1024),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1019),
.B(n_1027),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_945),
.A2(n_957),
.B(n_1024),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_996),
.A2(n_830),
.B(n_957),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1031),
.A2(n_794),
.B1(n_971),
.B2(n_961),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1019),
.B(n_1027),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_1008),
.A2(n_1012),
.A3(n_986),
.B(n_950),
.Y(n_1177)
);

OR2x6_ASAP7_75t_L g1178 ( 
.A(n_923),
.B(n_879),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1019),
.A2(n_1037),
.B1(n_1038),
.B2(n_1027),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_1044),
.A2(n_1031),
.B(n_794),
.C(n_811),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_945),
.A2(n_957),
.B(n_1024),
.Y(n_1181)
);

AO22x1_ASAP7_75t_L g1182 ( 
.A1(n_1124),
.A2(n_1154),
.B1(n_1162),
.B2(n_1122),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_L g1183 ( 
.A1(n_1147),
.A2(n_1175),
.B1(n_1163),
.B2(n_1135),
.Y(n_1183)
);

INVx6_ASAP7_75t_L g1184 ( 
.A(n_1168),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1129),
.A2(n_1135),
.B1(n_1068),
.B2(n_1140),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_1077),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1129),
.A2(n_1068),
.B1(n_1126),
.B2(n_1120),
.Y(n_1187)
);

CKINVDCx20_ASAP7_75t_R g1188 ( 
.A(n_1115),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1116),
.A2(n_1159),
.B1(n_1170),
.B2(n_1120),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1116),
.A2(n_1159),
.B1(n_1170),
.B2(n_1051),
.Y(n_1190)
);

BUFx3_ASAP7_75t_L g1191 ( 
.A(n_1167),
.Y(n_1191)
);

BUFx2_ASAP7_75t_L g1192 ( 
.A(n_1151),
.Y(n_1192)
);

BUFx3_ASAP7_75t_L g1193 ( 
.A(n_1144),
.Y(n_1193)
);

OAI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1058),
.A2(n_1150),
.B1(n_1143),
.B2(n_1146),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1098),
.A2(n_1104),
.B1(n_1069),
.B2(n_1179),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_1158),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_SL g1197 ( 
.A1(n_1098),
.A2(n_1079),
.B1(n_1100),
.B2(n_1103),
.Y(n_1197)
);

BUFx4f_ASAP7_75t_SL g1198 ( 
.A(n_1096),
.Y(n_1198)
);

OAI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1118),
.A2(n_1133),
.B1(n_1172),
.B2(n_1153),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1052),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1179),
.A2(n_1100),
.B1(n_1064),
.B2(n_1059),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_1178),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1132),
.A2(n_1176),
.B1(n_1127),
.B2(n_1164),
.Y(n_1203)
);

INVx1_ASAP7_75t_SL g1204 ( 
.A(n_1050),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1178),
.Y(n_1205)
);

BUFx12f_ASAP7_75t_L g1206 ( 
.A(n_1112),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1127),
.A2(n_1128),
.B1(n_1164),
.B2(n_1166),
.Y(n_1207)
);

BUFx12f_ASAP7_75t_L g1208 ( 
.A(n_1081),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1056),
.Y(n_1209)
);

BUFx3_ASAP7_75t_L g1210 ( 
.A(n_1148),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_SL g1211 ( 
.A1(n_1161),
.A2(n_1092),
.B1(n_1050),
.B2(n_1160),
.Y(n_1211)
);

BUFx4f_ASAP7_75t_L g1212 ( 
.A(n_1148),
.Y(n_1212)
);

CKINVDCx20_ASAP7_75t_R g1213 ( 
.A(n_1097),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_1139),
.Y(n_1214)
);

CKINVDCx20_ASAP7_75t_R g1215 ( 
.A(n_1081),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1128),
.A2(n_1166),
.B1(n_1076),
.B2(n_1070),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1075),
.A2(n_1074),
.B1(n_1067),
.B2(n_1053),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_SL g1218 ( 
.A1(n_1055),
.A2(n_1160),
.B1(n_1152),
.B2(n_1156),
.Y(n_1218)
);

INVx3_ASAP7_75t_SL g1219 ( 
.A(n_1113),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1091),
.Y(n_1220)
);

BUFx2_ASAP7_75t_SL g1221 ( 
.A(n_1145),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1139),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1066),
.Y(n_1223)
);

BUFx12f_ASAP7_75t_L g1224 ( 
.A(n_1111),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1119),
.B(n_1121),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1102),
.Y(n_1226)
);

CKINVDCx11_ASAP7_75t_R g1227 ( 
.A(n_1168),
.Y(n_1227)
);

CKINVDCx11_ASAP7_75t_R g1228 ( 
.A(n_1168),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1108),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1054),
.B(n_1149),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1067),
.A2(n_1089),
.B1(n_1093),
.B2(n_1071),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1087),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_1054),
.B(n_1149),
.Y(n_1233)
);

INVx4_ASAP7_75t_L g1234 ( 
.A(n_1157),
.Y(n_1234)
);

CKINVDCx20_ASAP7_75t_R g1235 ( 
.A(n_1090),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_SL g1236 ( 
.A(n_1099),
.Y(n_1236)
);

CKINVDCx11_ASAP7_75t_R g1237 ( 
.A(n_1136),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1106),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1134),
.B(n_1180),
.Y(n_1239)
);

AOI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1083),
.A2(n_1137),
.B1(n_1047),
.B2(n_1065),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_1086),
.Y(n_1241)
);

BUFx2_ASAP7_75t_L g1242 ( 
.A(n_1073),
.Y(n_1242)
);

BUFx10_ASAP7_75t_L g1243 ( 
.A(n_1105),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_SL g1244 ( 
.A1(n_1138),
.A2(n_1169),
.B1(n_1093),
.B2(n_1130),
.Y(n_1244)
);

BUFx2_ASAP7_75t_SL g1245 ( 
.A(n_1110),
.Y(n_1245)
);

BUFx12f_ASAP7_75t_L g1246 ( 
.A(n_1105),
.Y(n_1246)
);

BUFx8_ASAP7_75t_L g1247 ( 
.A(n_1130),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1114),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_1107),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1072),
.A2(n_1078),
.B1(n_1088),
.B2(n_1130),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1085),
.Y(n_1251)
);

BUFx2_ASAP7_75t_L g1252 ( 
.A(n_1085),
.Y(n_1252)
);

OAI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1094),
.A2(n_1095),
.B1(n_1101),
.B2(n_1072),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1080),
.Y(n_1254)
);

BUFx2_ASAP7_75t_SL g1255 ( 
.A(n_1109),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1048),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_SL g1257 ( 
.A1(n_1084),
.A2(n_1142),
.B1(n_1173),
.B2(n_1171),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1117),
.A2(n_1181),
.B1(n_1125),
.B2(n_1062),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1049),
.A2(n_1063),
.B1(n_1174),
.B2(n_1123),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1131),
.Y(n_1260)
);

CKINVDCx20_ASAP7_75t_R g1261 ( 
.A(n_1061),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1141),
.A2(n_1155),
.B1(n_1165),
.B2(n_1177),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1141),
.A2(n_1155),
.B1(n_1165),
.B2(n_1177),
.Y(n_1263)
);

CKINVDCx20_ASAP7_75t_R g1264 ( 
.A(n_1177),
.Y(n_1264)
);

INVx6_ASAP7_75t_L g1265 ( 
.A(n_1168),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_1115),
.Y(n_1266)
);

BUFx4f_ASAP7_75t_SL g1267 ( 
.A(n_1115),
.Y(n_1267)
);

BUFx12f_ASAP7_75t_L g1268 ( 
.A(n_1112),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1144),
.Y(n_1269)
);

INVx1_ASAP7_75t_SL g1270 ( 
.A(n_1050),
.Y(n_1270)
);

INVx2_ASAP7_75t_SL g1271 ( 
.A(n_1148),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1147),
.A2(n_1031),
.B1(n_1175),
.B2(n_1163),
.Y(n_1272)
);

INVx5_ASAP7_75t_L g1273 ( 
.A(n_1178),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1058),
.B(n_1118),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_SL g1275 ( 
.A1(n_1126),
.A2(n_1154),
.B(n_1124),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_SL g1276 ( 
.A1(n_1126),
.A2(n_1154),
.B(n_1124),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_SL g1277 ( 
.A1(n_1124),
.A2(n_1031),
.B1(n_1162),
.B2(n_1154),
.Y(n_1277)
);

INVx1_ASAP7_75t_SL g1278 ( 
.A(n_1050),
.Y(n_1278)
);

AOI22xp5_ASAP7_75t_SL g1279 ( 
.A1(n_1124),
.A2(n_1031),
.B1(n_1162),
.B2(n_1154),
.Y(n_1279)
);

INVxp67_ASAP7_75t_SL g1280 ( 
.A(n_1060),
.Y(n_1280)
);

INVx4_ASAP7_75t_SL g1281 ( 
.A(n_1178),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1058),
.B(n_1118),
.Y(n_1282)
);

OAI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1126),
.A2(n_794),
.B1(n_1031),
.B2(n_754),
.Y(n_1283)
);

BUFx4f_ASAP7_75t_SL g1284 ( 
.A(n_1115),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1057),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_1151),
.Y(n_1286)
);

AOI22xp5_ASAP7_75t_SL g1287 ( 
.A1(n_1124),
.A2(n_1031),
.B1(n_1162),
.B2(n_1154),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1082),
.B(n_961),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1147),
.A2(n_1031),
.B1(n_1175),
.B2(n_1163),
.Y(n_1289)
);

CKINVDCx11_ASAP7_75t_R g1290 ( 
.A(n_1115),
.Y(n_1290)
);

BUFx10_ASAP7_75t_L g1291 ( 
.A(n_1112),
.Y(n_1291)
);

INVxp67_ASAP7_75t_SL g1292 ( 
.A(n_1060),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1251),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1223),
.Y(n_1294)
);

INVx3_ASAP7_75t_L g1295 ( 
.A(n_1241),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_1290),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1189),
.A2(n_1258),
.B(n_1256),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1232),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1189),
.B(n_1207),
.Y(n_1299)
);

OA21x2_ASAP7_75t_L g1300 ( 
.A1(n_1231),
.A2(n_1250),
.B(n_1258),
.Y(n_1300)
);

BUFx2_ASAP7_75t_L g1301 ( 
.A(n_1261),
.Y(n_1301)
);

NAND2xp33_ASAP7_75t_R g1302 ( 
.A(n_1242),
.B(n_1254),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1281),
.B(n_1238),
.Y(n_1303)
);

AND2x4_ASAP7_75t_L g1304 ( 
.A(n_1281),
.B(n_1202),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1252),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1190),
.B(n_1264),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1207),
.B(n_1248),
.Y(n_1307)
);

OA21x2_ASAP7_75t_L g1308 ( 
.A1(n_1231),
.A2(n_1250),
.B(n_1262),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1190),
.B(n_1225),
.Y(n_1309)
);

CKINVDCx6p67_ASAP7_75t_R g1310 ( 
.A(n_1227),
.Y(n_1310)
);

OAI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1187),
.A2(n_1185),
.B(n_1289),
.Y(n_1311)
);

INVx3_ASAP7_75t_L g1312 ( 
.A(n_1260),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1187),
.A2(n_1289),
.B1(n_1272),
.B2(n_1203),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1203),
.B(n_1194),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1240),
.B(n_1244),
.Y(n_1315)
);

INVxp67_ASAP7_75t_L g1316 ( 
.A(n_1280),
.Y(n_1316)
);

HB1xp67_ASAP7_75t_L g1317 ( 
.A(n_1247),
.Y(n_1317)
);

BUFx2_ASAP7_75t_L g1318 ( 
.A(n_1247),
.Y(n_1318)
);

BUFx2_ASAP7_75t_L g1319 ( 
.A(n_1247),
.Y(n_1319)
);

OR2x2_ASAP7_75t_L g1320 ( 
.A(n_1239),
.B(n_1262),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1263),
.B(n_1185),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1200),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1209),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1259),
.A2(n_1217),
.B(n_1263),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1259),
.A2(n_1217),
.B(n_1216),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1246),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1292),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1272),
.A2(n_1183),
.B1(n_1283),
.B2(n_1237),
.Y(n_1328)
);

OA21x2_ASAP7_75t_L g1329 ( 
.A1(n_1216),
.A2(n_1201),
.B(n_1195),
.Y(n_1329)
);

CKINVDCx6p67_ASAP7_75t_R g1330 ( 
.A(n_1227),
.Y(n_1330)
);

OR2x2_ASAP7_75t_L g1331 ( 
.A(n_1201),
.B(n_1183),
.Y(n_1331)
);

BUFx6f_ASAP7_75t_L g1332 ( 
.A(n_1273),
.Y(n_1332)
);

INVxp67_ASAP7_75t_L g1333 ( 
.A(n_1220),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1253),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1195),
.A2(n_1205),
.B(n_1202),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1288),
.B(n_1237),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1281),
.B(n_1205),
.Y(n_1337)
);

INVxp67_ASAP7_75t_L g1338 ( 
.A(n_1269),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1285),
.Y(n_1339)
);

OR2x2_ASAP7_75t_L g1340 ( 
.A(n_1204),
.B(n_1278),
.Y(n_1340)
);

NOR2x1_ASAP7_75t_L g1341 ( 
.A(n_1245),
.B(n_1199),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1226),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_1290),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1274),
.B(n_1282),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1197),
.B(n_1229),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1246),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1243),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1222),
.A2(n_1257),
.B(n_1275),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1270),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1230),
.B(n_1233),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1196),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1276),
.A2(n_1277),
.B(n_1287),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1214),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1230),
.B(n_1233),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1214),
.Y(n_1355)
);

CKINVDCx6p67_ASAP7_75t_R g1356 ( 
.A(n_1310),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1352),
.B(n_1279),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1301),
.B(n_1219),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1344),
.B(n_1219),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1301),
.B(n_1193),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_SL g1361 ( 
.A1(n_1352),
.A2(n_1236),
.B(n_1234),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_1303),
.B(n_1295),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1298),
.Y(n_1363)
);

OA21x2_ASAP7_75t_L g1364 ( 
.A1(n_1325),
.A2(n_1233),
.B(n_1249),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1344),
.B(n_1182),
.Y(n_1365)
);

O2A1O1Ixp33_ASAP7_75t_SL g1366 ( 
.A1(n_1311),
.A2(n_1235),
.B(n_1215),
.C(n_1228),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1311),
.A2(n_1235),
.B(n_1192),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1327),
.B(n_1286),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1336),
.B(n_1186),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_SL g1370 ( 
.A(n_1296),
.B(n_1212),
.Y(n_1370)
);

AO21x2_ASAP7_75t_L g1371 ( 
.A1(n_1297),
.A2(n_1211),
.B(n_1224),
.Y(n_1371)
);

CKINVDCx20_ASAP7_75t_R g1372 ( 
.A(n_1343),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1314),
.B(n_1218),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1314),
.B(n_1236),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1313),
.B(n_1255),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1325),
.A2(n_1271),
.B(n_1234),
.Y(n_1376)
);

O2A1O1Ixp33_ASAP7_75t_L g1377 ( 
.A1(n_1313),
.A2(n_1331),
.B(n_1328),
.C(n_1297),
.Y(n_1377)
);

A2O1A1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1341),
.A2(n_1331),
.B(n_1315),
.C(n_1306),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1333),
.B(n_1191),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1322),
.B(n_1191),
.Y(n_1380)
);

NOR2x1_ASAP7_75t_SL g1381 ( 
.A(n_1332),
.B(n_1208),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1316),
.B(n_1221),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1345),
.B(n_1309),
.Y(n_1383)
);

OAI211xp5_ASAP7_75t_L g1384 ( 
.A1(n_1341),
.A2(n_1228),
.B(n_1210),
.C(n_1213),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1345),
.B(n_1208),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1310),
.A2(n_1213),
.B1(n_1212),
.B2(n_1188),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1336),
.B(n_1291),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1315),
.A2(n_1321),
.B1(n_1309),
.B2(n_1299),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1307),
.B(n_1184),
.Y(n_1389)
);

AOI221x1_ASAP7_75t_SL g1390 ( 
.A1(n_1307),
.A2(n_1291),
.B1(n_1198),
.B2(n_1206),
.C(n_1268),
.Y(n_1390)
);

OA21x2_ASAP7_75t_L g1391 ( 
.A1(n_1325),
.A2(n_1184),
.B(n_1265),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_SL g1392 ( 
.A(n_1310),
.B(n_1206),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1330),
.A2(n_1188),
.B1(n_1265),
.B2(n_1210),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1350),
.B(n_1268),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1354),
.B(n_1266),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1299),
.B(n_1265),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1346),
.B(n_1267),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_1316),
.B(n_1284),
.Y(n_1398)
);

OA21x2_ASAP7_75t_L g1399 ( 
.A1(n_1324),
.A2(n_1334),
.B(n_1348),
.Y(n_1399)
);

AO21x1_ASAP7_75t_L g1400 ( 
.A1(n_1302),
.A2(n_1339),
.B(n_1342),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1347),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_1330),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1330),
.A2(n_1346),
.B1(n_1326),
.B2(n_1329),
.Y(n_1403)
);

OAI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1348),
.A2(n_1329),
.B(n_1335),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1333),
.B(n_1294),
.Y(n_1405)
);

OR2x6_ASAP7_75t_L g1406 ( 
.A(n_1324),
.B(n_1335),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1321),
.A2(n_1319),
.B(n_1318),
.C(n_1317),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1303),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1322),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1406),
.B(n_1300),
.Y(n_1410)
);

AND2x4_ASAP7_75t_L g1411 ( 
.A(n_1408),
.B(n_1312),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1406),
.B(n_1300),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1401),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1406),
.B(n_1300),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1409),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1399),
.B(n_1305),
.Y(n_1416)
);

AND3x1_ASAP7_75t_SL g1417 ( 
.A(n_1357),
.B(n_1353),
.C(n_1355),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1363),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1357),
.A2(n_1329),
.B1(n_1349),
.B2(n_1320),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1376),
.Y(n_1420)
);

INVx1_ASAP7_75t_SL g1421 ( 
.A(n_1368),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1383),
.B(n_1322),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1399),
.Y(n_1423)
);

NOR2xp67_ASAP7_75t_L g1424 ( 
.A(n_1403),
.B(n_1295),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1405),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1400),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1372),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1404),
.B(n_1300),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1383),
.B(n_1323),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1364),
.B(n_1300),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1376),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1376),
.Y(n_1432)
);

OAI21xp5_ASAP7_75t_SL g1433 ( 
.A1(n_1377),
.A2(n_1337),
.B(n_1304),
.Y(n_1433)
);

NAND3xp33_ASAP7_75t_L g1434 ( 
.A(n_1375),
.B(n_1378),
.C(n_1388),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1391),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1391),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1418),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1434),
.A2(n_1375),
.B1(n_1367),
.B2(n_1371),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1423),
.Y(n_1439)
);

INVx5_ASAP7_75t_SL g1440 ( 
.A(n_1411),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1410),
.B(n_1391),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1423),
.Y(n_1442)
);

INVxp67_ASAP7_75t_L g1443 ( 
.A(n_1426),
.Y(n_1443)
);

AOI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1434),
.A2(n_1371),
.B1(n_1378),
.B2(n_1374),
.Y(n_1444)
);

NAND4xp25_ASAP7_75t_L g1445 ( 
.A(n_1419),
.B(n_1374),
.C(n_1365),
.D(n_1390),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1410),
.B(n_1362),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1415),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1410),
.B(n_1308),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1412),
.B(n_1308),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1422),
.B(n_1293),
.Y(n_1450)
);

INVx3_ASAP7_75t_SL g1451 ( 
.A(n_1427),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1431),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1415),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1412),
.B(n_1308),
.Y(n_1454)
);

INVx2_ASAP7_75t_SL g1455 ( 
.A(n_1411),
.Y(n_1455)
);

AND2x4_ASAP7_75t_SL g1456 ( 
.A(n_1411),
.B(n_1332),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1412),
.B(n_1308),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1414),
.B(n_1308),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1424),
.B(n_1407),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1413),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1429),
.B(n_1380),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1413),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1420),
.Y(n_1463)
);

INVxp67_ASAP7_75t_L g1464 ( 
.A(n_1426),
.Y(n_1464)
);

AND3x1_ASAP7_75t_L g1465 ( 
.A(n_1433),
.B(n_1392),
.C(n_1370),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1441),
.B(n_1414),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1447),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1441),
.B(n_1414),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1443),
.B(n_1416),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1441),
.B(n_1428),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1448),
.B(n_1428),
.Y(n_1471)
);

CKINVDCx16_ASAP7_75t_R g1472 ( 
.A(n_1444),
.Y(n_1472)
);

INVxp33_ASAP7_75t_L g1473 ( 
.A(n_1459),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1448),
.B(n_1428),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1448),
.B(n_1430),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1449),
.B(n_1430),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1455),
.B(n_1436),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1449),
.B(n_1430),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1449),
.B(n_1435),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1454),
.B(n_1435),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1439),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1447),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1443),
.B(n_1425),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1437),
.Y(n_1484)
);

INVx3_ASAP7_75t_L g1485 ( 
.A(n_1440),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1453),
.Y(n_1486)
);

NAND4xp25_ASAP7_75t_L g1487 ( 
.A(n_1444),
.B(n_1419),
.C(n_1373),
.D(n_1385),
.Y(n_1487)
);

AND2x4_ASAP7_75t_SL g1488 ( 
.A(n_1446),
.B(n_1356),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1439),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1464),
.B(n_1425),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1464),
.B(n_1416),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1439),
.Y(n_1492)
);

INVx2_ASAP7_75t_SL g1493 ( 
.A(n_1456),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1442),
.Y(n_1494)
);

AND2x4_ASAP7_75t_SL g1495 ( 
.A(n_1446),
.B(n_1356),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1463),
.B(n_1416),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1453),
.Y(n_1497)
);

INVxp67_ASAP7_75t_SL g1498 ( 
.A(n_1463),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1450),
.B(n_1429),
.Y(n_1499)
);

AND2x4_ASAP7_75t_SL g1500 ( 
.A(n_1446),
.B(n_1411),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1488),
.B(n_1440),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1467),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1467),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1488),
.B(n_1440),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1467),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1472),
.A2(n_1438),
.B1(n_1465),
.B2(n_1459),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1488),
.B(n_1440),
.Y(n_1507)
);

NOR3x1_ASAP7_75t_L g1508 ( 
.A(n_1487),
.B(n_1445),
.C(n_1384),
.Y(n_1508)
);

INVx1_ASAP7_75t_SL g1509 ( 
.A(n_1488),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1473),
.B(n_1451),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1496),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1482),
.Y(n_1512)
);

A2O1A1Ixp33_ASAP7_75t_L g1513 ( 
.A1(n_1473),
.A2(n_1438),
.B(n_1445),
.C(n_1433),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1482),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1472),
.B(n_1421),
.Y(n_1515)
);

INVx3_ASAP7_75t_L g1516 ( 
.A(n_1485),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1482),
.Y(n_1517)
);

OAI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1487),
.A2(n_1465),
.B(n_1424),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_SL g1519 ( 
.A(n_1485),
.B(n_1402),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1499),
.B(n_1460),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1486),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1486),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1496),
.Y(n_1523)
);

OAI21xp33_ASAP7_75t_L g1524 ( 
.A1(n_1499),
.A2(n_1458),
.B(n_1457),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1486),
.Y(n_1525)
);

INVx3_ASAP7_75t_L g1526 ( 
.A(n_1485),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1483),
.B(n_1460),
.Y(n_1527)
);

BUFx2_ASAP7_75t_L g1528 ( 
.A(n_1485),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1495),
.B(n_1455),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1497),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1483),
.B(n_1421),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1490),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1497),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1490),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1495),
.B(n_1440),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1469),
.B(n_1462),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1495),
.B(n_1440),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1497),
.Y(n_1538)
);

NOR2xp67_ASAP7_75t_L g1539 ( 
.A(n_1485),
.B(n_1455),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1496),
.Y(n_1540)
);

NOR2x1p5_ASAP7_75t_SL g1541 ( 
.A(n_1469),
.B(n_1452),
.Y(n_1541)
);

OAI32xp33_ASAP7_75t_L g1542 ( 
.A1(n_1469),
.A2(n_1420),
.A3(n_1432),
.B1(n_1457),
.B2(n_1458),
.Y(n_1542)
);

OAI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1493),
.A2(n_1385),
.B(n_1361),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1502),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1513),
.B(n_1471),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1501),
.B(n_1495),
.Y(n_1546)
);

NOR2xp67_ASAP7_75t_SL g1547 ( 
.A(n_1518),
.B(n_1402),
.Y(n_1547)
);

NOR2xp67_ASAP7_75t_L g1548 ( 
.A(n_1506),
.B(n_1493),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1510),
.B(n_1451),
.Y(n_1549)
);

OAI22xp33_ASAP7_75t_SL g1550 ( 
.A1(n_1515),
.A2(n_1498),
.B1(n_1491),
.B2(n_1451),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1501),
.B(n_1500),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1508),
.B(n_1471),
.Y(n_1552)
);

AND2x4_ASAP7_75t_SL g1553 ( 
.A(n_1529),
.B(n_1358),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1504),
.B(n_1500),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_L g1555 ( 
.A(n_1519),
.B(n_1451),
.Y(n_1555)
);

AOI32xp33_ASAP7_75t_L g1556 ( 
.A1(n_1509),
.A2(n_1358),
.A3(n_1386),
.B1(n_1457),
.B2(n_1458),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_SL g1557 ( 
.A(n_1543),
.B(n_1493),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1532),
.B(n_1471),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1534),
.B(n_1474),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1531),
.B(n_1474),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1504),
.B(n_1500),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1528),
.B(n_1474),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1528),
.B(n_1470),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1516),
.B(n_1372),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1507),
.B(n_1500),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_SL g1566 ( 
.A(n_1507),
.B(n_1393),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1529),
.B(n_1498),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1520),
.B(n_1470),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1535),
.B(n_1470),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1535),
.B(n_1466),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1537),
.B(n_1466),
.Y(n_1571)
);

XNOR2x2_ASAP7_75t_L g1572 ( 
.A(n_1536),
.B(n_1397),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1516),
.B(n_1387),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1520),
.B(n_1466),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1537),
.B(n_1468),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1527),
.B(n_1468),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1527),
.B(n_1468),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1524),
.B(n_1511),
.Y(n_1578)
);

AOI21xp33_ASAP7_75t_L g1579 ( 
.A1(n_1516),
.A2(n_1491),
.B(n_1359),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1552),
.B(n_1511),
.Y(n_1580)
);

OAI21xp5_ASAP7_75t_SL g1581 ( 
.A1(n_1545),
.A2(n_1556),
.B(n_1549),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1544),
.Y(n_1582)
);

O2A1O1Ixp33_ASAP7_75t_L g1583 ( 
.A1(n_1550),
.A2(n_1542),
.B(n_1366),
.C(n_1536),
.Y(n_1583)
);

XNOR2xp5_ASAP7_75t_L g1584 ( 
.A(n_1557),
.B(n_1572),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_L g1585 ( 
.A(n_1564),
.B(n_1526),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1550),
.A2(n_1548),
.B(n_1555),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1567),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1578),
.B(n_1523),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_SL g1589 ( 
.A(n_1548),
.B(n_1529),
.Y(n_1589)
);

AOI32xp33_ASAP7_75t_L g1590 ( 
.A1(n_1572),
.A2(n_1526),
.A3(n_1479),
.B1(n_1480),
.B2(n_1523),
.Y(n_1590)
);

INVx1_ASAP7_75t_SL g1591 ( 
.A(n_1546),
.Y(n_1591)
);

AOI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1566),
.A2(n_1539),
.B1(n_1526),
.B2(n_1389),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1567),
.B(n_1540),
.Y(n_1593)
);

INVx2_ASAP7_75t_SL g1594 ( 
.A(n_1553),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1544),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1567),
.B(n_1540),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1570),
.Y(n_1597)
);

AOI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1556),
.A2(n_1366),
.B(n_1542),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_SL g1599 ( 
.A(n_1546),
.B(n_1440),
.Y(n_1599)
);

AOI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1579),
.A2(n_1491),
.B(n_1397),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1562),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1576),
.B(n_1461),
.Y(n_1602)
);

AOI21xp33_ASAP7_75t_SL g1603 ( 
.A1(n_1573),
.A2(n_1369),
.B(n_1398),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1563),
.Y(n_1604)
);

INVx1_ASAP7_75t_SL g1605 ( 
.A(n_1591),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1582),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1587),
.B(n_1553),
.Y(n_1607)
);

AOI221xp5_ASAP7_75t_L g1608 ( 
.A1(n_1590),
.A2(n_1547),
.B1(n_1577),
.B2(n_1559),
.C(n_1558),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1594),
.B(n_1551),
.Y(n_1609)
);

AOI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1584),
.A2(n_1547),
.B1(n_1551),
.B2(n_1554),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1595),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1581),
.B(n_1569),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1586),
.A2(n_1574),
.B1(n_1568),
.B2(n_1560),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1580),
.B(n_1569),
.Y(n_1614)
);

OAI221xp5_ASAP7_75t_L g1615 ( 
.A1(n_1586),
.A2(n_1565),
.B1(n_1561),
.B2(n_1554),
.C(n_1575),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1589),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1601),
.B(n_1570),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1604),
.B(n_1571),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1593),
.Y(n_1619)
);

O2A1O1Ixp33_ASAP7_75t_L g1620 ( 
.A1(n_1583),
.A2(n_1575),
.B(n_1571),
.C(n_1565),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1596),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1598),
.A2(n_1561),
.B1(n_1329),
.B2(n_1396),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1597),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1605),
.B(n_1612),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1623),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1623),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1609),
.B(n_1585),
.Y(n_1627)
);

XNOR2x2_ASAP7_75t_L g1628 ( 
.A(n_1610),
.B(n_1598),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1609),
.B(n_1603),
.Y(n_1629)
);

AOI222xp33_ASAP7_75t_L g1630 ( 
.A1(n_1613),
.A2(n_1541),
.B1(n_1599),
.B2(n_1583),
.C1(n_1600),
.C2(n_1480),
.Y(n_1630)
);

NOR4xp25_ASAP7_75t_L g1631 ( 
.A(n_1606),
.B(n_1588),
.C(n_1602),
.D(n_1502),
.Y(n_1631)
);

XOR2x2_ASAP7_75t_SL g1632 ( 
.A(n_1614),
.B(n_1592),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_SL g1633 ( 
.A(n_1622),
.B(n_1600),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1619),
.B(n_1541),
.Y(n_1634)
);

NAND2xp33_ASAP7_75t_SL g1635 ( 
.A(n_1633),
.B(n_1627),
.Y(n_1635)
);

NOR3xp33_ASAP7_75t_L g1636 ( 
.A(n_1624),
.B(n_1616),
.C(n_1621),
.Y(n_1636)
);

AOI21xp5_ASAP7_75t_L g1637 ( 
.A1(n_1631),
.A2(n_1620),
.B(n_1622),
.Y(n_1637)
);

NOR3x1_ASAP7_75t_L g1638 ( 
.A(n_1629),
.B(n_1615),
.C(n_1617),
.Y(n_1638)
);

NOR3xp33_ASAP7_75t_L g1639 ( 
.A(n_1625),
.B(n_1618),
.C(n_1608),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1626),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1631),
.B(n_1607),
.Y(n_1641)
);

INVxp67_ASAP7_75t_L g1642 ( 
.A(n_1628),
.Y(n_1642)
);

OAI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1630),
.A2(n_1607),
.B(n_1611),
.Y(n_1643)
);

NOR3xp33_ASAP7_75t_SL g1644 ( 
.A(n_1634),
.B(n_1379),
.C(n_1407),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1632),
.B(n_1479),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1642),
.B(n_1351),
.Y(n_1646)
);

OAI211xp5_ASAP7_75t_L g1647 ( 
.A1(n_1637),
.A2(n_1338),
.B(n_1533),
.C(n_1530),
.Y(n_1647)
);

AOI221xp5_ASAP7_75t_L g1648 ( 
.A1(n_1639),
.A2(n_1538),
.B1(n_1533),
.B2(n_1530),
.C(n_1525),
.Y(n_1648)
);

NOR3xp33_ASAP7_75t_SL g1649 ( 
.A(n_1635),
.B(n_1505),
.C(n_1503),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1640),
.Y(n_1650)
);

OAI222xp33_ASAP7_75t_L g1651 ( 
.A1(n_1645),
.A2(n_1538),
.B1(n_1525),
.B2(n_1522),
.C1(n_1521),
.C2(n_1517),
.Y(n_1651)
);

NAND3xp33_ASAP7_75t_L g1652 ( 
.A(n_1649),
.B(n_1636),
.C(n_1641),
.Y(n_1652)
);

AOI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1646),
.A2(n_1643),
.B1(n_1644),
.B2(n_1638),
.Y(n_1653)
);

AOI221xp5_ASAP7_75t_L g1654 ( 
.A1(n_1647),
.A2(n_1512),
.B1(n_1521),
.B2(n_1517),
.C(n_1514),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1650),
.Y(n_1655)
);

AOI211xp5_ASAP7_75t_L g1656 ( 
.A1(n_1651),
.A2(n_1338),
.B(n_1360),
.C(n_1340),
.Y(n_1656)
);

AOI221xp5_ASAP7_75t_SL g1657 ( 
.A1(n_1648),
.A2(n_1522),
.B1(n_1514),
.B2(n_1512),
.C(n_1505),
.Y(n_1657)
);

NAND4xp75_ASAP7_75t_L g1658 ( 
.A(n_1655),
.B(n_1503),
.C(n_1479),
.D(n_1480),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1652),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1653),
.B(n_1395),
.Y(n_1660)
);

NAND4xp75_ASAP7_75t_L g1661 ( 
.A(n_1657),
.B(n_1478),
.C(n_1476),
.D(n_1475),
.Y(n_1661)
);

A2O1A1Ixp33_ASAP7_75t_L g1662 ( 
.A1(n_1656),
.A2(n_1477),
.B(n_1326),
.C(n_1492),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1659),
.B(n_1475),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1660),
.B(n_1654),
.Y(n_1664)
);

AO211x2_ASAP7_75t_L g1665 ( 
.A1(n_1658),
.A2(n_1484),
.B(n_1355),
.C(n_1353),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1663),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1666),
.Y(n_1667)
);

XNOR2xp5_ASAP7_75t_L g1668 ( 
.A(n_1667),
.B(n_1664),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1667),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1669),
.A2(n_1665),
.B1(n_1661),
.B2(n_1662),
.Y(n_1670)
);

CKINVDCx20_ASAP7_75t_R g1671 ( 
.A(n_1668),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1671),
.A2(n_1394),
.B(n_1481),
.Y(n_1672)
);

AOI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1670),
.A2(n_1477),
.B1(n_1494),
.B2(n_1492),
.Y(n_1673)
);

XOR2xp5_ASAP7_75t_L g1674 ( 
.A(n_1673),
.B(n_1381),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1674),
.B(n_1672),
.Y(n_1675)
);

OR3x2_ASAP7_75t_L g1676 ( 
.A(n_1675),
.B(n_1382),
.C(n_1326),
.Y(n_1676)
);

OAI221xp5_ASAP7_75t_R g1677 ( 
.A1(n_1676),
.A2(n_1417),
.B1(n_1494),
.B2(n_1492),
.C(n_1489),
.Y(n_1677)
);

AOI211xp5_ASAP7_75t_L g1678 ( 
.A1(n_1677),
.A2(n_1494),
.B(n_1492),
.C(n_1489),
.Y(n_1678)
);


endmodule