module fake_aes_12696_n_638 (n_117, n_44, n_133, n_149, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_125, n_9, n_161, n_10, n_177, n_130, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_169, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_46, n_31, n_58, n_122, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_182, n_166, n_162, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_638);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_125;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_169;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_182;
input n_166;
input n_162;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_638;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_431;
wire n_484;
wire n_496;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_612;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_627;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_202;
wire n_386;
wire n_432;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_205;
wire n_330;
wire n_587;
wire n_387;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_616;
wire n_365;
wire n_541;
wire n_315;
wire n_363;
wire n_409;
wire n_295;
wire n_263;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_553;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_524;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_602;
wire n_198;
wire n_424;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_187;
wire n_375;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_444;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_421;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g184 ( .A(n_157), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_137), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_160), .Y(n_186) );
NOR2xp67_ASAP7_75t_L g187 ( .A(n_131), .B(n_168), .Y(n_187) );
INVx1_ASAP7_75t_SL g188 ( .A(n_99), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_152), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_70), .Y(n_190) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_144), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_32), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_62), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_163), .Y(n_194) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_14), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_151), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_78), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_178), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_123), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_57), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_139), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_33), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_29), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_48), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_27), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_155), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_83), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_45), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_95), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_34), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_162), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_7), .B(n_81), .Y(n_212) );
INVxp33_ASAP7_75t_L g213 ( .A(n_135), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_119), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_107), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_126), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_42), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_60), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_24), .B(n_171), .Y(n_219) );
INVx1_ASAP7_75t_SL g220 ( .A(n_5), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_0), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_117), .Y(n_222) );
INVx3_ASAP7_75t_L g223 ( .A(n_146), .Y(n_223) );
INVx1_ASAP7_75t_SL g224 ( .A(n_100), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_8), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_143), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_127), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_61), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_36), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_102), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_149), .Y(n_231) );
CKINVDCx14_ASAP7_75t_R g232 ( .A(n_132), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_170), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_133), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_141), .Y(n_235) );
INVx2_ASAP7_75t_SL g236 ( .A(n_31), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_72), .Y(n_237) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_35), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_65), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_121), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_20), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_158), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_88), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_91), .Y(n_244) );
CKINVDCx16_ASAP7_75t_R g245 ( .A(n_93), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_74), .Y(n_246) );
NOR2xp67_ASAP7_75t_L g247 ( .A(n_159), .B(n_90), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_174), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_136), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g250 ( .A(n_82), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_71), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_53), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_147), .Y(n_253) );
BUFx10_ASAP7_75t_L g254 ( .A(n_5), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_43), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_76), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_150), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_118), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_59), .Y(n_259) );
INVx2_ASAP7_75t_SL g260 ( .A(n_175), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_86), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_124), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_172), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_148), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_105), .Y(n_265) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_154), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_129), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_56), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_109), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_75), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_130), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_166), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_145), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_25), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_116), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_38), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_26), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_161), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_177), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_169), .Y(n_280) );
CKINVDCx20_ASAP7_75t_R g281 ( .A(n_8), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_51), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_110), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_128), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_167), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_89), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_6), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_111), .Y(n_288) );
CKINVDCx16_ASAP7_75t_R g289 ( .A(n_58), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_153), .B(n_156), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_46), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_14), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_39), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_73), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_164), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_108), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_40), .Y(n_297) );
INVx1_ASAP7_75t_SL g298 ( .A(n_165), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_142), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_176), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_173), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_179), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_225), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_213), .B(n_0), .Y(n_304) );
AOI22x1_ASAP7_75t_SL g305 ( .A1(n_281), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_305) );
NOR2x1_ASAP7_75t_L g306 ( .A(n_223), .B(n_18), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_287), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_254), .Y(n_308) );
AND2x4_ASAP7_75t_L g309 ( .A(n_223), .B(n_1), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_236), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_292), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_184), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_203), .Y(n_313) );
CKINVDCx14_ASAP7_75t_R g314 ( .A(n_232), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_260), .Y(n_315) );
AOI22xp33_ASAP7_75t_SL g316 ( .A1(n_220), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_185), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_190), .B(n_4), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_186), .Y(n_319) );
INVx5_ASAP7_75t_L g320 ( .A(n_203), .Y(n_320) );
AND2x2_ASAP7_75t_SL g321 ( .A(n_245), .B(n_19), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_199), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_196), .Y(n_323) );
BUFx8_ASAP7_75t_L g324 ( .A(n_212), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_197), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_198), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_289), .B(n_6), .Y(n_327) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_203), .Y(n_328) );
INVxp67_ASAP7_75t_SL g329 ( .A(n_327), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_322), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_312), .B(n_218), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_320), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g333 ( .A1(n_321), .A2(n_221), .B1(n_195), .B2(n_230), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_314), .Y(n_334) );
CKINVDCx6p67_ASAP7_75t_R g335 ( .A(n_321), .Y(n_335) );
NAND3xp33_ASAP7_75t_L g336 ( .A(n_304), .B(n_302), .C(n_208), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_309), .B(n_227), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_320), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_316), .A2(n_250), .B1(n_288), .B2(n_220), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_320), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_309), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_320), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_318), .Y(n_343) );
NAND2xp5_ASAP7_75t_SL g344 ( .A(n_308), .B(n_189), .Y(n_344) );
INVx3_ASAP7_75t_L g345 ( .A(n_318), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_317), .B(n_233), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_319), .B(n_271), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_329), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_329), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_334), .Y(n_350) );
INVx2_ASAP7_75t_SL g351 ( .A(n_341), .Y(n_351) );
NAND2xp5_ASAP7_75t_SL g352 ( .A(n_336), .B(n_324), .Y(n_352) );
A2O1A1Ixp33_ASAP7_75t_L g353 ( .A1(n_343), .A2(n_345), .B(n_346), .C(n_331), .Y(n_353) );
INVxp67_ASAP7_75t_L g354 ( .A(n_331), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_337), .B(n_314), .Y(n_355) );
NAND2xp5_ASAP7_75t_SL g356 ( .A(n_337), .B(n_310), .Y(n_356) );
BUFx3_ASAP7_75t_L g357 ( .A(n_330), .Y(n_357) );
INVx2_ASAP7_75t_SL g358 ( .A(n_346), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_344), .B(n_323), .Y(n_359) );
OAI22xp5_ASAP7_75t_L g360 ( .A1(n_335), .A2(n_316), .B1(n_307), .B2(n_311), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_333), .B(n_254), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_347), .B(n_325), .Y(n_362) );
NAND2xp33_ASAP7_75t_L g363 ( .A(n_347), .B(n_290), .Y(n_363) );
AND2x4_ASAP7_75t_L g364 ( .A(n_332), .B(n_315), .Y(n_364) );
NAND2xp33_ASAP7_75t_L g365 ( .A(n_338), .B(n_306), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_339), .B(n_326), .Y(n_366) );
INVx8_ASAP7_75t_L g367 ( .A(n_339), .Y(n_367) );
CKINVDCx10_ASAP7_75t_R g368 ( .A(n_350), .Y(n_368) );
NOR2xp33_ASAP7_75t_R g369 ( .A(n_367), .B(n_191), .Y(n_369) );
AOI21xp5_ASAP7_75t_L g370 ( .A1(n_363), .A2(n_342), .B(n_340), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_357), .Y(n_371) );
NAND3xp33_ASAP7_75t_L g372 ( .A(n_366), .B(n_305), .C(n_303), .Y(n_372) );
O2A1O1Ixp33_ASAP7_75t_L g373 ( .A1(n_360), .A2(n_209), .B(n_210), .C(n_204), .Y(n_373) );
AOI21xp5_ASAP7_75t_L g374 ( .A1(n_353), .A2(n_222), .B(n_216), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_354), .B(n_224), .Y(n_375) );
A2O1A1Ixp33_ASAP7_75t_L g376 ( .A1(n_348), .A2(n_239), .B(n_242), .C(n_240), .Y(n_376) );
NAND2xp5_ASAP7_75t_SL g377 ( .A(n_358), .B(n_192), .Y(n_377) );
CKINVDCx8_ASAP7_75t_R g378 ( .A(n_367), .Y(n_378) );
O2A1O1Ixp33_ASAP7_75t_L g379 ( .A1(n_360), .A2(n_243), .B(n_248), .C(n_246), .Y(n_379) );
AO21x2_ASAP7_75t_L g380 ( .A1(n_365), .A2(n_253), .B(n_251), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_349), .Y(n_381) );
NAND2xp5_ASAP7_75t_SL g382 ( .A(n_351), .B(n_193), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_352), .B(n_255), .Y(n_383) );
OAI22xp5_ASAP7_75t_L g384 ( .A1(n_362), .A2(n_261), .B1(n_262), .B2(n_256), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_359), .B(n_194), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_367), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_361), .B(n_7), .Y(n_387) );
O2A1O1Ixp33_ASAP7_75t_L g388 ( .A1(n_356), .A2(n_275), .B(n_279), .C(n_278), .Y(n_388) );
AOI21xp5_ASAP7_75t_L g389 ( .A1(n_355), .A2(n_267), .B(n_263), .Y(n_389) );
AOI221x1_ASAP7_75t_L g390 ( .A1(n_374), .A2(n_286), .B1(n_268), .B2(n_273), .C(n_277), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_375), .B(n_364), .Y(n_391) );
A2O1A1Ixp33_ASAP7_75t_L g392 ( .A1(n_373), .A2(n_379), .B(n_389), .C(n_388), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_381), .B(n_364), .Y(n_393) );
OAI21xp5_ASAP7_75t_L g394 ( .A1(n_376), .A2(n_301), .B(n_247), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_371), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_387), .B(n_283), .Y(n_396) );
BUFx2_ASAP7_75t_L g397 ( .A(n_369), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_384), .B(n_200), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_384), .B(n_284), .Y(n_399) );
OAI21x1_ASAP7_75t_L g400 ( .A1(n_382), .A2(n_285), .B(n_187), .Y(n_400) );
AO21x1_ASAP7_75t_L g401 ( .A1(n_383), .A2(n_219), .B(n_313), .Y(n_401) );
AOI21xp5_ASAP7_75t_L g402 ( .A1(n_385), .A2(n_298), .B(n_188), .Y(n_402) );
AOI21xp5_ASAP7_75t_L g403 ( .A1(n_377), .A2(n_202), .B(n_201), .Y(n_403) );
OAI21xp5_ASAP7_75t_L g404 ( .A1(n_383), .A2(n_206), .B(n_205), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_372), .B(n_9), .Y(n_405) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_380), .A2(n_211), .B(n_207), .Y(n_406) );
AO31x2_ASAP7_75t_L g407 ( .A1(n_380), .A2(n_328), .A3(n_313), .B(n_266), .Y(n_407) );
OAI21xp5_ASAP7_75t_L g408 ( .A1(n_386), .A2(n_215), .B(n_214), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_378), .B(n_226), .Y(n_409) );
O2A1O1Ixp5_ASAP7_75t_L g410 ( .A1(n_368), .A2(n_265), .B(n_228), .C(n_300), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_381), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_378), .A2(n_266), .B1(n_229), .B2(n_258), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_381), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_381), .Y(n_414) );
OAI21x1_ASAP7_75t_L g415 ( .A1(n_370), .A2(n_229), .B(n_217), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_391), .B(n_9), .Y(n_416) );
BUFx3_ASAP7_75t_L g417 ( .A(n_397), .Y(n_417) );
OAI21x1_ASAP7_75t_SL g418 ( .A1(n_401), .A2(n_10), .B(n_11), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_414), .Y(n_419) );
OAI221xp5_ASAP7_75t_L g420 ( .A1(n_392), .A2(n_266), .B1(n_258), .B2(n_217), .C(n_297), .Y(n_420) );
AND2x6_ASAP7_75t_SL g421 ( .A(n_409), .B(n_11), .Y(n_421) );
A2O1A1Ixp33_ASAP7_75t_L g422 ( .A1(n_394), .A2(n_258), .B(n_231), .C(n_299), .Y(n_422) );
A2O1A1Ixp33_ASAP7_75t_L g423 ( .A1(n_394), .A2(n_269), .B(n_235), .C(n_296), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_413), .Y(n_424) );
AOI22x1_ASAP7_75t_SL g425 ( .A1(n_410), .A2(n_272), .B1(n_237), .B2(n_238), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_393), .Y(n_426) );
AO21x2_ASAP7_75t_L g427 ( .A1(n_415), .A2(n_328), .B(n_313), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_398), .A2(n_270), .B1(n_295), .B2(n_294), .Y(n_428) );
OAI221xp5_ASAP7_75t_L g429 ( .A1(n_396), .A2(n_259), .B1(n_293), .B2(n_291), .C(n_282), .Y(n_429) );
AND2x2_ASAP7_75t_SL g430 ( .A(n_399), .B(n_12), .Y(n_430) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_412), .Y(n_431) );
AOI21xp5_ASAP7_75t_L g432 ( .A1(n_396), .A2(n_241), .B(n_234), .Y(n_432) );
INVx3_ASAP7_75t_L g433 ( .A(n_395), .Y(n_433) );
AO31x2_ASAP7_75t_L g434 ( .A1(n_390), .A2(n_13), .A3(n_15), .B(n_16), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_407), .Y(n_435) );
NAND2x1p5_ASAP7_75t_L g436 ( .A(n_400), .B(n_15), .Y(n_436) );
BUFx2_ASAP7_75t_L g437 ( .A(n_404), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_399), .Y(n_438) );
OAI21x1_ASAP7_75t_L g439 ( .A1(n_406), .A2(n_113), .B(n_183), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_407), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g441 ( .A1(n_404), .A2(n_280), .B1(n_276), .B2(n_274), .Y(n_441) );
OAI21xp5_ASAP7_75t_L g442 ( .A1(n_402), .A2(n_264), .B(n_257), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_408), .B(n_17), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_403), .B(n_244), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_414), .Y(n_445) );
INVx6_ASAP7_75t_L g446 ( .A(n_405), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_414), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_397), .Y(n_448) );
OAI21xp5_ASAP7_75t_L g449 ( .A1(n_392), .A2(n_252), .B(n_249), .Y(n_449) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_395), .Y(n_450) );
OAI21x1_ASAP7_75t_L g451 ( .A1(n_415), .A2(n_104), .B(n_21), .Y(n_451) );
O2A1O1Ixp33_ASAP7_75t_SL g452 ( .A1(n_392), .A2(n_103), .B(n_22), .C(n_23), .Y(n_452) );
OAI21x1_ASAP7_75t_L g453 ( .A1(n_415), .A2(n_112), .B(n_28), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_411), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_419), .Y(n_455) );
OA21x2_ASAP7_75t_L g456 ( .A1(n_440), .A2(n_114), .B(n_30), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_424), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_445), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g459 ( .A(n_448), .Y(n_459) );
BUFx3_ASAP7_75t_L g460 ( .A(n_417), .Y(n_460) );
BUFx4f_ASAP7_75t_SL g461 ( .A(n_431), .Y(n_461) );
BUFx3_ASAP7_75t_L g462 ( .A(n_450), .Y(n_462) );
NAND2x1p5_ASAP7_75t_L g463 ( .A(n_430), .B(n_17), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_447), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_438), .Y(n_465) );
BUFx3_ASAP7_75t_L g466 ( .A(n_450), .Y(n_466) );
INVx3_ASAP7_75t_L g467 ( .A(n_450), .Y(n_467) );
OAI22xp33_ASAP7_75t_L g468 ( .A1(n_437), .A2(n_37), .B1(n_41), .B2(n_44), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_427), .Y(n_469) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_426), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_433), .Y(n_471) );
AO31x2_ASAP7_75t_L g472 ( .A1(n_422), .A2(n_423), .A3(n_452), .B(n_416), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_434), .Y(n_473) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_443), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_434), .Y(n_475) );
INVx2_ASAP7_75t_SL g476 ( .A(n_446), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_436), .Y(n_477) );
INVx3_ASAP7_75t_L g478 ( .A(n_446), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_418), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_449), .B(n_47), .Y(n_480) );
BUFx6f_ASAP7_75t_L g481 ( .A(n_451), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_425), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_439), .Y(n_483) );
BUFx3_ASAP7_75t_L g484 ( .A(n_453), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_421), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_420), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_442), .Y(n_487) );
BUFx2_ASAP7_75t_L g488 ( .A(n_441), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_429), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_444), .Y(n_490) );
OAI21x1_ASAP7_75t_L g491 ( .A1(n_432), .A2(n_49), .B(n_50), .Y(n_491) );
AO31x2_ASAP7_75t_L g492 ( .A1(n_428), .A2(n_52), .A3(n_54), .B(n_55), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_419), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_454), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_454), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_419), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_454), .B(n_182), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_454), .Y(n_498) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_440), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_419), .Y(n_500) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_440), .Y(n_501) );
BUFx3_ASAP7_75t_L g502 ( .A(n_417), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_435), .Y(n_503) );
INVx6_ASAP7_75t_L g504 ( .A(n_450), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_454), .B(n_181), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_419), .Y(n_506) );
AND2x6_ASAP7_75t_L g507 ( .A(n_438), .B(n_63), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_435), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_419), .Y(n_509) );
INVx8_ASAP7_75t_L g510 ( .A(n_507), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_455), .Y(n_511) );
BUFx2_ASAP7_75t_L g512 ( .A(n_460), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_490), .B(n_64), .Y(n_513) );
NOR2x1_ASAP7_75t_L g514 ( .A(n_502), .B(n_66), .Y(n_514) );
INVxp67_ASAP7_75t_L g515 ( .A(n_499), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_470), .B(n_67), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_474), .B(n_68), .Y(n_517) );
BUFx2_ASAP7_75t_L g518 ( .A(n_461), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_464), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_493), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_463), .A2(n_69), .B1(n_77), .B2(n_79), .Y(n_521) );
NOR2x1p5_ASAP7_75t_L g522 ( .A(n_485), .B(n_80), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_465), .B(n_84), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_465), .B(n_85), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_457), .B(n_87), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_496), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_458), .B(n_180), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_500), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_506), .B(n_92), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_503), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_509), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_494), .B(n_94), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_495), .B(n_96), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_498), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_501), .Y(n_535) );
AND2x4_ASAP7_75t_L g536 ( .A(n_462), .B(n_97), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_478), .B(n_98), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_476), .B(n_101), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_488), .B(n_106), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_487), .B(n_115), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_471), .Y(n_541) );
INVx2_ASAP7_75t_SL g542 ( .A(n_459), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_482), .B(n_120), .Y(n_543) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_508), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_461), .B(n_122), .Y(n_545) );
AND2x4_ASAP7_75t_L g546 ( .A(n_466), .B(n_125), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_497), .Y(n_547) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_475), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_477), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_505), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_479), .Y(n_551) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_473), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_489), .B(n_134), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_469), .Y(n_554) );
BUFx3_ASAP7_75t_L g555 ( .A(n_504), .Y(n_555) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_467), .Y(n_556) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_544), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_511), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_512), .B(n_504), .Y(n_559) );
INVx3_ASAP7_75t_L g560 ( .A(n_510), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_519), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_520), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_549), .B(n_483), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_522), .A2(n_510), .B1(n_518), .B2(n_486), .Y(n_564) );
AND2x4_ASAP7_75t_L g565 ( .A(n_515), .B(n_484), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_534), .B(n_492), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_526), .Y(n_567) );
AND2x4_ASAP7_75t_L g568 ( .A(n_535), .B(n_507), .Y(n_568) );
AOI21xp33_ASAP7_75t_L g569 ( .A1(n_539), .A2(n_468), .B(n_480), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_528), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_531), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_541), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_547), .B(n_492), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_550), .B(n_492), .Y(n_574) );
NAND2xp33_ASAP7_75t_L g575 ( .A(n_510), .B(n_507), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_551), .B(n_472), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_517), .B(n_456), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g578 ( .A(n_542), .Y(n_578) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_554), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_530), .B(n_468), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_516), .B(n_481), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_548), .B(n_481), .Y(n_582) );
INVxp67_ASAP7_75t_L g583 ( .A(n_556), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_557), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_558), .Y(n_585) );
BUFx2_ASAP7_75t_L g586 ( .A(n_560), .Y(n_586) );
INVx2_ASAP7_75t_SL g587 ( .A(n_578), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_561), .Y(n_588) );
AND2x2_ASAP7_75t_SL g589 ( .A(n_575), .B(n_545), .Y(n_589) );
BUFx2_ASAP7_75t_L g590 ( .A(n_560), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_562), .B(n_552), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_559), .B(n_543), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_567), .Y(n_593) );
INVxp67_ASAP7_75t_SL g594 ( .A(n_579), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_570), .B(n_552), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_571), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_572), .B(n_523), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_581), .B(n_555), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_563), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_574), .B(n_524), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_583), .B(n_523), .Y(n_601) );
AND2x4_ASAP7_75t_L g602 ( .A(n_568), .B(n_514), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_585), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_599), .B(n_576), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_584), .B(n_583), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_587), .B(n_592), .Y(n_606) );
NAND2x1p5_ASAP7_75t_L g607 ( .A(n_589), .B(n_536), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_598), .B(n_565), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_588), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_594), .B(n_566), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_593), .Y(n_611) );
BUFx2_ASAP7_75t_L g612 ( .A(n_586), .Y(n_612) );
NAND2x1p5_ASAP7_75t_L g613 ( .A(n_590), .B(n_536), .Y(n_613) );
INVx1_ASAP7_75t_SL g614 ( .A(n_612), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_603), .Y(n_615) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_605), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_607), .A2(n_564), .B1(n_602), .B2(n_597), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_608), .B(n_596), .Y(n_618) );
AOI222xp33_ASAP7_75t_L g619 ( .A1(n_614), .A2(n_606), .B1(n_604), .B2(n_610), .C1(n_611), .C2(n_609), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_616), .B(n_610), .Y(n_620) );
AOI21xp33_ASAP7_75t_L g621 ( .A1(n_617), .A2(n_597), .B(n_601), .Y(n_621) );
OAI221xp5_ASAP7_75t_L g622 ( .A1(n_621), .A2(n_607), .B1(n_615), .B2(n_613), .C(n_521), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_619), .A2(n_618), .B1(n_613), .B2(n_600), .Y(n_623) );
NAND4xp75_ASAP7_75t_L g624 ( .A(n_623), .B(n_620), .C(n_513), .D(n_569), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_622), .B(n_595), .Y(n_625) );
NOR2x1_ASAP7_75t_L g626 ( .A(n_624), .B(n_546), .Y(n_626) );
NOR2x1_ASAP7_75t_L g627 ( .A(n_625), .B(n_538), .Y(n_627) );
NOR3xp33_ASAP7_75t_L g628 ( .A(n_626), .B(n_537), .C(n_553), .Y(n_628) );
AND2x4_ASAP7_75t_L g629 ( .A(n_627), .B(n_591), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_629), .Y(n_630) );
OAI21xp33_ASAP7_75t_SL g631 ( .A1(n_630), .A2(n_628), .B(n_591), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_631), .Y(n_632) );
OAI22x1_ASAP7_75t_L g633 ( .A1(n_632), .A2(n_525), .B1(n_540), .B2(n_529), .Y(n_633) );
AOI21xp33_ASAP7_75t_SL g634 ( .A1(n_633), .A2(n_138), .B(n_140), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_634), .A2(n_491), .B(n_533), .Y(n_635) );
OAI22xp33_ASAP7_75t_L g636 ( .A1(n_635), .A2(n_527), .B1(n_580), .B2(n_582), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_636), .B(n_532), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_637), .A2(n_573), .B1(n_577), .B2(n_582), .Y(n_638) );
endmodule