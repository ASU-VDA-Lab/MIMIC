module real_jpeg_14555_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx10_ASAP7_75t_L g124 ( 
.A(n_0),
.Y(n_124)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_3),
.A2(n_66),
.B1(n_67),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_3),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_3),
.A2(n_35),
.B1(n_37),
.B2(n_71),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_71),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_71),
.Y(n_276)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_6),
.A2(n_46),
.B1(n_47),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_6),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_6),
.A2(n_58),
.B1(n_66),
.B2(n_67),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_58),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_6),
.A2(n_35),
.B1(n_37),
.B2(n_58),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_8),
.A2(n_46),
.B1(n_47),
.B2(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_8),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_8),
.A2(n_66),
.B1(n_67),
.B2(n_108),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_108),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_8),
.A2(n_35),
.B1(n_37),
.B2(n_108),
.Y(n_203)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_10),
.A2(n_66),
.B1(n_67),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_10),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_104),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_104),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_10),
.A2(n_35),
.B1(n_37),
.B2(n_104),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_11),
.A2(n_66),
.B1(n_67),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_11),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_73),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_11),
.A2(n_35),
.B1(n_37),
.B2(n_73),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_73),
.Y(n_247)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_13),
.A2(n_66),
.B1(n_67),
.B2(n_101),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_13),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_13),
.A2(n_63),
.B(n_66),
.C(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_13),
.B(n_88),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_13),
.B(n_46),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_SL g188 ( 
.A1(n_13),
.A2(n_46),
.B(n_173),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_13),
.B(n_31),
.C(n_37),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_101),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_13),
.A2(n_122),
.B1(n_123),
.B2(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_13),
.B(n_49),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_110),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_14),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_110),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_14),
.A2(n_35),
.B1(n_37),
.B2(n_110),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_14),
.A2(n_66),
.B1(n_67),
.B2(n_110),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_15),
.A2(n_40),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_15),
.A2(n_35),
.B1(n_37),
.B2(n_40),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_15),
.A2(n_40),
.B1(n_66),
.B2(n_67),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_92),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_90),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_84),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_19),
.B(n_84),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_74),
.C(n_78),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_20),
.A2(n_74),
.B1(n_309),
.B2(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_20),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_59),
.B2(n_60),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_41),
.B2(n_42),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_23),
.B(n_74),
.C(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_23),
.A2(n_24),
.B1(n_79),
.B2(n_80),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_24),
.B(n_41),
.C(n_59),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_34),
.B(n_38),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_25),
.A2(n_38),
.B(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_25),
.A2(n_166),
.B(n_168),
.Y(n_165)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_26),
.B(n_114),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_26),
.A2(n_115),
.B1(n_167),
.B2(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_26),
.A2(n_115),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_26),
.A2(n_115),
.B1(n_190),
.B2(n_200),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_26),
.A2(n_115),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_26),
.A2(n_247),
.B(n_269),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_34),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_28),
.A2(n_29),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

NAND3xp33_ASAP7_75t_SL g174 ( 
.A(n_28),
.B(n_47),
.C(n_51),
.Y(n_174)
);

INVx5_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_29),
.A2(n_52),
.B(n_172),
.C(n_174),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_29),
.B(n_197),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_32),
.B1(n_35),
.B2(n_37),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_34),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_34),
.A2(n_149),
.B(n_150),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_34),
.B(n_101),
.Y(n_214)
);

INVx5_ASAP7_75t_SL g37 ( 
.A(n_35),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_35),
.B(n_209),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_37),
.B(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_39),
.B(n_115),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_53),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_43),
.A2(n_55),
.B(n_109),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_49),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_44),
.A2(n_49),
.B(n_54),
.Y(n_85)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_45),
.A2(n_55),
.B(n_83),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_47),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_46),
.A2(n_64),
.B(n_101),
.Y(n_129)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_49),
.B(n_57),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_49),
.A2(n_54),
.B1(n_82),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_50),
.A2(n_55),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_50),
.A2(n_55),
.B1(n_107),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_50),
.A2(n_55),
.B1(n_138),
.B2(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_50),
.A2(n_53),
.B(n_276),
.Y(n_275)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_81),
.B(n_83),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_70),
.B2(n_72),
.Y(n_60)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_61),
.A2(n_72),
.B(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_61),
.A2(n_62),
.B1(n_103),
.B2(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_61),
.A2(n_62),
.B1(n_143),
.B2(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_61),
.A2(n_254),
.B(n_278),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_61),
.A2(n_87),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_70),
.B(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_63),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_74),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_74),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_76),
.A2(n_88),
.B1(n_100),
.B2(n_102),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_88),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_78),
.B(n_312),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx24_ASAP7_75t_SL g321 ( 
.A(n_84),
.Y(n_321)
);

FAx1_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_86),
.CI(n_89),
.CON(n_84),
.SN(n_84)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_88),
.B(n_279),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_303),
.B(n_317),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_284),
.B(n_302),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_259),
.B(n_283),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_156),
.B(n_237),
.C(n_258),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_139),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_97),
.B(n_139),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_117),
.C(n_130),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_98),
.B(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_105),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_99),
.B(n_111),
.C(n_116),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_101),
.B(n_123),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_111),
.B1(n_112),
.B2(n_116),
.Y(n_105)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_113),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_117),
.A2(n_118),
.B1(n_130),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_127),
.B2(n_128),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_127),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_121),
.A2(n_154),
.B(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_121),
.A2(n_124),
.B1(n_202),
.B2(n_204),
.Y(n_201)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_122),
.A2(n_152),
.B(n_153),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_122),
.A2(n_123),
.B1(n_203),
.B2(n_211),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_122),
.A2(n_205),
.B(n_221),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_122),
.A2(n_123),
.B(n_266),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_134),
.Y(n_154)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_124),
.A2(n_125),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_124),
.B(n_177),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_126),
.Y(n_152)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.C(n_137),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_132),
.B1(n_135),
.B2(n_136),
.Y(n_164)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_133),
.B(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_137),
.B(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_146),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_140),
.B(n_147),
.C(n_155),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_145),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_142),
.B(n_144),
.C(n_145),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_155),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_148),
.B(n_151),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_149),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_150),
.B(n_168),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_235),
.B(n_236),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_178),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_159),
.B(n_162),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.C(n_169),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_165),
.A2(n_169),
.B1(n_170),
.B2(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_171),
.A2(n_175),
.B1(n_176),
.B2(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_171),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_177),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_191),
.B(n_234),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_180),
.B(n_183),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.C(n_189),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_184),
.B(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_186),
.A2(n_187),
.B1(n_189),
.B2(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_228),
.B(n_233),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_217),
.B(n_227),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_206),
.B(n_216),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_201),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_201),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_198),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_212),
.B(n_215),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_213),
.B(n_214),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_219),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_223),
.C(n_226),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_221),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_225),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_232),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_232),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_257),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_257),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_241),
.C(n_249),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_249),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_245),
.B2(n_248),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_248),
.Y(n_272)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_245),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_252),
.C(n_256),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_255),
.B2(n_256),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_255),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_261),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_282),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_270),
.B1(n_280),
.B2(n_281),
.Y(n_262)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_263),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_263),
.B(n_281),
.C(n_282),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_267),
.B2(n_268),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_264),
.A2(n_265),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_267),
.Y(n_295)
);

AOI21xp33_ASAP7_75t_L g310 ( 
.A1(n_265),
.A2(n_295),
.B(n_297),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_270),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_275),
.C(n_277),
.Y(n_287)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_276),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_279),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_301),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_301),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_288),
.B2(n_300),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_289),
.C(n_294),
.Y(n_315)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_288),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_294),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_292),
.B(n_293),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_290),
.B(n_292),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_306),
.C(n_310),
.Y(n_305)
);

FAx1_ASAP7_75t_SL g316 ( 
.A(n_293),
.B(n_306),
.CI(n_310),
.CON(n_316),
.SN(n_316)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_314),
.Y(n_303)
);

AOI21xp33_ASAP7_75t_L g317 ( 
.A1(n_304),
.A2(n_318),
.B(n_319),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_311),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_311),
.Y(n_319)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_316),
.Y(n_318)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_316),
.Y(n_320)
);


endmodule