module fake_jpeg_4744_n_331 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx3_ASAP7_75t_SL g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_SL g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_37),
.B(n_35),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_33),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_48),
.Y(n_60)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_50),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_21),
.Y(n_74)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_52),
.A2(n_18),
.B1(n_17),
.B2(n_16),
.Y(n_73)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_53),
.B(n_54),
.Y(n_107)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_55),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_20),
.C(n_26),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_57),
.B(n_87),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_52),
.A2(n_35),
.B1(n_17),
.B2(n_16),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_58),
.A2(n_96),
.B1(n_99),
.B2(n_102),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_17),
.B1(n_16),
.B2(n_35),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_59),
.A2(n_78),
.B1(n_88),
.B2(n_101),
.Y(n_105)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_42),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g115 ( 
.A(n_61),
.Y(n_115)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_38),
.B(n_26),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_64),
.B(n_65),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_24),
.Y(n_65)
);

INVx5_ASAP7_75t_SL g67 ( 
.A(n_36),
.Y(n_67)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_36),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_68),
.Y(n_124)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_24),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_71),
.B(n_75),
.Y(n_120)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_73),
.A2(n_86),
.B1(n_89),
.B2(n_97),
.Y(n_125)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_25),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_34),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_76),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_25),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_81),
.Y(n_121)
);

AO22x1_ASAP7_75t_SL g78 ( 
.A1(n_43),
.A2(n_20),
.B1(n_32),
.B2(n_34),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_31),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_82),
.Y(n_103)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_44),
.B(n_31),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_46),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_44),
.B(n_20),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_91),
.A2(n_93),
.B(n_100),
.C(n_22),
.Y(n_129)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

AOI21xp33_ASAP7_75t_SL g93 ( 
.A1(n_47),
.A2(n_32),
.B(n_22),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_49),
.A2(n_30),
.B1(n_18),
.B2(n_33),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_36),
.B(n_30),
.Y(n_98)
);

AO21x1_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_14),
.B(n_22),
.Y(n_114)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_37),
.B(n_29),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g101 ( 
.A1(n_50),
.A2(n_32),
.B1(n_27),
.B2(n_23),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_93),
.A2(n_27),
.B1(n_23),
.B2(n_15),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_112),
.B1(n_113),
.B2(n_116),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_78),
.A2(n_27),
.B1(n_23),
.B2(n_15),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_78),
.A2(n_62),
.B1(n_73),
.B2(n_55),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_79),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_62),
.A2(n_27),
.B1(n_23),
.B2(n_15),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_68),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_91),
.A2(n_22),
.B1(n_15),
.B2(n_19),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_57),
.C(n_91),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_138),
.C(n_141),
.Y(n_178)
);

HAxp5_ASAP7_75t_SL g207 ( 
.A(n_135),
.B(n_13),
.CON(n_207),
.SN(n_207)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_60),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_147),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_66),
.C(n_90),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_123),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_140),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_123),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_61),
.C(n_56),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_145),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_89),
.Y(n_143)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_144),
.B(n_162),
.Y(n_206)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_86),
.Y(n_146)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_63),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_149),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_120),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_99),
.Y(n_150)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_105),
.A2(n_112),
.B1(n_116),
.B2(n_129),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_151),
.A2(n_153),
.B1(n_171),
.B2(n_1),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_117),
.A2(n_80),
.B1(n_82),
.B2(n_53),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_152),
.A2(n_108),
.B1(n_104),
.B2(n_126),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_105),
.A2(n_80),
.B1(n_101),
.B2(n_67),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_157),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_22),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_155),
.A2(n_158),
.B(n_160),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_109),
.B(n_97),
.Y(n_156)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_21),
.B(n_22),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_161),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_117),
.A2(n_21),
.B(n_84),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_14),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_110),
.B(n_94),
.Y(n_163)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_121),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_165),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_122),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_166),
.B(n_167),
.Y(n_193)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_111),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_110),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_168),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_0),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_118),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_114),
.B(n_94),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_132),
.C(n_114),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_108),
.A2(n_84),
.B1(n_70),
.B2(n_3),
.Y(n_171)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_187),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_176),
.A2(n_191),
.B1(n_207),
.B2(n_154),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_179),
.B(n_162),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_185),
.B(n_190),
.Y(n_236)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_147),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_149),
.B(n_118),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_166),
.A2(n_104),
.B1(n_128),
.B2(n_103),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_197),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_136),
.A2(n_128),
.B1(n_70),
.B2(n_127),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_194),
.A2(n_198),
.B1(n_203),
.B2(n_205),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_134),
.B(n_127),
.C(n_103),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_157),
.C(n_155),
.Y(n_221)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_208),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_167),
.B(n_13),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_201),
.B(n_202),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_168),
.B(n_13),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_136),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_203)
);

NAND2x1_ASAP7_75t_SL g204 ( 
.A(n_170),
.B(n_2),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_204),
.A2(n_5),
.B(n_6),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_151),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_153),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_138),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_12),
.Y(n_238)
);

BUFx5_ASAP7_75t_L g210 ( 
.A(n_161),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_210),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_213),
.B(n_229),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_198),
.A2(n_144),
.B1(n_141),
.B2(n_164),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_216),
.A2(n_219),
.B1(n_233),
.B2(n_214),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_183),
.B(n_165),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_222),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_208),
.A2(n_164),
.B1(n_158),
.B2(n_137),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_197),
.A2(n_205),
.B1(n_194),
.B2(n_203),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_178),
.B(n_144),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_221),
.C(n_224),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_189),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_231),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_180),
.B(n_206),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_178),
.B(n_162),
.C(n_155),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_226),
.C(n_228),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_148),
.C(n_140),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_145),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_172),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_230),
.Y(n_260)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_188),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_199),
.A2(n_159),
.B1(n_139),
.B2(n_161),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_234),
.A2(n_238),
.B(n_185),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_196),
.B(n_174),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_181),
.B(n_196),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_239),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_212),
.A2(n_200),
.B(n_232),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_241),
.B(n_242),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_234),
.A2(n_200),
.B(n_204),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_195),
.C(n_180),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_250),
.C(n_261),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_216),
.A2(n_214),
.B1(n_219),
.B2(n_226),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_246),
.A2(n_255),
.B1(n_236),
.B2(n_229),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_239),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_248),
.A2(n_249),
.B1(n_259),
.B2(n_222),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_187),
.C(n_179),
.Y(n_250)
);

NAND3xp33_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_204),
.C(n_181),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_253),
.B(n_5),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_254),
.A2(n_12),
.B1(n_6),
.B2(n_7),
.Y(n_278)
);

OA21x2_ASAP7_75t_L g255 ( 
.A1(n_211),
.A2(n_190),
.B(n_191),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_225),
.A2(n_186),
.B(n_192),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_223),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_233),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_221),
.B(n_193),
.C(n_186),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_236),
.B(n_184),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_184),
.C(n_182),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_264),
.A2(n_270),
.B1(n_271),
.B2(n_273),
.Y(n_286)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_251),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_268),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_244),
.Y(n_291)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_251),
.Y(n_268)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_269),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_249),
.A2(n_237),
.B1(n_231),
.B2(n_173),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_240),
.A2(n_173),
.B1(n_174),
.B2(n_230),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_258),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_246),
.A2(n_182),
.B1(n_175),
.B2(n_227),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_262),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_275),
.Y(n_294)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_262),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_215),
.C(n_6),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_280),
.C(n_250),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_278),
.A2(n_252),
.B1(n_263),
.B2(n_247),
.Y(n_287)
);

AOI321xp33_ASAP7_75t_L g284 ( 
.A1(n_279),
.A2(n_254),
.A3(n_253),
.B1(n_242),
.B2(n_248),
.C(n_247),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_243),
.B(n_215),
.C(n_8),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_281),
.B(n_241),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_270),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_295),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_284),
.A2(n_272),
.B(n_279),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_287),
.Y(n_297)
);

XNOR2x1_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_243),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_291),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_259),
.B1(n_244),
.B2(n_261),
.Y(n_289)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_289),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_290),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_258),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_266),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_266),
.C(n_277),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_296),
.A2(n_304),
.B(n_307),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_299),
.B(n_303),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_301),
.B(n_290),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_285),
.A2(n_260),
.B1(n_255),
.B2(n_273),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_302),
.A2(n_282),
.B1(n_287),
.B2(n_298),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_291),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_276),
.C(n_280),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_256),
.C(n_271),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_306),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_10),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_297),
.A2(n_284),
.B(n_294),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_310),
.A2(n_313),
.B1(n_315),
.B2(n_304),
.Y(n_317)
);

A2O1A1Ixp33_ASAP7_75t_SL g312 ( 
.A1(n_296),
.A2(n_286),
.B(n_255),
.C(n_288),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_312),
.A2(n_316),
.B1(n_7),
.B2(n_8),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_305),
.C(n_303),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_307),
.A2(n_255),
.B1(n_257),
.B2(n_260),
.Y(n_315)
);

NOR2x1_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_7),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_319),
.C(n_321),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_318),
.A2(n_320),
.B1(n_310),
.B2(n_312),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_316),
.A2(n_301),
.B1(n_305),
.B2(n_299),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_312),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_320),
.A2(n_322),
.B(n_311),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_324),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_308),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_325),
.B(n_321),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_326),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_327),
.Y(n_331)
);


endmodule