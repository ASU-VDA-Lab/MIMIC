module fake_ariane_523_n_1971 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1971);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1971;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_279;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_212;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_604;
wire n_439;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_1126;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g204 ( 
.A(n_16),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_189),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_150),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_5),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_81),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_135),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_188),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_121),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_57),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_162),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_43),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_198),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_61),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_167),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_23),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_125),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_13),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_144),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_45),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_86),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_40),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_115),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_66),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_156),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_53),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_36),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_14),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_54),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_186),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_6),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_99),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_53),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_49),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_129),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_159),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_185),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_69),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_119),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_120),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_76),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_90),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_60),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_106),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_39),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_175),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_158),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_25),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_173),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_127),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_107),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_164),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_199),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_36),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_134),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_181),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_20),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_97),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_203),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_113),
.Y(n_263)
);

INVxp67_ASAP7_75t_SL g264 ( 
.A(n_26),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_85),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_26),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_182),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_171),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_124),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_47),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_21),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_154),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_75),
.Y(n_273)
);

BUFx2_ASAP7_75t_SL g274 ( 
.A(n_38),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_118),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_84),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_7),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_201),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_196),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_83),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_21),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_123),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_22),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_143),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_184),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_92),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_35),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_139),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_131),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_146),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_122),
.Y(n_291)
);

BUFx10_ASAP7_75t_L g292 ( 
.A(n_191),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_0),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_157),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_57),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_147),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_95),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_47),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_73),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_93),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_91),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_151),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_48),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_78),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_73),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_22),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_174),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_179),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_195),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_192),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_9),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_7),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_10),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_137),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_34),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_165),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_110),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_11),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_200),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_160),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_42),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_172),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_41),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_103),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_148),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_41),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_112),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_9),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_65),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_46),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_128),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_169),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_96),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_35),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_11),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_60),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_6),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_34),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_59),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_10),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_62),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_177),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_142),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_77),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_161),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_5),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_155),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_72),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_50),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_138),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_15),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_23),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_136),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_194),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_117),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_89),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_78),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_82),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_202),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_37),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_44),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_16),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_80),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_52),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_132),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_74),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_149),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_178),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_87),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_28),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_176),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_27),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_140),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_187),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_45),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_76),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_133),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_166),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_111),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_37),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_105),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_3),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_75),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_193),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_170),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_31),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_88),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_19),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_168),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_30),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_43),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_94),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_70),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_29),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_141),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_19),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_20),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_15),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_77),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_126),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_40),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_153),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_42),
.Y(n_403)
);

BUFx10_ASAP7_75t_L g404 ( 
.A(n_33),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_2),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_1),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_183),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_68),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_102),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_237),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_289),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_237),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_221),
.B(n_0),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_289),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_210),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_252),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_259),
.Y(n_417)
);

NOR2xp67_ASAP7_75t_L g418 ( 
.A(n_237),
.B(n_1),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_344),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_393),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_393),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_276),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_221),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_223),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_205),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_223),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_406),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_309),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_406),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_205),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_355),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_292),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_328),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_209),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g435 ( 
.A(n_344),
.Y(n_435)
);

INVxp67_ASAP7_75t_SL g436 ( 
.A(n_344),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_209),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_214),
.B(n_2),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_381),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_292),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_204),
.Y(n_441)
);

INVxp33_ASAP7_75t_SL g442 ( 
.A(n_337),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_407),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_292),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_204),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_213),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_239),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_251),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_213),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_292),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_266),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_328),
.Y(n_452)
);

INVxp33_ASAP7_75t_SL g453 ( 
.A(n_242),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_274),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_217),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_217),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_273),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_383),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_231),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_231),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_234),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_312),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_234),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_344),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_383),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_246),
.Y(n_466)
);

NOR2xp67_ASAP7_75t_L g467 ( 
.A(n_366),
.B(n_3),
.Y(n_467)
);

BUFx6f_ASAP7_75t_SL g468 ( 
.A(n_207),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_388),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_246),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_270),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_388),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_215),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_219),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_270),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_277),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_326),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_225),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_277),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_382),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_281),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_281),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_274),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_207),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_293),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_224),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_224),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_293),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_227),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_305),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_404),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_305),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_229),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_404),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_306),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_306),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_214),
.B(n_4),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_315),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_230),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_315),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_232),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_330),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_236),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_216),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_330),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_216),
.B(n_4),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_404),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_338),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_404),
.Y(n_509)
);

INVx1_ASAP7_75t_SL g510 ( 
.A(n_208),
.Y(n_510)
);

INVxp67_ASAP7_75t_SL g511 ( 
.A(n_344),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_338),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_241),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_341),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_341),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_244),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_346),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_248),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_257),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_260),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_346),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_348),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_271),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_419),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_435),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_464),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_419),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_419),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_436),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_434),
.B(n_299),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_464),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_511),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_447),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_447),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_447),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_510),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_434),
.B(n_299),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_437),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_410),
.B(n_412),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_453),
.B(n_454),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_433),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_465),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_447),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_513),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_465),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_504),
.B(n_329),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_504),
.B(n_368),
.Y(n_547)
);

BUFx8_ASAP7_75t_L g548 ( 
.A(n_468),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_418),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_441),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_445),
.Y(n_551)
);

INVx4_ASAP7_75t_L g552 ( 
.A(n_447),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_446),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_449),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_455),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_456),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_459),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_413),
.B(n_460),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_461),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_420),
.B(n_218),
.Y(n_560)
);

OA21x2_ASAP7_75t_L g561 ( 
.A1(n_438),
.A2(n_226),
.B(n_218),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_463),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_421),
.B(n_466),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_470),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_471),
.Y(n_565)
);

NAND2xp33_ASAP7_75t_L g566 ( 
.A(n_413),
.B(n_344),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_518),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_475),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_476),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_479),
.B(n_329),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_481),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_482),
.B(n_334),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_485),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_488),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_490),
.B(n_334),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_492),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_495),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_496),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_498),
.B(n_226),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_502),
.B(n_348),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_505),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_508),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_512),
.B(n_228),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_514),
.Y(n_584)
);

OA21x2_ASAP7_75t_L g585 ( 
.A1(n_497),
.A2(n_243),
.B(n_228),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_515),
.Y(n_586)
);

INVx4_ASAP7_75t_L g587 ( 
.A(n_468),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_517),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_415),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_521),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_452),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_522),
.Y(n_592)
);

NAND2xp33_ASAP7_75t_L g593 ( 
.A(n_425),
.B(n_253),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_506),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_500),
.Y(n_595)
);

AND2x6_ASAP7_75t_L g596 ( 
.A(n_423),
.B(n_253),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_467),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_483),
.B(n_243),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_453),
.B(n_249),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_468),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_424),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_432),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_426),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_432),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_452),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_427),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_440),
.B(n_249),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_429),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_519),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_440),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_444),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_484),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_525),
.B(n_444),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_611),
.B(n_411),
.Y(n_614)
);

INVx4_ASAP7_75t_SL g615 ( 
.A(n_596),
.Y(n_615)
);

BUFx10_ASAP7_75t_L g616 ( 
.A(n_540),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_525),
.B(n_450),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_524),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_611),
.B(n_607),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_524),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_524),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_607),
.B(n_411),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_540),
.B(n_414),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_595),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_538),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_538),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_529),
.B(n_450),
.Y(n_627)
);

AND2x6_ASAP7_75t_L g628 ( 
.A(n_602),
.B(n_250),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_548),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_524),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_596),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_563),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_536),
.B(n_458),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_602),
.B(n_414),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_524),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_529),
.B(n_532),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_563),
.Y(n_637)
);

INVx4_ASAP7_75t_SL g638 ( 
.A(n_596),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_552),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_599),
.A2(n_430),
.B1(n_442),
.B2(n_458),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_563),
.Y(n_641)
);

BUFx8_ASAP7_75t_SL g642 ( 
.A(n_567),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_550),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_532),
.B(n_520),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_594),
.B(n_473),
.Y(n_645)
);

AND3x2_ASAP7_75t_L g646 ( 
.A(n_536),
.B(n_264),
.C(n_351),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_527),
.Y(n_647)
);

INVx8_ASAP7_75t_L g648 ( 
.A(n_596),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_527),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_550),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_527),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_554),
.Y(n_652)
);

INVx4_ASAP7_75t_SL g653 ( 
.A(n_596),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_527),
.Y(n_654)
);

AND2x6_ASAP7_75t_L g655 ( 
.A(n_602),
.B(n_604),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_602),
.B(n_250),
.Y(n_656)
);

OR2x6_ASAP7_75t_L g657 ( 
.A(n_558),
.B(n_351),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_596),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_561),
.A2(n_487),
.B1(n_486),
.B2(n_472),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_527),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_548),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_599),
.B(n_473),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_602),
.B(n_256),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_594),
.B(n_474),
.Y(n_664)
);

NAND2x1p5_ASAP7_75t_L g665 ( 
.A(n_587),
.B(n_265),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_594),
.B(n_474),
.Y(n_666)
);

OAI22xp33_ASAP7_75t_SL g667 ( 
.A1(n_598),
.A2(n_472),
.B1(n_469),
.B2(n_478),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_528),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_552),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_528),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_528),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_548),
.Y(n_672)
);

INVx4_ASAP7_75t_L g673 ( 
.A(n_596),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_528),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_594),
.B(n_478),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_548),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_528),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_548),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_602),
.B(n_256),
.Y(n_679)
);

OAI22x1_ASAP7_75t_L g680 ( 
.A1(n_567),
.A2(n_469),
.B1(n_541),
.B2(n_542),
.Y(n_680)
);

INVx6_ASAP7_75t_L g681 ( 
.A(n_587),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_554),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_554),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_602),
.B(n_258),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_558),
.B(n_489),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_551),
.Y(n_686)
);

BUFx10_ASAP7_75t_L g687 ( 
.A(n_602),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_604),
.B(n_258),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_593),
.B(n_489),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_594),
.B(n_493),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_593),
.B(n_493),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_526),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_604),
.B(n_263),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_554),
.Y(n_694)
);

CKINVDCx16_ASAP7_75t_R g695 ( 
.A(n_544),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_554),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_553),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_526),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_558),
.B(n_530),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_554),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_594),
.B(n_499),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_564),
.Y(n_702)
);

BUFx10_ASAP7_75t_L g703 ( 
.A(n_604),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_564),
.Y(n_704)
);

AND2x6_ASAP7_75t_L g705 ( 
.A(n_604),
.B(n_263),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_594),
.B(n_499),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_555),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_526),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_531),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_600),
.B(n_501),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_600),
.B(n_501),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_558),
.B(n_352),
.Y(n_712)
);

NAND3xp33_ASAP7_75t_L g713 ( 
.A(n_595),
.B(n_516),
.C(n_503),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_568),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_552),
.Y(n_715)
);

AND2x2_ASAP7_75t_SL g716 ( 
.A(n_566),
.B(n_604),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_552),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_568),
.Y(n_718)
);

OAI21xp33_ASAP7_75t_SL g719 ( 
.A1(n_598),
.A2(n_360),
.B(n_352),
.Y(n_719)
);

INVx2_ASAP7_75t_SL g720 ( 
.A(n_542),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_555),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_545),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_531),
.Y(n_723)
);

BUFx6f_ASAP7_75t_SL g724 ( 
.A(n_604),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_552),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_571),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_604),
.B(n_267),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_610),
.B(n_267),
.Y(n_728)
);

BUFx2_ASAP7_75t_L g729 ( 
.A(n_545),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_541),
.B(n_503),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_531),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_610),
.B(n_286),
.Y(n_732)
);

INVx4_ASAP7_75t_L g733 ( 
.A(n_596),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_554),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_L g735 ( 
.A(n_610),
.B(n_239),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_571),
.Y(n_736)
);

NOR2x1p5_ASAP7_75t_L g737 ( 
.A(n_609),
.B(n_516),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_558),
.B(n_360),
.Y(n_738)
);

INVx4_ASAP7_75t_L g739 ( 
.A(n_596),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_573),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_559),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_559),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_559),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_610),
.B(n_286),
.Y(n_744)
);

BUFx4f_ASAP7_75t_L g745 ( 
.A(n_596),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_559),
.Y(n_746)
);

AND3x2_ASAP7_75t_L g747 ( 
.A(n_591),
.B(n_605),
.C(n_567),
.Y(n_747)
);

OR2x6_ASAP7_75t_L g748 ( 
.A(n_603),
.B(n_362),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_561),
.A2(n_362),
.B1(n_372),
.B2(n_370),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_574),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_574),
.Y(n_751)
);

AND3x2_ASAP7_75t_L g752 ( 
.A(n_591),
.B(n_372),
.C(n_370),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_582),
.Y(n_753)
);

INVx5_ASAP7_75t_L g754 ( 
.A(n_543),
.Y(n_754)
);

AND2x6_ASAP7_75t_L g755 ( 
.A(n_610),
.B(n_294),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_610),
.B(n_549),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_555),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_530),
.B(n_390),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_559),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_610),
.B(n_559),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_584),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_745),
.B(n_610),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_695),
.Y(n_763)
);

HB1xp67_ASAP7_75t_L g764 ( 
.A(n_729),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_619),
.B(n_609),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_699),
.B(n_603),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_662),
.B(n_549),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_625),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_745),
.B(n_605),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_642),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_745),
.B(n_559),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_689),
.A2(n_566),
.B1(n_547),
.B2(n_561),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_644),
.B(n_555),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_624),
.B(n_555),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_624),
.B(n_556),
.Y(n_775)
);

INVxp67_ASAP7_75t_L g776 ( 
.A(n_633),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_622),
.B(n_601),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_626),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_691),
.B(n_556),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_616),
.B(n_645),
.Y(n_780)
);

NOR3xp33_ASAP7_75t_L g781 ( 
.A(n_730),
.B(n_606),
.C(n_601),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_633),
.B(n_720),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_692),
.Y(n_783)
);

AND2x2_ASAP7_75t_SL g784 ( 
.A(n_716),
.B(n_561),
.Y(n_784)
);

NAND2x1p5_ASAP7_75t_L g785 ( 
.A(n_629),
.B(n_661),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_623),
.B(n_664),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_666),
.B(n_556),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_685),
.A2(n_547),
.B1(n_585),
.B2(n_523),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_722),
.B(n_685),
.Y(n_789)
);

NOR2x1p5_ASAP7_75t_L g790 ( 
.A(n_713),
.B(n_589),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_643),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_699),
.B(n_603),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_675),
.B(n_556),
.Y(n_793)
);

OAI21xp33_ASAP7_75t_L g794 ( 
.A1(n_614),
.A2(n_597),
.B(n_608),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_690),
.B(n_556),
.Y(n_795)
);

OR2x2_ASAP7_75t_L g796 ( 
.A(n_722),
.B(n_589),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_640),
.B(n_612),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_707),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_698),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_650),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_701),
.B(n_584),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_706),
.B(n_586),
.Y(n_802)
);

INVxp33_ASAP7_75t_L g803 ( 
.A(n_642),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_631),
.B(n_559),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_616),
.B(n_608),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_631),
.B(n_577),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_708),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_758),
.B(n_612),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_631),
.B(n_577),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_721),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_613),
.B(n_586),
.Y(n_811)
);

BUFx6f_ASAP7_75t_SL g812 ( 
.A(n_629),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_636),
.B(n_617),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_627),
.B(n_588),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_686),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_710),
.B(n_588),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_708),
.Y(n_817)
);

OR2x2_ASAP7_75t_L g818 ( 
.A(n_680),
.B(n_590),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_697),
.B(n_590),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_658),
.B(n_577),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_658),
.B(n_577),
.Y(n_821)
);

NOR3xp33_ASAP7_75t_L g822 ( 
.A(n_667),
.B(n_539),
.C(n_390),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_709),
.Y(n_823)
);

NAND2xp33_ASAP7_75t_L g824 ( 
.A(n_655),
.B(n_577),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_702),
.B(n_530),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_704),
.B(n_546),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_711),
.B(n_557),
.Y(n_827)
);

NOR3xp33_ASAP7_75t_L g828 ( 
.A(n_719),
.B(n_637),
.C(n_632),
.Y(n_828)
);

OR2x2_ASAP7_75t_L g829 ( 
.A(n_680),
.B(n_579),
.Y(n_829)
);

NAND3xp33_ASAP7_75t_L g830 ( 
.A(n_756),
.B(n_557),
.C(n_585),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_758),
.B(n_491),
.Y(n_831)
);

AOI221xp5_ASAP7_75t_L g832 ( 
.A1(n_641),
.A2(n_580),
.B1(n_579),
.B2(n_583),
.C(n_287),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_737),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_714),
.B(n_546),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_748),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_718),
.B(n_546),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_749),
.A2(n_585),
.B1(n_537),
.B2(n_565),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_659),
.B(n_494),
.Y(n_838)
);

OAI221xp5_ASAP7_75t_L g839 ( 
.A1(n_657),
.A2(n_583),
.B1(n_560),
.B2(n_539),
.C(n_295),
.Y(n_839)
);

AOI221xp5_ASAP7_75t_L g840 ( 
.A1(n_738),
.A2(n_580),
.B1(n_298),
.B2(n_283),
.C(n_303),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_657),
.A2(n_585),
.B1(n_537),
.B2(n_557),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_738),
.B(n_507),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_747),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_726),
.B(n_587),
.Y(n_844)
);

OR2x6_ASAP7_75t_L g845 ( 
.A(n_657),
.B(n_570),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_736),
.B(n_587),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_760),
.A2(n_560),
.B(n_562),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_657),
.B(n_509),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_SL g849 ( 
.A(n_661),
.B(n_416),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_723),
.Y(n_850)
);

BUFx3_ASAP7_75t_L g851 ( 
.A(n_672),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_634),
.A2(n_537),
.B1(n_557),
.B2(n_562),
.Y(n_852)
);

AO221x1_ASAP7_75t_L g853 ( 
.A1(n_639),
.A2(n_253),
.B1(n_367),
.B2(n_359),
.C(n_324),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_721),
.B(n_557),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_740),
.B(n_587),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_673),
.B(n_577),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_712),
.B(n_748),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_634),
.A2(n_537),
.B1(n_557),
.B2(n_562),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_757),
.B(n_577),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_673),
.B(n_581),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_731),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_750),
.B(n_537),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_751),
.B(n_581),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_753),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_761),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_733),
.B(n_581),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_618),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_757),
.B(n_581),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_733),
.B(n_565),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_618),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_748),
.B(n_565),
.Y(n_871)
);

HB1xp67_ASAP7_75t_L g872 ( 
.A(n_748),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_731),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_620),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_620),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_621),
.B(n_569),
.Y(n_876)
);

OR2x2_ASAP7_75t_L g877 ( 
.A(n_665),
.B(n_580),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_621),
.B(n_569),
.Y(n_878)
);

BUFx10_ASAP7_75t_L g879 ( 
.A(n_752),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_716),
.A2(n_576),
.B1(n_578),
.B2(n_569),
.Y(n_880)
);

CKINVDCx20_ASAP7_75t_R g881 ( 
.A(n_672),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_733),
.B(n_576),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_639),
.A2(n_311),
.B1(n_313),
.B2(n_304),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_SL g884 ( 
.A1(n_665),
.A2(n_451),
.B1(n_457),
.B2(n_448),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_739),
.B(n_576),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_676),
.B(n_417),
.Y(n_886)
);

OAI22xp33_ASAP7_75t_L g887 ( 
.A1(n_739),
.A2(n_592),
.B1(n_578),
.B2(n_321),
.Y(n_887)
);

OAI22xp33_ASAP7_75t_L g888 ( 
.A1(n_739),
.A2(n_592),
.B1(n_578),
.B2(n_323),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_630),
.B(n_592),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_639),
.B(n_570),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_676),
.B(n_678),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_630),
.B(n_570),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_635),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_635),
.B(n_572),
.Y(n_894)
);

NOR2x1p5_ASAP7_75t_L g895 ( 
.A(n_678),
.B(n_318),
.Y(n_895)
);

OAI22xp33_ASAP7_75t_SL g896 ( 
.A1(n_656),
.A2(n_339),
.B1(n_408),
.B2(n_405),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_647),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_687),
.B(n_294),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_649),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_649),
.B(n_651),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_669),
.B(n_572),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_651),
.Y(n_902)
);

NOR3xp33_ASAP7_75t_L g903 ( 
.A(n_656),
.B(n_336),
.C(n_335),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_669),
.B(n_575),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_687),
.B(n_296),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_654),
.B(n_575),
.Y(n_906)
);

BUFx12f_ASAP7_75t_SL g907 ( 
.A(n_652),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_654),
.Y(n_908)
);

AND2x6_ASAP7_75t_SL g909 ( 
.A(n_646),
.B(n_575),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_660),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_663),
.A2(n_373),
.B1(n_300),
.B2(n_307),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_669),
.B(n_715),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_660),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_779),
.A2(n_760),
.B(n_684),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_L g915 ( 
.A1(n_788),
.A2(n_428),
.B1(n_431),
.B2(n_422),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_L g916 ( 
.A1(n_765),
.A2(n_715),
.B1(n_725),
.B2(n_717),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_787),
.A2(n_684),
.B(n_679),
.Y(n_917)
);

OR2x2_ASAP7_75t_SL g918 ( 
.A(n_796),
.B(n_439),
.Y(n_918)
);

AO21x1_ASAP7_75t_L g919 ( 
.A1(n_786),
.A2(n_688),
.B(n_679),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_791),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_793),
.A2(n_795),
.B(n_813),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_891),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_764),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_765),
.A2(n_443),
.B1(n_693),
.B2(n_688),
.Y(n_924)
);

AOI22xp5_ASAP7_75t_L g925 ( 
.A1(n_777),
.A2(n_693),
.B1(n_728),
.B2(n_727),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_800),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_801),
.A2(n_728),
.B(n_727),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_777),
.A2(n_744),
.B1(n_732),
.B2(n_705),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_776),
.A2(n_670),
.B(n_671),
.C(n_668),
.Y(n_929)
);

AOI21x1_ASAP7_75t_L g930 ( 
.A1(n_771),
.A2(n_744),
.B(n_732),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_845),
.B(n_615),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_816),
.B(n_668),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_767),
.A2(n_671),
.B(n_674),
.C(n_670),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_816),
.B(n_674),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_912),
.A2(n_703),
.B(n_735),
.Y(n_935)
);

O2A1O1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_782),
.A2(n_677),
.B(n_717),
.C(n_715),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_912),
.A2(n_735),
.B(n_725),
.Y(n_937)
);

OAI321xp33_ASAP7_75t_L g938 ( 
.A1(n_839),
.A2(n_392),
.A3(n_300),
.B1(n_307),
.B2(n_316),
.C(n_319),
.Y(n_938)
);

INVx5_ASAP7_75t_L g939 ( 
.A(n_845),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_798),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_811),
.B(n_677),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_900),
.A2(n_725),
.B(n_717),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_802),
.A2(n_724),
.B(n_655),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_811),
.B(n_628),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_830),
.A2(n_759),
.B(n_742),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_805),
.B(n_628),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_845),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_805),
.B(n_462),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_847),
.A2(n_742),
.B(n_741),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_762),
.A2(n_724),
.B(n_655),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_798),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_780),
.B(n_628),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_780),
.B(n_628),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_831),
.B(n_477),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_814),
.B(n_628),
.Y(n_955)
);

OAI21xp5_ASAP7_75t_L g956 ( 
.A1(n_804),
.A2(n_809),
.B(n_806),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_762),
.A2(n_724),
.B(n_655),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_890),
.B(n_628),
.Y(n_958)
);

NAND3xp33_ASAP7_75t_L g959 ( 
.A(n_781),
.B(n_480),
.C(n_349),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_804),
.A2(n_655),
.B(n_648),
.Y(n_960)
);

AND2x2_ASAP7_75t_SL g961 ( 
.A(n_838),
.B(n_849),
.Y(n_961)
);

AOI22xp5_ASAP7_75t_L g962 ( 
.A1(n_789),
.A2(n_755),
.B1(n_705),
.B2(n_648),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_890),
.B(n_901),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_815),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_901),
.B(n_766),
.Y(n_965)
);

OAI21xp33_ASAP7_75t_L g966 ( 
.A1(n_832),
.A2(n_357),
.B(n_340),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_799),
.Y(n_967)
);

CKINVDCx8_ASAP7_75t_R g968 ( 
.A(n_770),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_766),
.B(n_705),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_792),
.B(n_705),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_773),
.B(n_648),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_894),
.A2(n_759),
.B(n_746),
.C(n_743),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_806),
.A2(n_655),
.B(n_648),
.Y(n_973)
);

NAND2x1p5_ASAP7_75t_L g974 ( 
.A(n_891),
.B(n_652),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_809),
.A2(n_743),
.B(n_741),
.Y(n_975)
);

AOI33xp33_ASAP7_75t_L g976 ( 
.A1(n_840),
.A2(n_575),
.A3(n_395),
.B1(n_392),
.B2(n_384),
.B3(n_400),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_820),
.A2(n_746),
.B(n_683),
.Y(n_977)
);

INVx4_ASAP7_75t_L g978 ( 
.A(n_851),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_886),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_792),
.B(n_705),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_842),
.B(n_652),
.Y(n_981)
);

AOI21x1_ASAP7_75t_L g982 ( 
.A1(n_771),
.A2(n_535),
.B(n_322),
.Y(n_982)
);

HB1xp67_ASAP7_75t_L g983 ( 
.A(n_877),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_821),
.A2(n_683),
.B(n_682),
.Y(n_984)
);

AOI21x1_ASAP7_75t_L g985 ( 
.A1(n_876),
.A2(n_535),
.B(n_322),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_857),
.B(n_615),
.Y(n_986)
);

AOI21x1_ASAP7_75t_L g987 ( 
.A1(n_878),
.A2(n_535),
.B(n_324),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_797),
.B(n_682),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_848),
.B(n_682),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_799),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_851),
.Y(n_991)
);

BUFx8_ASAP7_75t_L g992 ( 
.A(n_812),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_821),
.A2(n_683),
.B(n_682),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_SL g994 ( 
.A(n_763),
.B(n_755),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_772),
.A2(n_904),
.B1(n_775),
.B2(n_774),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_856),
.A2(n_696),
.B(n_694),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_SL g997 ( 
.A(n_884),
.B(n_755),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_860),
.A2(n_696),
.B(n_694),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_833),
.B(n_694),
.Y(n_999)
);

AOI21x1_ASAP7_75t_L g1000 ( 
.A1(n_889),
.A2(n_359),
.B(n_316),
.Y(n_1000)
);

AND2x4_ASAP7_75t_L g1001 ( 
.A(n_895),
.B(n_615),
.Y(n_1001)
);

AND2x6_ASAP7_75t_L g1002 ( 
.A(n_841),
.B(n_615),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_835),
.B(n_696),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_808),
.B(n_755),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_769),
.B(n_638),
.Y(n_1005)
);

CKINVDCx8_ASAP7_75t_R g1006 ( 
.A(n_909),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_904),
.B(n_575),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_794),
.A2(n_384),
.B(n_373),
.C(n_371),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_769),
.B(n_696),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_828),
.B(n_700),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_817),
.Y(n_1011)
);

BUFx2_ASAP7_75t_SL g1012 ( 
.A(n_812),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_864),
.B(n_700),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_810),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_829),
.B(n_700),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_872),
.B(n_734),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_865),
.B(n_734),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_768),
.B(n_778),
.Y(n_1018)
);

AO21x1_ASAP7_75t_L g1019 ( 
.A1(n_827),
.A2(n_367),
.B(n_238),
.Y(n_1019)
);

O2A1O1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_825),
.A2(n_235),
.B(n_238),
.C(n_268),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_906),
.Y(n_1021)
);

A2O1A1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_827),
.A2(n_358),
.B(n_354),
.C(n_290),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_892),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_866),
.A2(n_754),
.B(n_534),
.Y(n_1024)
);

INVxp67_ASAP7_75t_SL g1025 ( 
.A(n_810),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_826),
.B(n_638),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_896),
.B(n_638),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_866),
.A2(n_754),
.B(n_534),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_L g1029 ( 
.A1(n_784),
.A2(n_653),
.B1(n_386),
.B2(n_399),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_824),
.A2(n_754),
.B(n_534),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_859),
.A2(n_534),
.B(n_533),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_818),
.B(n_361),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_834),
.B(n_653),
.Y(n_1033)
);

AOI21x1_ASAP7_75t_L g1034 ( 
.A1(n_863),
.A2(n_681),
.B(n_653),
.Y(n_1034)
);

OAI21xp33_ASAP7_75t_L g1035 ( 
.A1(n_883),
.A2(n_375),
.B(n_364),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_859),
.A2(n_533),
.B(n_543),
.Y(n_1036)
);

NAND2xp33_ASAP7_75t_L g1037 ( 
.A(n_844),
.B(n_376),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_887),
.B(n_888),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_868),
.A2(n_533),
.B(n_543),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_836),
.B(n_653),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_819),
.B(n_681),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_867),
.A2(n_391),
.B(n_396),
.C(n_397),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_870),
.A2(n_403),
.B(n_401),
.C(n_394),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_874),
.A2(n_902),
.B(n_893),
.C(n_875),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_785),
.Y(n_1045)
);

NOR2x1_ASAP7_75t_L g1046 ( 
.A(n_790),
.B(n_288),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_868),
.A2(n_533),
.B(n_543),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_862),
.B(n_681),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_871),
.B(n_380),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_854),
.A2(n_533),
.B(n_543),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_908),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_869),
.A2(n_379),
.B(n_398),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_843),
.B(n_8),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_903),
.B(n_206),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_869),
.A2(n_310),
.B(n_409),
.Y(n_1055)
);

AOI21xp33_ASAP7_75t_L g1056 ( 
.A1(n_913),
.A2(n_363),
.B(n_302),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_882),
.A2(n_308),
.B(n_402),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_897),
.A2(n_910),
.B(n_899),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_897),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_881),
.B(n_211),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_784),
.A2(n_314),
.B1(n_389),
.B2(n_387),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_822),
.B(n_212),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_899),
.A2(n_543),
.B(n_385),
.Y(n_1063)
);

INVx4_ASAP7_75t_L g1064 ( 
.A(n_785),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_837),
.B(n_220),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_846),
.A2(n_301),
.B1(n_378),
.B2(n_233),
.Y(n_1066)
);

BUFx2_ASAP7_75t_L g1067 ( 
.A(n_907),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_837),
.B(n_222),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_855),
.A2(n_317),
.B1(n_240),
.B2(n_374),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_882),
.B(n_12),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_911),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_910),
.A2(n_543),
.B(n_297),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_885),
.A2(n_291),
.B(n_369),
.Y(n_1073)
);

INVx4_ASAP7_75t_L g1074 ( 
.A(n_879),
.Y(n_1074)
);

AO21x1_ASAP7_75t_L g1075 ( 
.A1(n_898),
.A2(n_377),
.B(n_239),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_885),
.A2(n_285),
.B(n_365),
.Y(n_1076)
);

NAND2x1p5_ASAP7_75t_L g1077 ( 
.A(n_905),
.B(n_239),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_905),
.A2(n_284),
.B(n_356),
.Y(n_1078)
);

AO32x1_ASAP7_75t_L g1079 ( 
.A1(n_995),
.A2(n_853),
.A3(n_850),
.B1(n_861),
.B2(n_873),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_925),
.A2(n_963),
.B(n_938),
.C(n_1052),
.Y(n_1080)
);

CKINVDCx8_ASAP7_75t_R g1081 ( 
.A(n_1012),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_948),
.B(n_803),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_965),
.A2(n_880),
.B1(n_858),
.B2(n_852),
.Y(n_1083)
);

INVxp67_ASAP7_75t_L g1084 ( 
.A(n_923),
.Y(n_1084)
);

AO21x1_ASAP7_75t_L g1085 ( 
.A1(n_1038),
.A2(n_823),
.B(n_807),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1021),
.B(n_783),
.Y(n_1086)
);

OAI21xp33_ASAP7_75t_L g1087 ( 
.A1(n_1035),
.A2(n_245),
.B(n_353),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_932),
.B(n_879),
.Y(n_1088)
);

OR2x6_ASAP7_75t_L g1089 ( 
.A(n_931),
.B(n_239),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_920),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_954),
.B(n_983),
.Y(n_1091)
);

CKINVDCx20_ASAP7_75t_R g1092 ( 
.A(n_968),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_949),
.A2(n_945),
.B(n_1034),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_931),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1023),
.B(n_14),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_934),
.A2(n_320),
.B(n_350),
.Y(n_1096)
);

NAND3xp33_ASAP7_75t_SL g1097 ( 
.A(n_924),
.B(n_247),
.C(n_254),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_SL g1098 ( 
.A1(n_999),
.A2(n_17),
.B(n_18),
.C(n_24),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_926),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_1060),
.B(n_255),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_1062),
.A2(n_17),
.B(n_18),
.C(n_24),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_988),
.B(n_25),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_928),
.A2(n_325),
.B(n_347),
.C(n_345),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_979),
.B(n_261),
.Y(n_1104)
);

O2A1O1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_1042),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_981),
.B(n_1071),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_1074),
.B(n_262),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_959),
.B(n_269),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_992),
.Y(n_1109)
);

NAND2xp33_ASAP7_75t_L g1110 ( 
.A(n_1002),
.B(n_941),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1018),
.B(n_32),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_1067),
.Y(n_1112)
);

O2A1O1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_1043),
.A2(n_46),
.B(n_48),
.C(n_49),
.Y(n_1113)
);

NAND2xp33_ASAP7_75t_R g1114 ( 
.A(n_1001),
.B(n_272),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_947),
.Y(n_1115)
);

O2A1O1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_966),
.A2(n_51),
.B(n_52),
.C(n_54),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_1064),
.Y(n_1117)
);

BUFx4f_ASAP7_75t_L g1118 ( 
.A(n_922),
.Y(n_1118)
);

NAND2x1_ASAP7_75t_L g1119 ( 
.A(n_940),
.B(n_377),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_992),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_944),
.A2(n_327),
.B(n_343),
.C(n_342),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1007),
.B(n_51),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1041),
.A2(n_282),
.B(n_333),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_916),
.A2(n_280),
.B(n_332),
.Y(n_1124)
);

BUFx8_ASAP7_75t_L g1125 ( 
.A(n_1053),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_915),
.B(n_55),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_922),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1048),
.A2(n_331),
.B(n_279),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_976),
.A2(n_278),
.B(n_275),
.C(n_377),
.Y(n_1129)
);

BUFx8_ASAP7_75t_L g1130 ( 
.A(n_1001),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_964),
.B(n_55),
.Y(n_1131)
);

NAND2x1_ASAP7_75t_L g1132 ( 
.A(n_940),
.B(n_377),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_935),
.A2(n_377),
.B(n_239),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_937),
.A2(n_377),
.B(n_109),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_1058),
.A2(n_975),
.B(n_957),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_918),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_SL g1137 ( 
.A(n_997),
.B(n_56),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_1015),
.A2(n_56),
.B(n_58),
.C(n_59),
.Y(n_1138)
);

INVx2_ASAP7_75t_SL g1139 ( 
.A(n_991),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_989),
.B(n_58),
.Y(n_1140)
);

AOI21x1_ASAP7_75t_L g1141 ( 
.A1(n_985),
.A2(n_108),
.B(n_190),
.Y(n_1141)
);

O2A1O1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_1054),
.A2(n_61),
.B(n_62),
.C(n_63),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1059),
.B(n_63),
.Y(n_1143)
);

AOI22x1_ASAP7_75t_L g1144 ( 
.A1(n_942),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1070),
.A2(n_64),
.B1(n_67),
.B2(n_68),
.Y(n_1145)
);

OR2x2_ASAP7_75t_L g1146 ( 
.A(n_1032),
.B(n_67),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_961),
.B(n_69),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_967),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_SL g1149 ( 
.A1(n_936),
.A2(n_70),
.B(n_71),
.C(n_72),
.Y(n_1149)
);

AOI221xp5_ASAP7_75t_L g1150 ( 
.A1(n_1070),
.A2(n_71),
.B1(n_74),
.B2(n_79),
.C(n_98),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1051),
.B(n_100),
.Y(n_1151)
);

CKINVDCx14_ASAP7_75t_R g1152 ( 
.A(n_922),
.Y(n_1152)
);

OAI21xp33_ASAP7_75t_SL g1153 ( 
.A1(n_956),
.A2(n_101),
.B(n_104),
.Y(n_1153)
);

NAND3xp33_ASAP7_75t_L g1154 ( 
.A(n_1008),
.B(n_114),
.C(n_116),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_SL g1155 ( 
.A1(n_1006),
.A2(n_130),
.B1(n_145),
.B2(n_152),
.Y(n_1155)
);

AOI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_1061),
.A2(n_1068),
.B1(n_1065),
.B2(n_939),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_994),
.B(n_163),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1058),
.A2(n_197),
.B(n_950),
.Y(n_1158)
);

AOI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1016),
.A2(n_1003),
.B1(n_978),
.B2(n_946),
.Y(n_1159)
);

NAND2x1p5_ASAP7_75t_L g1160 ( 
.A(n_1064),
.B(n_1045),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_990),
.B(n_1011),
.Y(n_1161)
);

NOR2x1_ASAP7_75t_SL g1162 ( 
.A(n_1005),
.B(n_1010),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_958),
.A2(n_1029),
.B1(n_1013),
.B2(n_1017),
.Y(n_1163)
);

O2A1O1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_1037),
.A2(n_929),
.B(n_1049),
.C(n_933),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_991),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_952),
.A2(n_953),
.B(n_971),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_R g1167 ( 
.A(n_991),
.B(n_1045),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_943),
.A2(n_914),
.B(n_977),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1044),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1002),
.B(n_951),
.Y(n_1170)
);

OAI22x1_ASAP7_75t_L g1171 ( 
.A1(n_1046),
.A2(n_1027),
.B1(n_962),
.B2(n_986),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1014),
.B(n_1056),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1014),
.Y(n_1173)
);

O2A1O1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_955),
.A2(n_1057),
.B(n_1055),
.C(n_1066),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_974),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_1045),
.Y(n_1176)
);

BUFx3_ASAP7_75t_L g1177 ( 
.A(n_974),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1004),
.B(n_980),
.Y(n_1178)
);

INVx6_ASAP7_75t_L g1179 ( 
.A(n_1002),
.Y(n_1179)
);

OR2x6_ASAP7_75t_L g1180 ( 
.A(n_969),
.B(n_970),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_1025),
.Y(n_1181)
);

INVxp33_ASAP7_75t_L g1182 ( 
.A(n_1009),
.Y(n_1182)
);

BUFx4f_ASAP7_75t_L g1183 ( 
.A(n_1002),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_930),
.Y(n_1184)
);

NOR3xp33_ASAP7_75t_SL g1185 ( 
.A(n_1078),
.B(n_1069),
.C(n_1076),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1000),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_919),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_987),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_984),
.A2(n_998),
.B(n_996),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1031),
.Y(n_1190)
);

OAI21xp33_ASAP7_75t_SL g1191 ( 
.A1(n_1026),
.A2(n_1033),
.B(n_1040),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_927),
.B(n_917),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_982),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1073),
.B(n_1076),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_1077),
.Y(n_1195)
);

BUFx4f_ASAP7_75t_L g1196 ( 
.A(n_1077),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_960),
.B(n_973),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_917),
.B(n_1022),
.Y(n_1198)
);

AOI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1075),
.A2(n_993),
.B1(n_1063),
.B2(n_1072),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1020),
.B(n_1031),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_972),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1050),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1036),
.B(n_1039),
.Y(n_1203)
);

O2A1O1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_1047),
.A2(n_1072),
.B(n_1063),
.C(n_1028),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1024),
.B(n_1028),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1030),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_1030),
.B(n_939),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_963),
.B(n_765),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_948),
.B(n_831),
.Y(n_1209)
);

AOI221x1_ASAP7_75t_L g1210 ( 
.A1(n_1145),
.A2(n_1080),
.B1(n_1140),
.B2(n_1138),
.C(n_1198),
.Y(n_1210)
);

OR2x6_ASAP7_75t_L g1211 ( 
.A(n_1179),
.B(n_1089),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1090),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1208),
.A2(n_1197),
.B(n_1168),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1099),
.Y(n_1214)
);

AOI221xp5_ASAP7_75t_SL g1215 ( 
.A1(n_1145),
.A2(n_1105),
.B1(n_1113),
.B2(n_1101),
.C(n_1142),
.Y(n_1215)
);

NAND3xp33_ASAP7_75t_L g1216 ( 
.A(n_1150),
.B(n_1137),
.C(n_1100),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_1092),
.Y(n_1217)
);

INVxp67_ASAP7_75t_L g1218 ( 
.A(n_1091),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1158),
.A2(n_1135),
.B(n_1093),
.Y(n_1219)
);

OA21x2_ASAP7_75t_L g1220 ( 
.A1(n_1189),
.A2(n_1203),
.B(n_1205),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1137),
.A2(n_1097),
.B1(n_1106),
.B2(n_1082),
.Y(n_1221)
);

AOI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1203),
.A2(n_1192),
.B(n_1205),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1174),
.A2(n_1172),
.B(n_1116),
.C(n_1194),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1088),
.B(n_1084),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_1126),
.B(n_1115),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1088),
.A2(n_1102),
.B(n_1087),
.C(n_1108),
.Y(n_1226)
);

O2A1O1Ixp33_ASAP7_75t_SL g1227 ( 
.A1(n_1122),
.A2(n_1121),
.B(n_1149),
.C(n_1103),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1166),
.A2(n_1191),
.B(n_1206),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1163),
.A2(n_1200),
.B(n_1122),
.Y(n_1229)
);

INVx2_ASAP7_75t_SL g1230 ( 
.A(n_1118),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1102),
.A2(n_1164),
.B(n_1111),
.C(n_1183),
.Y(n_1231)
);

NOR3xp33_ASAP7_75t_SL g1232 ( 
.A(n_1109),
.B(n_1131),
.C(n_1095),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_SL g1233 ( 
.A1(n_1098),
.A2(n_1131),
.B(n_1129),
.C(n_1170),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1118),
.Y(n_1234)
);

AOI221xp5_ASAP7_75t_SL g1235 ( 
.A1(n_1096),
.A2(n_1124),
.B1(n_1163),
.B2(n_1190),
.C(n_1143),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_1120),
.Y(n_1236)
);

OA21x2_ASAP7_75t_L g1237 ( 
.A1(n_1202),
.A2(n_1133),
.B(n_1193),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_L g1238 ( 
.A(n_1127),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1152),
.B(n_1182),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_1081),
.Y(n_1240)
);

AOI221xp5_ASAP7_75t_L g1241 ( 
.A1(n_1147),
.A2(n_1104),
.B1(n_1083),
.B2(n_1107),
.C(n_1156),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1112),
.B(n_1094),
.Y(n_1242)
);

NOR2xp67_ASAP7_75t_L g1243 ( 
.A(n_1139),
.B(n_1117),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1204),
.A2(n_1183),
.B(n_1134),
.Y(n_1244)
);

O2A1O1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_1153),
.A2(n_1143),
.B(n_1185),
.C(n_1173),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1159),
.B(n_1181),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1083),
.A2(n_1201),
.B(n_1184),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1136),
.B(n_1094),
.Y(n_1248)
);

AO31x2_ASAP7_75t_L g1249 ( 
.A1(n_1171),
.A2(n_1169),
.A3(n_1162),
.B(n_1151),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1127),
.Y(n_1250)
);

INVxp67_ASAP7_75t_L g1251 ( 
.A(n_1125),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1127),
.B(n_1117),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1123),
.A2(n_1128),
.B(n_1178),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1141),
.A2(n_1132),
.B(n_1119),
.Y(n_1254)
);

AOI221xp5_ASAP7_75t_SL g1255 ( 
.A1(n_1086),
.A2(n_1144),
.B1(n_1155),
.B2(n_1157),
.C(n_1161),
.Y(n_1255)
);

AOI221x1_ASAP7_75t_L g1256 ( 
.A1(n_1154),
.A2(n_1207),
.B1(n_1175),
.B2(n_1195),
.C(n_1148),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1079),
.A2(n_1196),
.B(n_1180),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1125),
.B(n_1176),
.Y(n_1258)
);

A2O1A1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1177),
.A2(n_1165),
.B(n_1195),
.C(n_1180),
.Y(n_1259)
);

AOI221xp5_ASAP7_75t_L g1260 ( 
.A1(n_1167),
.A2(n_1165),
.B1(n_1195),
.B2(n_1160),
.C(n_1114),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1130),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1090),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1090),
.Y(n_1263)
);

AO32x2_ASAP7_75t_L g1264 ( 
.A1(n_1145),
.A2(n_1163),
.A3(n_995),
.B1(n_1083),
.B2(n_884),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1110),
.A2(n_1208),
.B(n_921),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1158),
.A2(n_1135),
.B(n_1093),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_1118),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1110),
.A2(n_1208),
.B(n_921),
.Y(n_1268)
);

INVxp67_ASAP7_75t_SL g1269 ( 
.A(n_1181),
.Y(n_1269)
);

AO31x2_ASAP7_75t_L g1270 ( 
.A1(n_1085),
.A2(n_1019),
.A3(n_1194),
.B(n_1187),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1090),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1209),
.B(n_1091),
.Y(n_1272)
);

CKINVDCx11_ASAP7_75t_R g1273 ( 
.A(n_1092),
.Y(n_1273)
);

AO22x2_ASAP7_75t_L g1274 ( 
.A1(n_1126),
.A2(n_838),
.B1(n_1146),
.B2(n_1145),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1080),
.A2(n_1208),
.B(n_1198),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1110),
.A2(n_1208),
.B(n_921),
.Y(n_1276)
);

O2A1O1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1146),
.A2(n_662),
.B(n_623),
.C(n_765),
.Y(n_1277)
);

NAND3xp33_ASAP7_75t_SL g1278 ( 
.A(n_1146),
.B(n_662),
.C(n_567),
.Y(n_1278)
);

OAI22x1_ASAP7_75t_L g1279 ( 
.A1(n_1147),
.A2(n_948),
.B1(n_1126),
.B2(n_1146),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1208),
.B(n_765),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1158),
.A2(n_1135),
.B(n_1093),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1158),
.A2(n_1135),
.B(n_1093),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1208),
.B(n_765),
.Y(n_1283)
);

INVxp67_ASAP7_75t_SL g1284 ( 
.A(n_1181),
.Y(n_1284)
);

BUFx12f_ASAP7_75t_L g1285 ( 
.A(n_1109),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1209),
.B(n_948),
.Y(n_1286)
);

OR2x6_ASAP7_75t_L g1287 ( 
.A(n_1179),
.B(n_1089),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_SL g1288 ( 
.A1(n_1145),
.A2(n_948),
.B1(n_765),
.B2(n_662),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1208),
.B(n_765),
.Y(n_1289)
);

O2A1O1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1146),
.A2(n_662),
.B(n_623),
.C(n_765),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1110),
.A2(n_1208),
.B(n_921),
.Y(n_1291)
);

CKINVDCx20_ASAP7_75t_R g1292 ( 
.A(n_1092),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1090),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1208),
.A2(n_765),
.B1(n_662),
.B2(n_777),
.Y(n_1294)
);

BUFx10_ASAP7_75t_L g1295 ( 
.A(n_1109),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1158),
.A2(n_1135),
.B(n_1093),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1158),
.A2(n_1135),
.B(n_1093),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1090),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1158),
.A2(n_1135),
.B(n_1093),
.Y(n_1299)
);

AOI221x1_ASAP7_75t_L g1300 ( 
.A1(n_1145),
.A2(n_1080),
.B1(n_1140),
.B2(n_1138),
.C(n_1198),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1110),
.A2(n_1208),
.B(n_921),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1209),
.B(n_948),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1090),
.Y(n_1303)
);

AO32x2_ASAP7_75t_L g1304 ( 
.A1(n_1145),
.A2(n_1163),
.A3(n_995),
.B1(n_1083),
.B2(n_884),
.Y(n_1304)
);

INVxp67_ASAP7_75t_SL g1305 ( 
.A(n_1181),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1208),
.B(n_765),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1090),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1208),
.B(n_765),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_1208),
.B(n_1106),
.Y(n_1309)
);

AOI221xp5_ASAP7_75t_SL g1310 ( 
.A1(n_1080),
.A2(n_1145),
.B1(n_1138),
.B2(n_1113),
.C(n_1105),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1110),
.A2(n_1208),
.B(n_921),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1110),
.A2(n_1208),
.B(n_921),
.Y(n_1312)
);

OAI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1080),
.A2(n_1208),
.B(n_1198),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1179),
.Y(n_1314)
);

CKINVDCx11_ASAP7_75t_R g1315 ( 
.A(n_1092),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_SL g1316 ( 
.A1(n_1080),
.A2(n_724),
.B(n_1208),
.Y(n_1316)
);

AOI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1137),
.A2(n_948),
.B1(n_765),
.B2(n_1209),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1090),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1208),
.B(n_765),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1137),
.A2(n_948),
.B1(n_765),
.B2(n_1209),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_L g1321 ( 
.A(n_1209),
.B(n_948),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1090),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1080),
.A2(n_1208),
.B(n_1198),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1208),
.A2(n_765),
.B1(n_662),
.B2(n_777),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1112),
.Y(n_1325)
);

AOI221x1_ASAP7_75t_L g1326 ( 
.A1(n_1145),
.A2(n_1080),
.B1(n_1140),
.B2(n_1138),
.C(n_1198),
.Y(n_1326)
);

AOI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1137),
.A2(n_948),
.B1(n_765),
.B2(n_1209),
.Y(n_1327)
);

AOI31xp67_ASAP7_75t_L g1328 ( 
.A1(n_1197),
.A2(n_1188),
.A3(n_1199),
.B(n_1186),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1090),
.Y(n_1329)
);

AO31x2_ASAP7_75t_L g1330 ( 
.A1(n_1085),
.A2(n_1019),
.A3(n_1194),
.B(n_1187),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1090),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1110),
.A2(n_1208),
.B(n_921),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1208),
.A2(n_765),
.B1(n_662),
.B2(n_777),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1208),
.A2(n_765),
.B1(n_662),
.B2(n_777),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1209),
.B(n_1091),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1084),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1158),
.A2(n_1135),
.B(n_1093),
.Y(n_1337)
);

O2A1O1Ixp33_ASAP7_75t_SL g1338 ( 
.A1(n_1208),
.A2(n_1080),
.B(n_786),
.C(n_963),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_1092),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1110),
.A2(n_1208),
.B(n_921),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1208),
.B(n_765),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1208),
.B(n_765),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1110),
.A2(n_1208),
.B(n_921),
.Y(n_1343)
);

CKINVDCx6p67_ASAP7_75t_R g1344 ( 
.A(n_1092),
.Y(n_1344)
);

A2O1A1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1080),
.A2(n_777),
.B(n_689),
.C(n_691),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1208),
.B(n_765),
.Y(n_1346)
);

OAI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1317),
.A2(n_1327),
.B1(n_1320),
.B2(n_1216),
.Y(n_1347)
);

INVx8_ASAP7_75t_L g1348 ( 
.A(n_1292),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1272),
.B(n_1335),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1214),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1280),
.B(n_1283),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_SL g1352 ( 
.A1(n_1288),
.A2(n_1320),
.B1(n_1317),
.B2(n_1327),
.Y(n_1352)
);

INVx3_ASAP7_75t_L g1353 ( 
.A(n_1234),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1274),
.A2(n_1279),
.B1(n_1294),
.B2(n_1324),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1333),
.A2(n_1334),
.B1(n_1277),
.B2(n_1290),
.Y(n_1355)
);

BUFx8_ASAP7_75t_L g1356 ( 
.A(n_1285),
.Y(n_1356)
);

INVx6_ASAP7_75t_L g1357 ( 
.A(n_1234),
.Y(n_1357)
);

CKINVDCx20_ASAP7_75t_R g1358 ( 
.A(n_1273),
.Y(n_1358)
);

BUFx10_ASAP7_75t_L g1359 ( 
.A(n_1236),
.Y(n_1359)
);

CKINVDCx6p67_ASAP7_75t_R g1360 ( 
.A(n_1315),
.Y(n_1360)
);

AOI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1286),
.A2(n_1321),
.B1(n_1302),
.B2(n_1241),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1278),
.A2(n_1313),
.B1(n_1323),
.B2(n_1275),
.Y(n_1362)
);

CKINVDCx6p67_ASAP7_75t_R g1363 ( 
.A(n_1339),
.Y(n_1363)
);

CKINVDCx11_ASAP7_75t_R g1364 ( 
.A(n_1295),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1275),
.A2(n_1323),
.B1(n_1313),
.B2(n_1341),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1217),
.Y(n_1366)
);

INVx2_ASAP7_75t_SL g1367 ( 
.A(n_1240),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1289),
.A2(n_1346),
.B1(n_1342),
.B2(n_1306),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1221),
.A2(n_1308),
.B1(n_1319),
.B2(n_1345),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1221),
.A2(n_1229),
.B1(n_1225),
.B2(n_1309),
.Y(n_1370)
);

CKINVDCx11_ASAP7_75t_R g1371 ( 
.A(n_1295),
.Y(n_1371)
);

INVx4_ASAP7_75t_L g1372 ( 
.A(n_1344),
.Y(n_1372)
);

INVxp67_ASAP7_75t_L g1373 ( 
.A(n_1269),
.Y(n_1373)
);

OAI22xp33_ASAP7_75t_SL g1374 ( 
.A1(n_1246),
.A2(n_1218),
.B1(n_1224),
.B2(n_1304),
.Y(n_1374)
);

BUFx3_ASAP7_75t_L g1375 ( 
.A(n_1325),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1226),
.A2(n_1231),
.B1(n_1305),
.B2(n_1284),
.Y(n_1376)
);

BUFx10_ASAP7_75t_L g1377 ( 
.A(n_1242),
.Y(n_1377)
);

CKINVDCx11_ASAP7_75t_R g1378 ( 
.A(n_1261),
.Y(n_1378)
);

INVx6_ASAP7_75t_L g1379 ( 
.A(n_1267),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1248),
.B(n_1336),
.Y(n_1380)
);

INVx1_ASAP7_75t_SL g1381 ( 
.A(n_1239),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1229),
.A2(n_1264),
.B1(n_1304),
.B2(n_1247),
.Y(n_1382)
);

OAI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1210),
.A2(n_1326),
.B1(n_1300),
.B2(n_1304),
.Y(n_1383)
);

BUFx2_ASAP7_75t_R g1384 ( 
.A(n_1258),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1264),
.A2(n_1247),
.B1(n_1293),
.B2(n_1303),
.Y(n_1385)
);

INVx6_ASAP7_75t_L g1386 ( 
.A(n_1238),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1264),
.A2(n_1318),
.B1(n_1271),
.B2(n_1262),
.Y(n_1387)
);

INVx6_ASAP7_75t_L g1388 ( 
.A(n_1238),
.Y(n_1388)
);

INVx1_ASAP7_75t_SL g1389 ( 
.A(n_1250),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1263),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1298),
.A2(n_1331),
.B1(n_1329),
.B2(n_1322),
.Y(n_1391)
);

CKINVDCx6p67_ASAP7_75t_R g1392 ( 
.A(n_1238),
.Y(n_1392)
);

BUFx8_ASAP7_75t_L g1393 ( 
.A(n_1230),
.Y(n_1393)
);

CKINVDCx20_ASAP7_75t_R g1394 ( 
.A(n_1251),
.Y(n_1394)
);

BUFx8_ASAP7_75t_L g1395 ( 
.A(n_1307),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_SL g1396 ( 
.A1(n_1310),
.A2(n_1257),
.B1(n_1211),
.B2(n_1287),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1211),
.A2(n_1287),
.B1(n_1260),
.B2(n_1253),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1314),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_1232),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1243),
.B(n_1252),
.Y(n_1400)
);

OAI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1265),
.A2(n_1268),
.B1(n_1340),
.B2(n_1332),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1276),
.A2(n_1343),
.B1(n_1291),
.B2(n_1301),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1328),
.Y(n_1403)
);

INVx6_ASAP7_75t_L g1404 ( 
.A(n_1259),
.Y(n_1404)
);

AOI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1310),
.A2(n_1255),
.B1(n_1215),
.B2(n_1338),
.Y(n_1405)
);

CKINVDCx11_ASAP7_75t_R g1406 ( 
.A(n_1255),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1311),
.A2(n_1312),
.B1(n_1215),
.B2(n_1244),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1222),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1316),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1237),
.A2(n_1228),
.B1(n_1213),
.B2(n_1220),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1223),
.B(n_1249),
.Y(n_1411)
);

INVxp67_ASAP7_75t_SL g1412 ( 
.A(n_1220),
.Y(n_1412)
);

INVx3_ASAP7_75t_L g1413 ( 
.A(n_1270),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1227),
.A2(n_1235),
.B1(n_1233),
.B2(n_1330),
.Y(n_1414)
);

INVx1_ASAP7_75t_SL g1415 ( 
.A(n_1254),
.Y(n_1415)
);

BUFx10_ASAP7_75t_L g1416 ( 
.A(n_1235),
.Y(n_1416)
);

INVx6_ASAP7_75t_L g1417 ( 
.A(n_1256),
.Y(n_1417)
);

CKINVDCx11_ASAP7_75t_R g1418 ( 
.A(n_1245),
.Y(n_1418)
);

AOI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1219),
.A2(n_1337),
.B1(n_1281),
.B2(n_1282),
.Y(n_1419)
);

OAI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1266),
.A2(n_1296),
.B1(n_1297),
.B2(n_1299),
.Y(n_1420)
);

CKINVDCx6p67_ASAP7_75t_R g1421 ( 
.A(n_1273),
.Y(n_1421)
);

BUFx12f_ASAP7_75t_L g1422 ( 
.A(n_1273),
.Y(n_1422)
);

BUFx8_ASAP7_75t_L g1423 ( 
.A(n_1285),
.Y(n_1423)
);

BUFx8_ASAP7_75t_L g1424 ( 
.A(n_1285),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1212),
.Y(n_1425)
);

BUFx12f_ASAP7_75t_L g1426 ( 
.A(n_1273),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1212),
.Y(n_1427)
);

CKINVDCx11_ASAP7_75t_R g1428 ( 
.A(n_1273),
.Y(n_1428)
);

OAI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1317),
.A2(n_1327),
.B1(n_1320),
.B2(n_1137),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1212),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1280),
.B(n_1283),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_SL g1432 ( 
.A1(n_1274),
.A2(n_1288),
.B1(n_1137),
.B2(n_1216),
.Y(n_1432)
);

INVx6_ASAP7_75t_SL g1433 ( 
.A(n_1295),
.Y(n_1433)
);

INVx1_ASAP7_75t_SL g1434 ( 
.A(n_1292),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_SL g1435 ( 
.A1(n_1274),
.A2(n_1288),
.B1(n_1137),
.B2(n_1216),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_1273),
.Y(n_1436)
);

AOI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1288),
.A2(n_948),
.B1(n_1320),
.B2(n_1317),
.Y(n_1437)
);

OAI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1317),
.A2(n_1327),
.B1(n_1320),
.B2(n_1137),
.Y(n_1438)
);

OAI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1317),
.A2(n_1327),
.B1(n_1320),
.B2(n_1137),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1274),
.A2(n_1288),
.B1(n_1216),
.B2(n_1279),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1274),
.A2(n_1288),
.B1(n_1216),
.B2(n_1279),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1288),
.A2(n_1317),
.B1(n_1327),
.B2(n_1320),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1280),
.B(n_1283),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1280),
.B(n_1283),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1274),
.A2(n_1288),
.B1(n_1216),
.B2(n_1279),
.Y(n_1445)
);

BUFx5_ASAP7_75t_L g1446 ( 
.A(n_1212),
.Y(n_1446)
);

AOI21xp33_ASAP7_75t_L g1447 ( 
.A1(n_1216),
.A2(n_1290),
.B(n_1277),
.Y(n_1447)
);

BUFx10_ASAP7_75t_L g1448 ( 
.A(n_1236),
.Y(n_1448)
);

INVx2_ASAP7_75t_SL g1449 ( 
.A(n_1240),
.Y(n_1449)
);

OAI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1317),
.A2(n_1327),
.B1(n_1320),
.B2(n_1137),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1274),
.A2(n_1288),
.B1(n_1216),
.B2(n_1279),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1274),
.A2(n_1288),
.B1(n_1216),
.B2(n_1279),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1274),
.A2(n_1288),
.B1(n_1216),
.B2(n_1279),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1212),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_SL g1455 ( 
.A1(n_1274),
.A2(n_1288),
.B1(n_1137),
.B2(n_1216),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1280),
.B(n_1283),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1325),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1274),
.A2(n_1288),
.B1(n_1216),
.B2(n_1279),
.Y(n_1458)
);

BUFx8_ASAP7_75t_L g1459 ( 
.A(n_1285),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_SL g1460 ( 
.A(n_1317),
.B(n_1320),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1280),
.B(n_1283),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1212),
.Y(n_1462)
);

BUFx12f_ASAP7_75t_L g1463 ( 
.A(n_1273),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1288),
.A2(n_1317),
.B1(n_1327),
.B2(n_1320),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1274),
.A2(n_1288),
.B1(n_838),
.B2(n_961),
.Y(n_1465)
);

OAI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1317),
.A2(n_1327),
.B1(n_1320),
.B2(n_1137),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1212),
.Y(n_1467)
);

CKINVDCx11_ASAP7_75t_R g1468 ( 
.A(n_1273),
.Y(n_1468)
);

AOI22xp5_ASAP7_75t_SL g1469 ( 
.A1(n_1286),
.A2(n_1321),
.B1(n_1302),
.B2(n_1147),
.Y(n_1469)
);

BUFx10_ASAP7_75t_L g1470 ( 
.A(n_1236),
.Y(n_1470)
);

INVx2_ASAP7_75t_SL g1471 ( 
.A(n_1240),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1212),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1274),
.A2(n_1288),
.B1(n_1216),
.B2(n_1279),
.Y(n_1473)
);

AOI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1288),
.A2(n_948),
.B1(n_1320),
.B2(n_1317),
.Y(n_1474)
);

INVx1_ASAP7_75t_SL g1475 ( 
.A(n_1292),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1212),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1274),
.A2(n_1288),
.B1(n_1216),
.B2(n_1279),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1408),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1402),
.A2(n_1410),
.B(n_1407),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1373),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1446),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1382),
.B(n_1411),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_1457),
.Y(n_1483)
);

BUFx2_ASAP7_75t_SL g1484 ( 
.A(n_1446),
.Y(n_1484)
);

AOI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1355),
.A2(n_1403),
.B(n_1369),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1446),
.Y(n_1486)
);

OAI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1437),
.A2(n_1474),
.B1(n_1361),
.B2(n_1464),
.Y(n_1487)
);

NOR2x1_ASAP7_75t_SL g1488 ( 
.A(n_1376),
.B(n_1442),
.Y(n_1488)
);

INVx3_ASAP7_75t_L g1489 ( 
.A(n_1416),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1373),
.B(n_1460),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1409),
.Y(n_1491)
);

BUFx2_ASAP7_75t_L g1492 ( 
.A(n_1412),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1350),
.Y(n_1493)
);

BUFx3_ASAP7_75t_L g1494 ( 
.A(n_1375),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1390),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1425),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1427),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1430),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1454),
.B(n_1462),
.Y(n_1499)
);

BUFx12f_ASAP7_75t_L g1500 ( 
.A(n_1428),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1468),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1467),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1412),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1472),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1476),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1385),
.B(n_1387),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1385),
.B(n_1387),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1413),
.Y(n_1508)
);

BUFx2_ASAP7_75t_L g1509 ( 
.A(n_1415),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1416),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1365),
.B(n_1349),
.Y(n_1511)
);

AOI221xp5_ASAP7_75t_L g1512 ( 
.A1(n_1347),
.A2(n_1383),
.B1(n_1447),
.B2(n_1354),
.C(n_1445),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1432),
.A2(n_1455),
.B1(n_1435),
.B2(n_1465),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1404),
.Y(n_1514)
);

OAI21xp33_ASAP7_75t_SL g1515 ( 
.A1(n_1405),
.A2(n_1362),
.B(n_1365),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1419),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1391),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_1404),
.Y(n_1518)
);

INVx2_ASAP7_75t_SL g1519 ( 
.A(n_1386),
.Y(n_1519)
);

OAI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1362),
.A2(n_1347),
.B(n_1466),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1389),
.Y(n_1521)
);

INVxp67_ASAP7_75t_L g1522 ( 
.A(n_1380),
.Y(n_1522)
);

INVxp67_ASAP7_75t_SL g1523 ( 
.A(n_1407),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1417),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1418),
.Y(n_1525)
);

OR2x6_ASAP7_75t_L g1526 ( 
.A(n_1417),
.B(n_1404),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1354),
.B(n_1370),
.Y(n_1527)
);

BUFx2_ASAP7_75t_L g1528 ( 
.A(n_1352),
.Y(n_1528)
);

INVx1_ASAP7_75t_SL g1529 ( 
.A(n_1348),
.Y(n_1529)
);

BUFx2_ASAP7_75t_L g1530 ( 
.A(n_1392),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1432),
.B(n_1435),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1455),
.B(n_1370),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1351),
.B(n_1431),
.Y(n_1533)
);

INVxp67_ASAP7_75t_SL g1534 ( 
.A(n_1401),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1400),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1406),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1401),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_1386),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1420),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1420),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1440),
.B(n_1441),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1374),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1414),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1440),
.B(n_1441),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1381),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1429),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1429),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1438),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1443),
.B(n_1444),
.Y(n_1549)
);

CKINVDCx11_ASAP7_75t_R g1550 ( 
.A(n_1358),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1445),
.B(n_1451),
.Y(n_1551)
);

AO21x2_ASAP7_75t_L g1552 ( 
.A1(n_1439),
.A2(n_1450),
.B(n_1466),
.Y(n_1552)
);

AOI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1439),
.A2(n_1450),
.B(n_1451),
.Y(n_1553)
);

INVx2_ASAP7_75t_SL g1554 ( 
.A(n_1388),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1396),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1452),
.B(n_1453),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1396),
.Y(n_1557)
);

BUFx2_ASAP7_75t_L g1558 ( 
.A(n_1395),
.Y(n_1558)
);

BUFx2_ASAP7_75t_SL g1559 ( 
.A(n_1377),
.Y(n_1559)
);

INVx3_ASAP7_75t_L g1560 ( 
.A(n_1377),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1458),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1473),
.Y(n_1562)
);

OA21x2_ASAP7_75t_L g1563 ( 
.A1(n_1477),
.A2(n_1397),
.B(n_1368),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1398),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1456),
.B(n_1461),
.Y(n_1565)
);

AND2x2_ASAP7_75t_SL g1566 ( 
.A(n_1372),
.B(n_1368),
.Y(n_1566)
);

BUFx2_ASAP7_75t_L g1567 ( 
.A(n_1395),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1353),
.Y(n_1568)
);

INVx1_ASAP7_75t_SL g1569 ( 
.A(n_1348),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1393),
.Y(n_1570)
);

CKINVDCx20_ASAP7_75t_R g1571 ( 
.A(n_1360),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1469),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1422),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1511),
.B(n_1366),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1511),
.B(n_1372),
.Y(n_1575)
);

OAI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1515),
.A2(n_1399),
.B(n_1471),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1528),
.B(n_1475),
.Y(n_1577)
);

OAI21x1_ASAP7_75t_SL g1578 ( 
.A1(n_1488),
.A2(n_1367),
.B(n_1449),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1483),
.B(n_1363),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1531),
.A2(n_1378),
.B1(n_1348),
.B2(n_1434),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1524),
.B(n_1436),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1565),
.B(n_1421),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1483),
.B(n_1384),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1483),
.B(n_1384),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_SL g1585 ( 
.A1(n_1531),
.A2(n_1463),
.B1(n_1426),
.B2(n_1379),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1522),
.B(n_1470),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1565),
.B(n_1393),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1494),
.B(n_1470),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1480),
.B(n_1493),
.Y(n_1589)
);

OA21x2_ASAP7_75t_L g1590 ( 
.A1(n_1479),
.A2(n_1379),
.B(n_1357),
.Y(n_1590)
);

BUFx3_ASAP7_75t_L g1591 ( 
.A(n_1530),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1524),
.B(n_1394),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1533),
.B(n_1364),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1482),
.B(n_1448),
.Y(n_1594)
);

INVx1_ASAP7_75t_SL g1595 ( 
.A(n_1529),
.Y(n_1595)
);

A2O1A1Ixp33_ASAP7_75t_L g1596 ( 
.A1(n_1553),
.A2(n_1433),
.B(n_1371),
.C(n_1424),
.Y(n_1596)
);

AOI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1532),
.A2(n_1356),
.B1(n_1423),
.B2(n_1424),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1549),
.B(n_1359),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_SL g1599 ( 
.A(n_1570),
.Y(n_1599)
);

O2A1O1Ixp33_ASAP7_75t_L g1600 ( 
.A1(n_1487),
.A2(n_1359),
.B(n_1448),
.C(n_1459),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1499),
.B(n_1534),
.Y(n_1601)
);

AOI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1520),
.A2(n_1356),
.B(n_1423),
.Y(n_1602)
);

AOI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1532),
.A2(n_1528),
.B1(n_1513),
.B2(n_1512),
.Y(n_1603)
);

A2O1A1Ixp33_ASAP7_75t_L g1604 ( 
.A1(n_1515),
.A2(n_1527),
.B(n_1544),
.C(n_1556),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1492),
.Y(n_1605)
);

AOI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1488),
.A2(n_1552),
.B(n_1523),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1490),
.B(n_1521),
.Y(n_1607)
);

AND3x1_ASAP7_75t_L g1608 ( 
.A(n_1536),
.B(n_1500),
.C(n_1550),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1535),
.B(n_1564),
.Y(n_1609)
);

OR2x6_ASAP7_75t_L g1610 ( 
.A(n_1526),
.B(n_1484),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_SL g1611 ( 
.A1(n_1544),
.A2(n_1556),
.B1(n_1551),
.B2(n_1541),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1502),
.B(n_1504),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1504),
.B(n_1505),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_L g1614 ( 
.A(n_1566),
.B(n_1510),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1505),
.B(n_1546),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1545),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1560),
.B(n_1552),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1495),
.B(n_1496),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1560),
.B(n_1546),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_SL g1620 ( 
.A(n_1500),
.B(n_1573),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1492),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1560),
.B(n_1547),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1495),
.Y(n_1623)
);

AO32x2_ASAP7_75t_L g1624 ( 
.A1(n_1519),
.A2(n_1538),
.A3(n_1554),
.B1(n_1507),
.B2(n_1506),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1548),
.B(n_1568),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1497),
.B(n_1498),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1537),
.B(n_1498),
.Y(n_1627)
);

NOR3xp33_ASAP7_75t_SL g1628 ( 
.A(n_1501),
.B(n_1516),
.C(n_1540),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1503),
.Y(n_1629)
);

AO21x2_ASAP7_75t_L g1630 ( 
.A1(n_1485),
.A2(n_1539),
.B(n_1516),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1489),
.B(n_1559),
.Y(n_1631)
);

OA21x2_ASAP7_75t_L g1632 ( 
.A1(n_1543),
.A2(n_1503),
.B(n_1508),
.Y(n_1632)
);

OAI22xp5_ASAP7_75t_SL g1633 ( 
.A1(n_1525),
.A2(n_1567),
.B1(n_1558),
.B2(n_1536),
.Y(n_1633)
);

INVx2_ASAP7_75t_SL g1634 ( 
.A(n_1568),
.Y(n_1634)
);

O2A1O1Ixp33_ASAP7_75t_SL g1635 ( 
.A1(n_1569),
.A2(n_1571),
.B(n_1489),
.C(n_1543),
.Y(n_1635)
);

INVxp33_ASAP7_75t_SL g1636 ( 
.A(n_1620),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1605),
.B(n_1478),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1624),
.B(n_1481),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1624),
.B(n_1617),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1624),
.B(n_1486),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1624),
.B(n_1486),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1632),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1632),
.Y(n_1643)
);

INVx1_ASAP7_75t_SL g1644 ( 
.A(n_1632),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1603),
.A2(n_1563),
.B1(n_1562),
.B2(n_1561),
.Y(n_1645)
);

BUFx2_ASAP7_75t_L g1646 ( 
.A(n_1621),
.Y(n_1646)
);

INVxp67_ASAP7_75t_SL g1647 ( 
.A(n_1621),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1629),
.B(n_1509),
.Y(n_1648)
);

OAI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1604),
.A2(n_1555),
.B1(n_1557),
.B2(n_1572),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1623),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1627),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1601),
.B(n_1619),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_SL g1653 ( 
.A(n_1606),
.B(n_1489),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1627),
.Y(n_1654)
);

BUFx3_ASAP7_75t_L g1655 ( 
.A(n_1578),
.Y(n_1655)
);

BUFx3_ASAP7_75t_L g1656 ( 
.A(n_1610),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1626),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1622),
.B(n_1625),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1589),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1618),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1616),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1607),
.Y(n_1662)
);

NOR2x1_ASAP7_75t_L g1663 ( 
.A(n_1631),
.B(n_1491),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1630),
.B(n_1634),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1643),
.Y(n_1665)
);

AOI221xp5_ASAP7_75t_L g1666 ( 
.A1(n_1649),
.A2(n_1604),
.B1(n_1580),
.B2(n_1576),
.C(n_1611),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1643),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1650),
.Y(n_1668)
);

AOI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1649),
.A2(n_1542),
.B1(n_1555),
.B2(n_1557),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1650),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1646),
.Y(n_1671)
);

AND4x1_ASAP7_75t_L g1672 ( 
.A(n_1663),
.B(n_1596),
.C(n_1602),
.D(n_1597),
.Y(n_1672)
);

INVxp67_ASAP7_75t_L g1673 ( 
.A(n_1664),
.Y(n_1673)
);

INVxp67_ASAP7_75t_L g1674 ( 
.A(n_1664),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1657),
.B(n_1594),
.Y(n_1675)
);

INVx4_ASAP7_75t_L g1676 ( 
.A(n_1655),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1643),
.Y(n_1677)
);

OAI211xp5_ASAP7_75t_SL g1678 ( 
.A1(n_1653),
.A2(n_1600),
.B(n_1598),
.C(n_1580),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1646),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1646),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1643),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1638),
.B(n_1640),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1638),
.B(n_1575),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1650),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1650),
.Y(n_1685)
);

INVx4_ASAP7_75t_L g1686 ( 
.A(n_1655),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1643),
.Y(n_1687)
);

AOI221xp5_ASAP7_75t_L g1688 ( 
.A1(n_1649),
.A2(n_1572),
.B1(n_1577),
.B2(n_1596),
.C(n_1628),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1638),
.B(n_1640),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1640),
.B(n_1594),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1651),
.B(n_1609),
.Y(n_1691)
);

INVx3_ASAP7_75t_L g1692 ( 
.A(n_1655),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1657),
.B(n_1574),
.Y(n_1693)
);

INVxp67_ASAP7_75t_SL g1694 ( 
.A(n_1642),
.Y(n_1694)
);

OAI31xp33_ASAP7_75t_L g1695 ( 
.A1(n_1645),
.A2(n_1614),
.A3(n_1542),
.B(n_1577),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1637),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1657),
.B(n_1614),
.Y(n_1697)
);

BUFx2_ASAP7_75t_L g1698 ( 
.A(n_1655),
.Y(n_1698)
);

NAND3xp33_ASAP7_75t_L g1699 ( 
.A(n_1661),
.B(n_1628),
.C(n_1585),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1641),
.B(n_1590),
.Y(n_1700)
);

INVx1_ASAP7_75t_SL g1701 ( 
.A(n_1648),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1637),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1639),
.B(n_1590),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1637),
.B(n_1615),
.Y(n_1704)
);

INVx3_ASAP7_75t_L g1705 ( 
.A(n_1655),
.Y(n_1705)
);

AOI221xp5_ASAP7_75t_L g1706 ( 
.A1(n_1639),
.A2(n_1525),
.B1(n_1608),
.B2(n_1517),
.C(n_1635),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1647),
.B(n_1612),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1639),
.B(n_1590),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_SL g1709 ( 
.A1(n_1639),
.A2(n_1525),
.B1(n_1514),
.B2(n_1518),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1652),
.B(n_1581),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1654),
.B(n_1613),
.Y(n_1711)
);

AOI33xp33_ASAP7_75t_L g1712 ( 
.A1(n_1644),
.A2(n_1595),
.A3(n_1586),
.B1(n_1583),
.B2(n_1584),
.B3(n_1579),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1665),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1710),
.B(n_1652),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1668),
.Y(n_1715)
);

HB1xp67_ASAP7_75t_L g1716 ( 
.A(n_1671),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1676),
.B(n_1663),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1701),
.B(n_1659),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1710),
.B(n_1652),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1678),
.B(n_1636),
.Y(n_1720)
);

BUFx2_ASAP7_75t_L g1721 ( 
.A(n_1676),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1670),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1697),
.B(n_1662),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1697),
.B(n_1662),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1710),
.B(n_1652),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1665),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1701),
.B(n_1659),
.Y(n_1727)
);

BUFx2_ASAP7_75t_L g1728 ( 
.A(n_1676),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1678),
.B(n_1636),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1696),
.B(n_1660),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1690),
.B(n_1658),
.Y(n_1731)
);

AND2x2_ASAP7_75t_SL g1732 ( 
.A(n_1688),
.B(n_1525),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1704),
.B(n_1654),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1704),
.B(n_1654),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1676),
.B(n_1663),
.Y(n_1735)
);

INVxp67_ASAP7_75t_SL g1736 ( 
.A(n_1673),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1665),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1670),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1684),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1690),
.B(n_1658),
.Y(n_1740)
);

AND2x4_ASAP7_75t_L g1741 ( 
.A(n_1686),
.B(n_1656),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1684),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1711),
.B(n_1654),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1690),
.B(n_1658),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1685),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1711),
.B(n_1654),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1675),
.B(n_1661),
.Y(n_1747)
);

BUFx2_ASAP7_75t_L g1748 ( 
.A(n_1686),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1682),
.B(n_1689),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1667),
.Y(n_1750)
);

NOR2x1_ASAP7_75t_L g1751 ( 
.A(n_1686),
.B(n_1699),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1682),
.B(n_1658),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1667),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1675),
.B(n_1648),
.Y(n_1754)
);

INVx1_ASAP7_75t_SL g1755 ( 
.A(n_1698),
.Y(n_1755)
);

INVxp67_ASAP7_75t_L g1756 ( 
.A(n_1699),
.Y(n_1756)
);

INVx1_ASAP7_75t_SL g1757 ( 
.A(n_1698),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1667),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1686),
.B(n_1656),
.Y(n_1759)
);

INVx3_ASAP7_75t_L g1760 ( 
.A(n_1692),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1696),
.B(n_1660),
.Y(n_1761)
);

AND2x4_ASAP7_75t_L g1762 ( 
.A(n_1749),
.B(n_1692),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1716),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1730),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1723),
.B(n_1702),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1756),
.B(n_1712),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1752),
.B(n_1682),
.Y(n_1767)
);

HB1xp67_ASAP7_75t_L g1768 ( 
.A(n_1736),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1724),
.B(n_1702),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1730),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1752),
.B(n_1689),
.Y(n_1771)
);

NOR3xp33_ASAP7_75t_L g1772 ( 
.A(n_1751),
.B(n_1688),
.C(n_1706),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1713),
.Y(n_1773)
);

INVxp67_ASAP7_75t_SL g1774 ( 
.A(n_1751),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1747),
.B(n_1693),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1761),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1720),
.B(n_1693),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1761),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1718),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1729),
.B(n_1671),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1732),
.B(n_1679),
.Y(n_1781)
);

INVx2_ASAP7_75t_SL g1782 ( 
.A(n_1741),
.Y(n_1782)
);

OAI221xp5_ASAP7_75t_L g1783 ( 
.A1(n_1743),
.A2(n_1695),
.B1(n_1666),
.B2(n_1706),
.C(n_1669),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1713),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1732),
.B(n_1679),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1754),
.B(n_1718),
.Y(n_1786)
);

AND2x4_ASAP7_75t_L g1787 ( 
.A(n_1749),
.B(n_1692),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1732),
.B(n_1755),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1755),
.B(n_1672),
.Y(n_1789)
);

INVx1_ASAP7_75t_SL g1790 ( 
.A(n_1757),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1731),
.B(n_1740),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1731),
.B(n_1689),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1754),
.B(n_1691),
.Y(n_1793)
);

NOR2x1p5_ASAP7_75t_SL g1794 ( 
.A(n_1713),
.B(n_1726),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1727),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1727),
.Y(n_1796)
);

AND2x4_ASAP7_75t_L g1797 ( 
.A(n_1741),
.B(n_1692),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1757),
.B(n_1680),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1715),
.Y(n_1799)
);

INVxp67_ASAP7_75t_L g1800 ( 
.A(n_1721),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1714),
.B(n_1719),
.Y(n_1801)
);

INVx5_ASAP7_75t_L g1802 ( 
.A(n_1721),
.Y(n_1802)
);

OAI21xp33_ASAP7_75t_SL g1803 ( 
.A1(n_1740),
.A2(n_1705),
.B(n_1683),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1726),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1726),
.Y(n_1805)
);

NOR2x1p5_ASAP7_75t_L g1806 ( 
.A(n_1741),
.B(n_1570),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1733),
.B(n_1734),
.Y(n_1807)
);

INVx3_ASAP7_75t_L g1808 ( 
.A(n_1717),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1733),
.B(n_1691),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1737),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1715),
.Y(n_1811)
);

INVxp67_ASAP7_75t_L g1812 ( 
.A(n_1728),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1773),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1799),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1790),
.B(n_1714),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1806),
.B(n_1741),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1791),
.B(n_1759),
.Y(n_1817)
);

AND2x4_ASAP7_75t_SL g1818 ( 
.A(n_1797),
.B(n_1759),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1811),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1786),
.B(n_1734),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1773),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1779),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1791),
.B(n_1759),
.Y(n_1823)
);

HB1xp67_ASAP7_75t_L g1824 ( 
.A(n_1768),
.Y(n_1824)
);

BUFx3_ASAP7_75t_L g1825 ( 
.A(n_1768),
.Y(n_1825)
);

NOR2xp33_ASAP7_75t_L g1826 ( 
.A(n_1789),
.B(n_1599),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1766),
.B(n_1719),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1786),
.B(n_1795),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1763),
.B(n_1725),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1796),
.B(n_1743),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1765),
.B(n_1746),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1789),
.B(n_1759),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1784),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1792),
.B(n_1744),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1772),
.B(n_1725),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1777),
.B(n_1744),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1765),
.B(n_1746),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1784),
.Y(n_1838)
);

BUFx2_ASAP7_75t_L g1839 ( 
.A(n_1774),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1800),
.B(n_1728),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_SL g1841 ( 
.A(n_1797),
.B(n_1717),
.Y(n_1841)
);

INVxp67_ASAP7_75t_L g1842 ( 
.A(n_1780),
.Y(n_1842)
);

AOI32xp33_ASAP7_75t_L g1843 ( 
.A1(n_1783),
.A2(n_1666),
.A3(n_1703),
.B1(n_1708),
.B2(n_1644),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1804),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1793),
.B(n_1707),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1804),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1805),
.Y(n_1847)
);

NOR3xp33_ASAP7_75t_L g1848 ( 
.A(n_1808),
.B(n_1633),
.C(n_1748),
.Y(n_1848)
);

INVx1_ASAP7_75t_SL g1849 ( 
.A(n_1782),
.Y(n_1849)
);

AOI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1788),
.A2(n_1695),
.B(n_1748),
.Y(n_1850)
);

INVx1_ASAP7_75t_SL g1851 ( 
.A(n_1782),
.Y(n_1851)
);

A2O1A1Ixp33_ASAP7_75t_L g1852 ( 
.A1(n_1794),
.A2(n_1708),
.B(n_1703),
.C(n_1700),
.Y(n_1852)
);

OAI22xp5_ASAP7_75t_L g1853 ( 
.A1(n_1801),
.A2(n_1709),
.B1(n_1735),
.B2(n_1717),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1824),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_SL g1855 ( 
.A(n_1843),
.B(n_1802),
.Y(n_1855)
);

NAND3xp33_ASAP7_75t_L g1856 ( 
.A(n_1843),
.B(n_1812),
.C(n_1802),
.Y(n_1856)
);

INVx2_ASAP7_75t_SL g1857 ( 
.A(n_1818),
.Y(n_1857)
);

OAI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1835),
.A2(n_1781),
.B1(n_1785),
.B2(n_1644),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1825),
.B(n_1764),
.Y(n_1859)
);

AND2x4_ASAP7_75t_L g1860 ( 
.A(n_1832),
.B(n_1825),
.Y(n_1860)
);

AOI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1826),
.A2(n_1708),
.B1(n_1703),
.B2(n_1645),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1817),
.Y(n_1862)
);

AOI222xp33_ASAP7_75t_L g1863 ( 
.A1(n_1839),
.A2(n_1842),
.B1(n_1827),
.B2(n_1852),
.C1(n_1822),
.C2(n_1853),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1828),
.Y(n_1864)
);

NAND3xp33_ASAP7_75t_L g1865 ( 
.A(n_1839),
.B(n_1802),
.C(n_1798),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1828),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1849),
.B(n_1770),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1832),
.B(n_1797),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1851),
.B(n_1776),
.Y(n_1869)
);

OAI22xp33_ASAP7_75t_L g1870 ( 
.A1(n_1850),
.A2(n_1822),
.B1(n_1820),
.B2(n_1815),
.Y(n_1870)
);

INVxp67_ASAP7_75t_SL g1871 ( 
.A(n_1840),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1836),
.B(n_1778),
.Y(n_1872)
);

OAI21xp5_ASAP7_75t_SL g1873 ( 
.A1(n_1848),
.A2(n_1672),
.B(n_1808),
.Y(n_1873)
);

OAI32xp33_ASAP7_75t_L g1874 ( 
.A1(n_1820),
.A2(n_1803),
.A3(n_1808),
.B1(n_1807),
.B2(n_1760),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1845),
.B(n_1775),
.Y(n_1875)
);

AOI221xp5_ASAP7_75t_L g1876 ( 
.A1(n_1814),
.A2(n_1819),
.B1(n_1846),
.B2(n_1833),
.C(n_1694),
.Y(n_1876)
);

OAI31xp33_ASAP7_75t_L g1877 ( 
.A1(n_1833),
.A2(n_1700),
.A3(n_1694),
.B(n_1681),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1814),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1817),
.B(n_1792),
.Y(n_1879)
);

INVx1_ASAP7_75t_SL g1880 ( 
.A(n_1818),
.Y(n_1880)
);

A2O1A1Ixp33_ASAP7_75t_SL g1881 ( 
.A1(n_1819),
.A2(n_1816),
.B(n_1760),
.C(n_1813),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1864),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1870),
.B(n_1834),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1871),
.B(n_1834),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1866),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1868),
.B(n_1823),
.Y(n_1886)
);

OR2x2_ASAP7_75t_L g1887 ( 
.A(n_1875),
.B(n_1829),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1878),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1871),
.B(n_1860),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1854),
.Y(n_1890)
);

OAI32xp33_ASAP7_75t_L g1891 ( 
.A1(n_1855),
.A2(n_1831),
.A3(n_1837),
.B1(n_1830),
.B2(n_1841),
.Y(n_1891)
);

OAI22xp33_ASAP7_75t_L g1892 ( 
.A1(n_1861),
.A2(n_1845),
.B1(n_1830),
.B2(n_1837),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1860),
.B(n_1823),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1859),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1867),
.Y(n_1895)
);

AOI22xp5_ASAP7_75t_L g1896 ( 
.A1(n_1870),
.A2(n_1821),
.B1(n_1838),
.B2(n_1813),
.Y(n_1896)
);

AOI22xp5_ASAP7_75t_L g1897 ( 
.A1(n_1863),
.A2(n_1838),
.B1(n_1844),
.B2(n_1821),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1869),
.Y(n_1898)
);

A2O1A1Ixp33_ASAP7_75t_L g1899 ( 
.A1(n_1855),
.A2(n_1856),
.B(n_1873),
.C(n_1881),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1872),
.Y(n_1900)
);

OAI32xp33_ASAP7_75t_L g1901 ( 
.A1(n_1865),
.A2(n_1831),
.A3(n_1816),
.B1(n_1807),
.B2(n_1760),
.Y(n_1901)
);

OAI21xp33_ASAP7_75t_L g1902 ( 
.A1(n_1880),
.A2(n_1857),
.B(n_1862),
.Y(n_1902)
);

AOI22xp5_ASAP7_75t_L g1903 ( 
.A1(n_1858),
.A2(n_1847),
.B1(n_1844),
.B2(n_1846),
.Y(n_1903)
);

OAI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1858),
.A2(n_1802),
.B1(n_1735),
.B2(n_1717),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1884),
.B(n_1879),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_SL g1906 ( 
.A(n_1889),
.B(n_1735),
.Y(n_1906)
);

AOI21xp33_ASAP7_75t_L g1907 ( 
.A1(n_1891),
.A2(n_1881),
.B(n_1876),
.Y(n_1907)
);

OAI21xp5_ASAP7_75t_L g1908 ( 
.A1(n_1899),
.A2(n_1874),
.B(n_1877),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_SL g1909 ( 
.A(n_1904),
.B(n_1893),
.Y(n_1909)
);

OR2x2_ASAP7_75t_L g1910 ( 
.A(n_1883),
.B(n_1809),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1887),
.Y(n_1911)
);

AND2x2_ASAP7_75t_SL g1912 ( 
.A(n_1883),
.B(n_1558),
.Y(n_1912)
);

OAI322xp33_ASAP7_75t_L g1913 ( 
.A1(n_1895),
.A2(n_1847),
.A3(n_1673),
.B1(n_1674),
.B2(n_1769),
.C1(n_1810),
.C2(n_1805),
.Y(n_1913)
);

AO22x2_ASAP7_75t_L g1914 ( 
.A1(n_1890),
.A2(n_1810),
.B1(n_1593),
.B2(n_1582),
.Y(n_1914)
);

O2A1O1Ixp33_ASAP7_75t_L g1915 ( 
.A1(n_1904),
.A2(n_1674),
.B(n_1687),
.C(n_1677),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1886),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1882),
.Y(n_1917)
);

OA211x2_ASAP7_75t_L g1918 ( 
.A1(n_1902),
.A2(n_1653),
.B(n_1587),
.C(n_1631),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1885),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1888),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_SL g1921 ( 
.A(n_1912),
.B(n_1908),
.Y(n_1921)
);

AOI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1907),
.A2(n_1908),
.B(n_1909),
.Y(n_1922)
);

OAI21xp33_ASAP7_75t_L g1923 ( 
.A1(n_1907),
.A2(n_1898),
.B(n_1894),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1911),
.Y(n_1924)
);

OAI21xp5_ASAP7_75t_L g1925 ( 
.A1(n_1905),
.A2(n_1897),
.B(n_1896),
.Y(n_1925)
);

NAND3xp33_ASAP7_75t_L g1926 ( 
.A(n_1917),
.B(n_1919),
.C(n_1920),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_SL g1927 ( 
.A(n_1916),
.B(n_1910),
.Y(n_1927)
);

NOR2xp33_ASAP7_75t_L g1928 ( 
.A(n_1906),
.B(n_1900),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1914),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_L g1930 ( 
.A(n_1913),
.B(n_1901),
.Y(n_1930)
);

NAND4xp25_ASAP7_75t_SL g1931 ( 
.A(n_1915),
.B(n_1903),
.C(n_1892),
.D(n_1771),
.Y(n_1931)
);

OAI22xp5_ASAP7_75t_L g1932 ( 
.A1(n_1922),
.A2(n_1921),
.B1(n_1930),
.B2(n_1927),
.Y(n_1932)
);

NOR3xp33_ASAP7_75t_L g1933 ( 
.A(n_1923),
.B(n_1913),
.C(n_1567),
.Y(n_1933)
);

AOI222xp33_ASAP7_75t_L g1934 ( 
.A1(n_1929),
.A2(n_1914),
.B1(n_1700),
.B2(n_1687),
.C1(n_1681),
.C2(n_1677),
.Y(n_1934)
);

XOR2x2_ASAP7_75t_SL g1935 ( 
.A(n_1924),
.B(n_1918),
.Y(n_1935)
);

O2A1O1Ixp33_ASAP7_75t_L g1936 ( 
.A1(n_1925),
.A2(n_1681),
.B(n_1677),
.C(n_1687),
.Y(n_1936)
);

AOI211xp5_ASAP7_75t_L g1937 ( 
.A1(n_1931),
.A2(n_1570),
.B(n_1735),
.C(n_1635),
.Y(n_1937)
);

OAI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1926),
.A2(n_1787),
.B(n_1762),
.Y(n_1938)
);

AOI211xp5_ASAP7_75t_L g1939 ( 
.A1(n_1932),
.A2(n_1928),
.B(n_1767),
.C(n_1771),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1935),
.Y(n_1940)
);

NOR3xp33_ASAP7_75t_SL g1941 ( 
.A(n_1938),
.B(n_1647),
.C(n_1707),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_SL g1942 ( 
.A(n_1933),
.B(n_1760),
.Y(n_1942)
);

AOI221xp5_ASAP7_75t_L g1943 ( 
.A1(n_1936),
.A2(n_1753),
.B1(n_1737),
.B2(n_1750),
.C(n_1758),
.Y(n_1943)
);

AOI221xp5_ASAP7_75t_L g1944 ( 
.A1(n_1937),
.A2(n_1753),
.B1(n_1737),
.B2(n_1750),
.C(n_1758),
.Y(n_1944)
);

OAI221xp5_ASAP7_75t_L g1945 ( 
.A1(n_1934),
.A2(n_1750),
.B1(n_1753),
.B2(n_1758),
.C(n_1709),
.Y(n_1945)
);

NOR2x1_ASAP7_75t_L g1946 ( 
.A(n_1932),
.B(n_1762),
.Y(n_1946)
);

OAI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1940),
.A2(n_1787),
.B1(n_1762),
.B2(n_1767),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1946),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1942),
.Y(n_1949)
);

NOR2x1_ASAP7_75t_L g1950 ( 
.A(n_1945),
.B(n_1787),
.Y(n_1950)
);

OR2x2_ASAP7_75t_L g1951 ( 
.A(n_1939),
.B(n_1680),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1941),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1944),
.B(n_1705),
.Y(n_1953)
);

CKINVDCx20_ASAP7_75t_R g1954 ( 
.A(n_1948),
.Y(n_1954)
);

AOI21xp5_ASAP7_75t_L g1955 ( 
.A1(n_1952),
.A2(n_1943),
.B(n_1722),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1949),
.B(n_1950),
.Y(n_1956)
);

OAI211xp5_ASAP7_75t_SL g1957 ( 
.A1(n_1951),
.A2(n_1705),
.B(n_1745),
.C(n_1742),
.Y(n_1957)
);

XNOR2x1_ASAP7_75t_L g1958 ( 
.A(n_1953),
.B(n_1592),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1954),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1956),
.B(n_1958),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1959),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1961),
.Y(n_1962)
);

AOI21xp5_ASAP7_75t_L g1963 ( 
.A1(n_1961),
.A2(n_1960),
.B(n_1955),
.Y(n_1963)
);

NOR2x1p5_ASAP7_75t_L g1964 ( 
.A(n_1962),
.B(n_1957),
.Y(n_1964)
);

BUFx2_ASAP7_75t_L g1965 ( 
.A(n_1963),
.Y(n_1965)
);

OAI22xp33_ASAP7_75t_L g1966 ( 
.A1(n_1965),
.A2(n_1947),
.B1(n_1705),
.B2(n_1745),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1966),
.B(n_1964),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1967),
.Y(n_1968)
);

INVxp67_ASAP7_75t_L g1969 ( 
.A(n_1968),
.Y(n_1969)
);

AOI221xp5_ASAP7_75t_L g1970 ( 
.A1(n_1969),
.A2(n_1588),
.B1(n_1742),
.B2(n_1739),
.C(n_1738),
.Y(n_1970)
);

AOI211xp5_ASAP7_75t_L g1971 ( 
.A1(n_1970),
.A2(n_1530),
.B(n_1591),
.C(n_1592),
.Y(n_1971)
);


endmodule