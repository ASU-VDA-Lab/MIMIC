module real_jpeg_26273_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_3),
.A2(n_21),
.B1(n_22),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_3),
.A2(n_33),
.B1(n_38),
.B2(n_42),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_3),
.A2(n_33),
.B1(n_53),
.B2(n_57),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_3),
.A2(n_33),
.B1(n_59),
.B2(n_67),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_4),
.A2(n_38),
.B1(n_42),
.B2(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_4),
.A2(n_45),
.B1(n_60),
.B2(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_4),
.A2(n_45),
.B1(n_53),
.B2(n_57),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_4),
.A2(n_56),
.B(n_104),
.C(n_105),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_4),
.B(n_52),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_4),
.A2(n_21),
.B1(n_22),
.B2(n_45),
.Y(n_124)
);

O2A1O1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_4),
.A2(n_57),
.B(n_78),
.C(n_133),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_4),
.B(n_22),
.C(n_41),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_4),
.B(n_84),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_4),
.B(n_30),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_4),
.B(n_43),
.Y(n_181)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_6),
.Y(n_78)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_8),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_58)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_8),
.A2(n_53),
.B1(n_57),
.B2(n_61),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_8),
.A2(n_38),
.B1(n_42),
.B2(n_61),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_8),
.A2(n_21),
.B1(n_22),
.B2(n_61),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_10),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_11),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_11),
.B(n_166),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_126),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_125),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_111),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_15),
.B(n_111),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_17),
.B1(n_88),
.B2(n_110),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_48),
.B1(n_86),
.B2(n_87),
.Y(n_17)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_34),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_25),
.B(n_27),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_20),
.A2(n_108),
.B(n_109),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_21),
.A2(n_22),
.B1(n_40),
.B2(n_41),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_22),
.B(n_177),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_25),
.B(n_32),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_25),
.B(n_124),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_25),
.A2(n_31),
.B(n_124),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_25),
.B(n_165),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_26),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_28),
.B(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_28),
.B(n_164),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_46),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_35),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_44),
.Y(n_35)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_36),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_36),
.B(n_47),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_43),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_37)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_38),
.A2(n_42),
.B1(n_78),
.B2(n_79),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_38),
.B(n_152),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_42),
.A2(n_45),
.B(n_79),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_43),
.B(n_139),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_44),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_45),
.A2(n_55),
.B(n_57),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_46),
.B(n_138),
.Y(n_157)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_69),
.C(n_74),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_49),
.A2(n_50),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_62),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_58),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_52),
.B(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_52)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_57),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_56),
.B1(n_59),
.B2(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_58),
.B(n_65),
.Y(n_99)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_69),
.A2(n_70),
.B1(n_74),
.B2(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_72),
.B(n_73),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_72),
.B(n_73),
.Y(n_136)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_82),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_81),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_76),
.B(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_76),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_80),
.B(n_81),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_83),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

INVxp67_ASAP7_75t_SL g92 ( 
.A(n_85),
.Y(n_92)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_102),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_96),
.B1(n_100),
.B2(n_101),
.Y(n_89)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_93),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_95),
.B(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_96),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_107),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_107),
.Y(n_117)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_109),
.B(n_171),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_117),
.C(n_118),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_112),
.A2(n_113),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_118),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_121),
.C(n_122),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_122),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_123),
.B(n_179),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_143),
.B(n_204),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_140),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_128),
.B(n_140),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.C(n_135),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_129),
.B(n_202),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_131),
.B(n_135),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_132),
.A2(n_134),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_132),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_134),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_199),
.B(n_203),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_186),
.B(n_198),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_168),
.B(n_185),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_153),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_147),
.B(n_153),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_150),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_148),
.A2(n_150),
.B1(n_151),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_160),
.B2(n_167),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_156),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_159),
.C(n_167),
.Y(n_187)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_157),
.Y(n_159)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_174),
.B(n_184),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_170),
.B(n_172),
.Y(n_184)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_180),
.B(n_183),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_181),
.B(n_182),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_187),
.B(n_188),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_195),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_193),
.C(n_195),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_200),
.B(n_201),
.Y(n_203)
);


endmodule