module fake_jpeg_2286_n_77 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_77);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_77;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_18),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_24),
.B(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_25),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_19),
.C(n_17),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_31),
.C(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_36),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_39),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_30),
.B1(n_29),
.B2(n_22),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_46),
.B1(n_33),
.B2(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_33),
.Y(n_50)
);

BUFx2_ASAP7_75t_SL g44 ( 
.A(n_38),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_44),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_30),
.B1(n_29),
.B2(n_32),
.Y(n_46)
);

AND2x6_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_10),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_47),
.B(n_21),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_48),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_52),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_23),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_51),
.B(n_27),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_45),
.Y(n_52)
);

OAI21x1_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_41),
.B(n_42),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_54),
.A2(n_3),
.B(n_4),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_55),
.B(n_57),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_41),
.B1(n_23),
.B2(n_21),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_60),
.B1(n_5),
.B2(n_6),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_32),
.C(n_41),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_58),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_SL g61 ( 
.A1(n_57),
.A2(n_59),
.B(n_60),
.C(n_53),
.Y(n_61)
);

NAND3xp33_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_62),
.C(n_63),
.Y(n_68)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_66),
.C(n_6),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_65),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_69),
.C(n_70),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

MAJx2_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_16),
.C(n_12),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_13),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_15),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_71),
.B(n_8),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_7),
.B(n_8),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_9),
.Y(n_77)
);


endmodule