module fake_netlist_6_1799_n_1736 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1736);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1736;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_93),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_34),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_150),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_157),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_26),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_37),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_127),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_2),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_101),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_81),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_77),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_122),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_94),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_91),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_39),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_78),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_38),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_41),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_9),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_15),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_7),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_118),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_5),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_66),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_71),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_125),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_126),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_44),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_44),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_80),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_30),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_36),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_9),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_39),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_69),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_123),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_165),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_129),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_11),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_121),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_70),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_149),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_144),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_26),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g214 ( 
.A(n_160),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_120),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_61),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_3),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_11),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_4),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_37),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_68),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_112),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_124),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_53),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_24),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_73),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_141),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_5),
.Y(n_228)
);

BUFx8_ASAP7_75t_SL g229 ( 
.A(n_50),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_97),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_25),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_86),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_4),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_131),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_90),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_41),
.Y(n_236)
);

BUFx10_ASAP7_75t_L g237 ( 
.A(n_48),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_103),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_85),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_153),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_48),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_46),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_18),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_65),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_58),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_13),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_107),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_33),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_75),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_158),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_117),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_27),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_156),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_47),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_146),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_147),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_163),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_30),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_99),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_32),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_16),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_19),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_98),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_15),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_47),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_46),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_82),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_22),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_132),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_138),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_2),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_10),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_74),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_43),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_106),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_7),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_51),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_12),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_19),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_111),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_109),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_67),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_24),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_22),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_0),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_20),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_96),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_135),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_143),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_28),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_100),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_34),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_84),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_83),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_6),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_64),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_17),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_28),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_63),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_152),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_134),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_31),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_50),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_116),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_57),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_56),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_137),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_55),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_53),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_108),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_62),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_29),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_0),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_42),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_29),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_89),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_27),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_17),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_76),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_36),
.Y(n_320)
);

BUFx10_ASAP7_75t_L g321 ( 
.A(n_54),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_159),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_115),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_133),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_3),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_52),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_164),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_148),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_79),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_155),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_202),
.Y(n_331)
);

NOR2xp67_ASAP7_75t_L g332 ( 
.A(n_297),
.B(n_1),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_203),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_167),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_167),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_229),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_172),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_172),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_168),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_269),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_202),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_171),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_288),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_190),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_322),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_190),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_192),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_186),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_166),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_186),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_186),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_186),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_327),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_189),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_238),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_192),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_256),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_178),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_193),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_193),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_194),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_237),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_194),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_291),
.B(n_1),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_196),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_291),
.B(n_6),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_205),
.B(n_8),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_205),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_197),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_210),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_169),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_210),
.B(n_8),
.Y(n_372)
);

NOR2xp67_ASAP7_75t_L g373 ( 
.A(n_297),
.B(n_10),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_186),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_223),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_237),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_223),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_232),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_199),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_227),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_227),
.B(n_12),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_170),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_201),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_239),
.Y(n_384)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_173),
.B(n_175),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_239),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_208),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_240),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_217),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_174),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_218),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_237),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_176),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_240),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_177),
.Y(n_395)
);

CKINVDCx14_ASAP7_75t_R g396 ( 
.A(n_321),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_249),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_219),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_180),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_321),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_224),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_259),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_233),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_236),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_182),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_249),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g407 ( 
.A(n_173),
.B(n_13),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_255),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_241),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_255),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_280),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_321),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_184),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_280),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_242),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_228),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_350),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_350),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_R g419 ( 
.A(n_358),
.B(n_195),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_348),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_333),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_340),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_371),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_351),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_351),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_402),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_352),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_343),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_352),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_382),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_345),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_390),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_348),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_374),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_393),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_378),
.B(n_232),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_402),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_339),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_374),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_416),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_395),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_399),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_353),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_416),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_405),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_402),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_339),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_402),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_402),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_385),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_385),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_413),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_336),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_334),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_335),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_355),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_357),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_336),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_337),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_338),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_344),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_349),
.B(n_287),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_342),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_396),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_346),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_364),
.B(n_287),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_347),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_342),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_365),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_356),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_362),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_359),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_366),
.B(n_282),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_360),
.B(n_282),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_361),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_363),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_365),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_368),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_369),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_369),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_376),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_370),
.B(n_179),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_375),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_379),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_379),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_377),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_380),
.Y(n_487)
);

CKINVDCx8_ASAP7_75t_R g488 ( 
.A(n_400),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_384),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_386),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_388),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_383),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_394),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_466),
.A2(n_367),
.B1(n_372),
.B2(n_381),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_473),
.B(n_397),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_436),
.B(n_406),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_L g497 ( 
.A1(n_462),
.A2(n_341),
.B1(n_331),
.B2(n_407),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_474),
.B(n_179),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_474),
.B(n_181),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_459),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_450),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_420),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_487),
.Y(n_503)
);

NAND3xp33_ASAP7_75t_L g504 ( 
.A(n_450),
.B(n_354),
.C(n_383),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_451),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_451),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_474),
.B(n_181),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_419),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_420),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_474),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_459),
.Y(n_511)
);

BUFx10_ASAP7_75t_L g512 ( 
.A(n_453),
.Y(n_512)
);

BUFx4f_ASAP7_75t_L g513 ( 
.A(n_487),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_465),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_433),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_490),
.B(n_204),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_465),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_490),
.B(n_408),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_438),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_433),
.Y(n_520)
);

INVx5_ASAP7_75t_L g521 ( 
.A(n_446),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_470),
.B(n_410),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_470),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_463),
.B(n_387),
.Y(n_524)
);

INVx4_ASAP7_75t_SL g525 ( 
.A(n_446),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_472),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_454),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_490),
.B(n_411),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_439),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_479),
.Y(n_530)
);

NAND3xp33_ASAP7_75t_L g531 ( 
.A(n_447),
.B(n_389),
.C(n_387),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_490),
.B(n_414),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_454),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_472),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_468),
.B(n_389),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_439),
.Y(n_536)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_487),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_475),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_475),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_446),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_478),
.B(n_391),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_469),
.B(n_391),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_449),
.B(n_398),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_446),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_454),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_449),
.B(n_398),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_482),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_482),
.A2(n_478),
.B1(n_491),
.B2(n_483),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_454),
.B(n_401),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_417),
.Y(n_550)
);

NAND2x1p5_ASAP7_75t_L g551 ( 
.A(n_482),
.B(n_296),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_454),
.B(n_401),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_483),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_489),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_491),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_477),
.B(n_403),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_446),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_447),
.B(n_392),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_493),
.Y(n_559)
);

BUFx8_ASAP7_75t_SL g560 ( 
.A(n_471),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_482),
.B(n_204),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_417),
.Y(n_562)
);

INVx6_ASAP7_75t_L g563 ( 
.A(n_489),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_487),
.B(n_245),
.Y(n_564)
);

OAI22xp33_ASAP7_75t_L g565 ( 
.A1(n_480),
.A2(n_313),
.B1(n_407),
.B2(n_373),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_487),
.B(n_245),
.Y(n_566)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_421),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_484),
.B(n_403),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_493),
.Y(n_569)
);

AND3x2_ASAP7_75t_L g570 ( 
.A(n_480),
.B(n_294),
.C(n_263),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_485),
.A2(n_415),
.B1(n_409),
.B2(n_404),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_455),
.B(n_296),
.Y(n_572)
);

OAI22xp33_ASAP7_75t_L g573 ( 
.A1(n_492),
.A2(n_332),
.B1(n_243),
.B2(n_277),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_489),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_422),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_455),
.B(n_404),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_489),
.Y(n_577)
);

OR2x2_ASAP7_75t_L g578 ( 
.A(n_481),
.B(n_412),
.Y(n_578)
);

NAND2xp33_ASAP7_75t_R g579 ( 
.A(n_423),
.B(n_409),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_440),
.B(n_444),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_426),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_489),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_460),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_460),
.B(n_415),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_487),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_426),
.B(n_198),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_426),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_461),
.A2(n_272),
.B1(n_228),
.B2(n_283),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_461),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_426),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_430),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_437),
.B(n_206),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_467),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_418),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_437),
.B(n_207),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_437),
.B(n_209),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_437),
.B(n_211),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_464),
.A2(n_251),
.B1(n_329),
.B2(n_324),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_467),
.B(n_246),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_476),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_476),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_432),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_486),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_L g604 ( 
.A(n_486),
.B(n_259),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_418),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_424),
.B(n_263),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_456),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_440),
.B(n_258),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_424),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_448),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g611 ( 
.A(n_481),
.B(n_225),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_425),
.B(n_294),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_425),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_444),
.B(n_427),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_448),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_429),
.A2(n_283),
.B1(n_272),
.B2(n_292),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_429),
.Y(n_617)
);

OAI22xp33_ASAP7_75t_L g618 ( 
.A1(n_488),
.A2(n_278),
.B1(n_261),
.B2(n_274),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_434),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_434),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_458),
.B(n_284),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_488),
.B(n_225),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_428),
.Y(n_623)
);

AND2x6_ASAP7_75t_L g624 ( 
.A(n_435),
.B(n_299),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_441),
.Y(n_625)
);

INVx6_ASAP7_75t_L g626 ( 
.A(n_442),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_445),
.B(n_252),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_452),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_457),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_431),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_443),
.Y(n_631)
);

AND2x6_ASAP7_75t_L g632 ( 
.A(n_466),
.B(n_299),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_466),
.B(n_212),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_466),
.B(n_252),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_474),
.B(n_300),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_466),
.B(n_215),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_466),
.B(n_325),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_420),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_459),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_459),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_466),
.B(n_325),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_459),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_459),
.Y(n_643)
);

INVx4_ASAP7_75t_L g644 ( 
.A(n_487),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_459),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g646 ( 
.A(n_611),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_494),
.B(n_547),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_550),
.Y(n_648)
);

O2A1O1Ixp33_ASAP7_75t_L g649 ( 
.A1(n_501),
.A2(n_264),
.B(n_292),
.C(n_326),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_501),
.B(n_286),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_541),
.B(n_183),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_580),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_632),
.B(n_300),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_504),
.B(n_298),
.Y(n_654)
);

INVx4_ASAP7_75t_L g655 ( 
.A(n_510),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_510),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_632),
.B(n_305),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_632),
.B(n_305),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_632),
.B(n_306),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_627),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_547),
.A2(n_330),
.B1(n_328),
.B2(n_323),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_632),
.B(n_306),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_541),
.B(n_530),
.Y(n_663)
);

INVxp67_ASAP7_75t_L g664 ( 
.A(n_558),
.Y(n_664)
);

NOR2xp67_ASAP7_75t_L g665 ( 
.A(n_508),
.B(n_221),
.Y(n_665)
);

NAND2x1_ASAP7_75t_L g666 ( 
.A(n_563),
.B(n_259),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_562),
.Y(n_667)
);

INVx1_ASAP7_75t_SL g668 ( 
.A(n_558),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_549),
.B(n_259),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_L g670 ( 
.A(n_624),
.B(n_222),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_495),
.B(n_319),
.Y(n_671)
);

NOR2xp67_ASAP7_75t_L g672 ( 
.A(n_508),
.B(n_226),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_580),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_505),
.B(n_302),
.Y(n_674)
);

BUFx8_ASAP7_75t_L g675 ( 
.A(n_607),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_633),
.B(n_319),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_552),
.B(n_259),
.Y(n_677)
);

NOR2xp67_ASAP7_75t_L g678 ( 
.A(n_531),
.B(n_230),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_636),
.B(n_496),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_594),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_627),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_594),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_635),
.B(n_216),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_530),
.B(n_185),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_500),
.Y(n_685)
);

INVxp67_ASAP7_75t_SL g686 ( 
.A(n_582),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_620),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_605),
.B(n_323),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_506),
.B(n_309),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_620),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_502),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_605),
.B(n_328),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_634),
.B(n_254),
.Y(n_693)
);

INVx8_ASAP7_75t_L g694 ( 
.A(n_624),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_513),
.A2(n_270),
.B(n_273),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_576),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_584),
.B(n_314),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_502),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_543),
.B(n_317),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_583),
.B(n_234),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_624),
.A2(n_275),
.B1(n_316),
.B2(n_235),
.Y(n_701)
);

INVx8_ASAP7_75t_L g702 ( 
.A(n_624),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_635),
.B(n_244),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_635),
.B(n_247),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_634),
.B(n_312),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_583),
.B(n_250),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_617),
.B(n_253),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_611),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_593),
.B(n_617),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_593),
.B(n_257),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_546),
.B(n_267),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_619),
.B(n_281),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_509),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_565),
.B(n_289),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_619),
.B(n_293),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_622),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_609),
.B(n_301),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_622),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_SL g719 ( 
.A(n_512),
.B(n_318),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_511),
.B(n_175),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_514),
.B(n_307),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_517),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_637),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_637),
.B(n_214),
.Y(n_724)
);

OAI21xp5_ASAP7_75t_L g725 ( 
.A1(n_498),
.A2(n_311),
.B(n_310),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_641),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_641),
.B(n_214),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_519),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_523),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_613),
.B(n_264),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_526),
.B(n_220),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_534),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_538),
.B(n_271),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_539),
.B(n_276),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_553),
.B(n_326),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_555),
.B(n_187),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_559),
.Y(n_737)
);

NAND3xp33_ASAP7_75t_L g738 ( 
.A(n_497),
.B(n_320),
.C(n_315),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_569),
.B(n_187),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_639),
.B(n_214),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_640),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_642),
.Y(n_742)
);

AO221x1_ASAP7_75t_L g743 ( 
.A1(n_573),
.A2(n_320),
.B1(n_315),
.B2(n_308),
.C(n_188),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_572),
.A2(n_308),
.B1(n_188),
.B2(n_303),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_579),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_509),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_643),
.B(n_265),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_645),
.B(n_304),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_610),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_614),
.B(n_265),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_522),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_581),
.B(n_304),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_581),
.B(n_304),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_589),
.B(n_303),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_515),
.Y(n_755)
);

INVxp33_ASAP7_75t_L g756 ( 
.A(n_560),
.Y(n_756)
);

INVxp67_ASAP7_75t_L g757 ( 
.A(n_621),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_515),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_600),
.B(n_295),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_601),
.B(n_295),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_513),
.A2(n_290),
.B(n_285),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_603),
.B(n_290),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_522),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_571),
.B(n_285),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_524),
.B(n_535),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_615),
.B(n_279),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_610),
.Y(n_767)
);

NAND2xp33_ASAP7_75t_L g768 ( 
.A(n_624),
.B(n_268),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_570),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_615),
.B(n_268),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_498),
.B(n_266),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_542),
.B(n_266),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_499),
.B(n_262),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_499),
.B(n_262),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_610),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_507),
.B(n_260),
.Y(n_776)
);

NOR2x1p5_ASAP7_75t_L g777 ( 
.A(n_578),
.B(n_260),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_556),
.B(n_248),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_561),
.A2(n_248),
.B1(n_231),
.B2(n_213),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_520),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_568),
.B(n_231),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_507),
.B(n_213),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_548),
.A2(n_200),
.B1(n_191),
.B2(n_60),
.Y(n_783)
);

A2O1A1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_608),
.A2(n_528),
.B(n_532),
.C(n_518),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_581),
.B(n_200),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_599),
.B(n_191),
.Y(n_786)
);

O2A1O1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_561),
.A2(n_14),
.B(n_16),
.C(n_18),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_590),
.B(n_59),
.Y(n_788)
);

BUFx6f_ASAP7_75t_SL g789 ( 
.A(n_512),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_590),
.B(n_72),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_628),
.B(n_14),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_520),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_618),
.B(n_598),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_638),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_567),
.Y(n_795)
);

NAND2xp33_ASAP7_75t_L g796 ( 
.A(n_610),
.B(n_87),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_590),
.B(n_162),
.Y(n_797)
);

O2A1O1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_606),
.A2(n_20),
.B(n_21),
.C(n_23),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_527),
.B(n_154),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_SL g800 ( 
.A(n_512),
.B(n_21),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_628),
.B(n_23),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_586),
.A2(n_88),
.B1(n_142),
.B2(n_139),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_533),
.B(n_151),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_626),
.Y(n_804)
);

AO21x1_ASAP7_75t_L g805 ( 
.A1(n_653),
.A2(n_551),
.B(n_566),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_679),
.B(n_551),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_696),
.B(n_533),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_697),
.B(n_772),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_691),
.Y(n_809)
);

NOR2x1_ASAP7_75t_L g810 ( 
.A(n_804),
.B(n_625),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_765),
.B(n_623),
.Y(n_811)
);

AND2x4_ASAP7_75t_L g812 ( 
.A(n_804),
.B(n_630),
.Y(n_812)
);

OAI21xp5_ASAP7_75t_L g813 ( 
.A1(n_647),
.A2(n_516),
.B(n_585),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_709),
.A2(n_513),
.B(n_503),
.Y(n_814)
);

NAND2xp33_ASAP7_75t_L g815 ( 
.A(n_694),
.B(n_587),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_648),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_697),
.B(n_545),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_691),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_765),
.B(n_630),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_793),
.A2(n_616),
.B1(n_588),
.B2(n_578),
.Y(n_820)
);

A2O1A1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_793),
.A2(n_595),
.B(n_597),
.C(n_592),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_784),
.A2(n_644),
.B(n_537),
.Y(n_822)
);

A2O1A1Ixp33_ASAP7_75t_L g823 ( 
.A1(n_772),
.A2(n_596),
.B(n_516),
.C(n_574),
.Y(n_823)
);

O2A1O1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_647),
.A2(n_612),
.B(n_606),
.C(n_566),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_764),
.A2(n_577),
.B1(n_564),
.B2(n_536),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_663),
.B(n_591),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_716),
.A2(n_545),
.B1(n_554),
.B2(n_563),
.Y(n_827)
);

NOR2x1p5_ASAP7_75t_L g828 ( 
.A(n_745),
.B(n_629),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_L g829 ( 
.A1(n_744),
.A2(n_626),
.B1(n_631),
.B2(n_602),
.Y(n_829)
);

NAND3xp33_ASAP7_75t_L g830 ( 
.A(n_778),
.B(n_612),
.C(n_564),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_768),
.A2(n_644),
.B(n_537),
.Y(n_831)
);

INVxp67_ASAP7_75t_L g832 ( 
.A(n_646),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_652),
.B(n_554),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_728),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_655),
.Y(n_835)
);

BUFx2_ASAP7_75t_L g836 ( 
.A(n_795),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_712),
.A2(n_503),
.B(n_540),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_778),
.B(n_544),
.Y(n_838)
);

O2A1O1Ixp33_ASAP7_75t_SL g839 ( 
.A1(n_790),
.A2(n_529),
.B(n_536),
.C(n_638),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_718),
.B(n_587),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_757),
.B(n_626),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_723),
.B(n_587),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_668),
.B(n_626),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_781),
.B(n_711),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_698),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_789),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_781),
.B(n_544),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_670),
.A2(n_557),
.B(n_540),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_664),
.B(n_575),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_698),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_648),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_655),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_656),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_711),
.B(n_544),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_699),
.B(n_587),
.Y(n_855)
);

NAND3xp33_ASAP7_75t_L g856 ( 
.A(n_714),
.B(n_575),
.C(n_604),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_675),
.Y(n_857)
);

O2A1O1Ixp33_ASAP7_75t_SL g858 ( 
.A1(n_790),
.A2(n_604),
.B(n_563),
.C(n_525),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_656),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_673),
.B(n_525),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_650),
.B(n_557),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_713),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_650),
.B(n_521),
.Y(n_863)
);

NOR2x1_ASAP7_75t_L g864 ( 
.A(n_665),
.B(n_560),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_708),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_L g866 ( 
.A1(n_744),
.A2(n_521),
.B1(n_31),
.B2(n_32),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_726),
.B(n_521),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_676),
.B(n_25),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_749),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_660),
.B(n_33),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_749),
.A2(n_92),
.B(n_130),
.Y(n_871)
);

A2O1A1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_764),
.A2(n_35),
.B(n_38),
.C(n_40),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_751),
.B(n_110),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_749),
.A2(n_136),
.B(n_128),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_763),
.B(n_35),
.Y(n_875)
);

NAND3xp33_ASAP7_75t_L g876 ( 
.A(n_714),
.B(n_40),
.C(n_42),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_681),
.B(n_43),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_749),
.A2(n_767),
.B(n_775),
.Y(n_878)
);

AO21x1_ASAP7_75t_L g879 ( 
.A1(n_657),
.A2(n_45),
.B(n_49),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_767),
.A2(n_95),
.B(n_114),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_685),
.B(n_45),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_713),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_791),
.B(n_119),
.Y(n_883)
);

AOI22x1_ASAP7_75t_L g884 ( 
.A1(n_667),
.A2(n_105),
.B1(n_104),
.B2(n_102),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_693),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_684),
.B(n_49),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_722),
.B(n_51),
.Y(n_887)
);

BUFx3_ASAP7_75t_L g888 ( 
.A(n_675),
.Y(n_888)
);

NAND2x1p5_ASAP7_75t_L g889 ( 
.A(n_767),
.B(n_52),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_746),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_775),
.Y(n_891)
);

A2O1A1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_654),
.A2(n_54),
.B(n_55),
.C(n_674),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_707),
.A2(n_715),
.B1(n_737),
.B2(n_742),
.Y(n_893)
);

NOR2x1_ASAP7_75t_L g894 ( 
.A(n_672),
.B(n_678),
.Y(n_894)
);

INVx3_ASAP7_75t_L g895 ( 
.A(n_775),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_746),
.Y(n_896)
);

BUFx4f_ASAP7_75t_L g897 ( 
.A(n_801),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_651),
.B(n_654),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_729),
.B(n_732),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_705),
.Y(n_900)
);

A2O1A1Ixp33_ASAP7_75t_L g901 ( 
.A1(n_674),
.A2(n_689),
.B(n_786),
.C(n_659),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_741),
.B(n_724),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_SL g903 ( 
.A1(n_719),
.A2(n_800),
.B1(n_727),
.B2(n_702),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_686),
.B(n_671),
.Y(n_904)
);

AND2x2_ASAP7_75t_SL g905 ( 
.A(n_779),
.B(n_689),
.Y(n_905)
);

AOI21xp33_ASAP7_75t_L g906 ( 
.A1(n_783),
.A2(n_662),
.B(n_658),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_688),
.B(n_692),
.Y(n_907)
);

AND2x6_ASAP7_75t_L g908 ( 
.A(n_802),
.B(n_720),
.Y(n_908)
);

OAI21xp5_ASAP7_75t_L g909 ( 
.A1(n_785),
.A2(n_680),
.B(n_690),
.Y(n_909)
);

BUFx4f_ASAP7_75t_L g910 ( 
.A(n_769),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_775),
.A2(n_669),
.B(n_677),
.Y(n_911)
);

AOI21x1_ASAP7_75t_L g912 ( 
.A1(n_677),
.A2(n_707),
.B(n_715),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_721),
.A2(n_683),
.B1(n_753),
.B2(n_752),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_694),
.A2(n_702),
.B(n_710),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_779),
.A2(n_750),
.B1(n_738),
.B2(n_774),
.Y(n_915)
);

NAND3xp33_ASAP7_75t_SL g916 ( 
.A(n_740),
.B(n_748),
.C(n_787),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_680),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_720),
.B(n_777),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_694),
.A2(n_702),
.B(n_706),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_720),
.Y(n_920)
);

AOI21xp33_ASAP7_75t_L g921 ( 
.A1(n_725),
.A2(n_717),
.B(n_703),
.Y(n_921)
);

OAI21xp33_ASAP7_75t_L g922 ( 
.A1(n_731),
.A2(n_734),
.B(n_733),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_740),
.B(n_748),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_700),
.A2(n_803),
.B(n_799),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_771),
.A2(n_776),
.B1(n_773),
.B2(n_782),
.Y(n_925)
);

BUFx8_ASAP7_75t_SL g926 ( 
.A(n_789),
.Y(n_926)
);

NOR2xp67_ASAP7_75t_L g927 ( 
.A(n_701),
.B(n_770),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_788),
.A2(n_797),
.B(n_682),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_687),
.B(n_766),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_703),
.A2(n_704),
.B(n_683),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_785),
.A2(n_755),
.B(n_758),
.Y(n_931)
);

AND2x6_ASAP7_75t_L g932 ( 
.A(n_755),
.B(n_758),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_735),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_780),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_780),
.Y(n_935)
);

AOI22xp33_ASAP7_75t_L g936 ( 
.A1(n_743),
.A2(n_661),
.B1(n_794),
.B2(n_792),
.Y(n_936)
);

OAI21x1_ASAP7_75t_L g937 ( 
.A1(n_792),
.A2(n_794),
.B(n_666),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_761),
.A2(n_730),
.B(n_747),
.Y(n_938)
);

NOR2xp67_ASAP7_75t_L g939 ( 
.A(n_736),
.B(n_739),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_704),
.A2(n_721),
.B(n_753),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_754),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_752),
.B(n_760),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_759),
.B(n_762),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_756),
.B(n_798),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_649),
.A2(n_695),
.B(n_796),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_647),
.A2(n_784),
.B(n_679),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_709),
.A2(n_513),
.B(n_679),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_697),
.A2(n_793),
.B(n_778),
.C(n_781),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_709),
.A2(n_513),
.B(n_679),
.Y(n_949)
);

AND2x2_ASAP7_75t_SL g950 ( 
.A(n_719),
.B(n_800),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_648),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_691),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_709),
.A2(n_513),
.B(n_679),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_709),
.A2(n_513),
.B(n_679),
.Y(n_954)
);

OR2x2_ASAP7_75t_L g955 ( 
.A(n_668),
.B(n_664),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_663),
.B(n_696),
.Y(n_956)
);

NOR3xp33_ASAP7_75t_L g957 ( 
.A(n_765),
.B(n_531),
.C(n_793),
.Y(n_957)
);

O2A1O1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_647),
.A2(n_772),
.B(n_781),
.C(n_778),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_793),
.A2(n_647),
.B1(n_679),
.B2(n_697),
.Y(n_959)
);

OAI21xp33_ASAP7_75t_SL g960 ( 
.A1(n_647),
.A2(n_679),
.B(n_673),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_793),
.A2(n_494),
.B1(n_744),
.B2(n_679),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_793),
.A2(n_494),
.B1(n_744),
.B2(n_679),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_663),
.B(n_696),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_663),
.B(n_696),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_L g965 ( 
.A1(n_647),
.A2(n_784),
.B(n_679),
.Y(n_965)
);

AOI22xp5_ASAP7_75t_L g966 ( 
.A1(n_793),
.A2(n_647),
.B1(n_679),
.B2(n_697),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_679),
.B(n_696),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_793),
.A2(n_494),
.B1(n_744),
.B2(n_679),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_709),
.A2(n_513),
.B(n_679),
.Y(n_969)
);

AO21x2_ASAP7_75t_L g970 ( 
.A1(n_653),
.A2(n_658),
.B(n_657),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_691),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_663),
.B(n_696),
.Y(n_972)
);

AND2x6_ASAP7_75t_L g973 ( 
.A(n_652),
.B(n_673),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_745),
.Y(n_974)
);

INVx1_ASAP7_75t_SL g975 ( 
.A(n_668),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_679),
.B(n_696),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_647),
.A2(n_772),
.B(n_781),
.C(n_778),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_663),
.B(n_696),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_795),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_806),
.A2(n_855),
.B(n_947),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_860),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_816),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_808),
.B(n_959),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_949),
.A2(n_954),
.B(n_953),
.Y(n_984)
);

AO31x2_ASAP7_75t_L g985 ( 
.A1(n_805),
.A2(n_948),
.A3(n_823),
.B(n_901),
.Y(n_985)
);

NOR2x1_ASAP7_75t_L g986 ( 
.A(n_841),
.B(n_843),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_946),
.A2(n_965),
.B(n_966),
.Y(n_987)
);

AO31x2_ASAP7_75t_L g988 ( 
.A1(n_879),
.A2(n_822),
.A3(n_821),
.B(n_844),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_972),
.B(n_978),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_809),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_946),
.A2(n_965),
.B(n_960),
.Y(n_991)
);

NOR2xp67_ASAP7_75t_SL g992 ( 
.A(n_835),
.B(n_852),
.Y(n_992)
);

INVx2_ASAP7_75t_SL g993 ( 
.A(n_836),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_958),
.A2(n_977),
.B(n_898),
.C(n_961),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_961),
.A2(n_968),
.B1(n_962),
.B2(n_905),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_962),
.A2(n_968),
.B(n_892),
.C(n_967),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_976),
.B(n_819),
.Y(n_997)
);

AO31x2_ASAP7_75t_L g998 ( 
.A1(n_969),
.A2(n_928),
.A3(n_861),
.B(n_930),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_851),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_957),
.A2(n_940),
.B(n_921),
.C(n_913),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_831),
.A2(n_815),
.B(n_924),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_854),
.A2(n_907),
.B(n_817),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_941),
.B(n_904),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_818),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_979),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_897),
.B(n_950),
.Y(n_1006)
);

OR2x2_ASAP7_75t_L g1007 ( 
.A(n_975),
.B(n_955),
.Y(n_1007)
);

OAI22x1_ASAP7_75t_L g1008 ( 
.A1(n_811),
.A2(n_886),
.B1(n_944),
.B2(n_975),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_845),
.Y(n_1009)
);

AO31x2_ASAP7_75t_L g1010 ( 
.A1(n_915),
.A2(n_911),
.A3(n_848),
.B(n_838),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_933),
.B(n_902),
.Y(n_1011)
);

AOI21x1_ASAP7_75t_L g1012 ( 
.A1(n_863),
.A2(n_912),
.B(n_927),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_837),
.A2(n_906),
.B(n_929),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_850),
.Y(n_1014)
);

O2A1O1Ixp5_ASAP7_75t_L g1015 ( 
.A1(n_945),
.A2(n_938),
.B(n_906),
.C(n_868),
.Y(n_1015)
);

AOI21xp33_ASAP7_75t_L g1016 ( 
.A1(n_915),
.A2(n_820),
.B(n_824),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_814),
.A2(n_919),
.B(n_914),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_813),
.A2(n_830),
.B(n_909),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_939),
.B(n_847),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_813),
.A2(n_931),
.B(n_925),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_812),
.B(n_918),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_970),
.A2(n_878),
.B(n_938),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_832),
.B(n_956),
.Y(n_1023)
);

INVxp67_ASAP7_75t_L g1024 ( 
.A(n_826),
.Y(n_1024)
);

OR2x2_ASAP7_75t_L g1025 ( 
.A(n_885),
.B(n_900),
.Y(n_1025)
);

BUFx12f_ASAP7_75t_L g1026 ( 
.A(n_846),
.Y(n_1026)
);

OAI21x1_ASAP7_75t_L g1027 ( 
.A1(n_917),
.A2(n_951),
.B(n_934),
.Y(n_1027)
);

NAND3xp33_ASAP7_75t_L g1028 ( 
.A(n_849),
.B(n_903),
.C(n_829),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_922),
.B(n_925),
.Y(n_1029)
);

OAI22x1_ASAP7_75t_L g1030 ( 
.A1(n_828),
.A2(n_876),
.B1(n_923),
.B2(n_918),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_893),
.B(n_942),
.Y(n_1031)
);

INVxp67_ASAP7_75t_L g1032 ( 
.A(n_834),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_865),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_891),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_812),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_899),
.B(n_807),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_970),
.A2(n_943),
.B(n_859),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_945),
.A2(n_858),
.B(n_897),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_973),
.B(n_935),
.Y(n_1039)
);

NAND3xp33_ASAP7_75t_SL g1040 ( 
.A(n_974),
.B(n_829),
.C(n_872),
.Y(n_1040)
);

OA21x2_ASAP7_75t_L g1041 ( 
.A1(n_936),
.A2(n_825),
.B(n_896),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_973),
.B(n_971),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_862),
.A2(n_882),
.B(n_890),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_952),
.Y(n_1044)
);

NOR2x1_ASAP7_75t_L g1045 ( 
.A(n_864),
.B(n_894),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_973),
.B(n_820),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_867),
.A2(n_839),
.B(n_883),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_963),
.B(n_964),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_842),
.A2(n_840),
.B(n_891),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_916),
.A2(n_856),
.B(n_877),
.C(n_870),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_973),
.B(n_873),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_873),
.B(n_833),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_810),
.B(n_920),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_889),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_869),
.A2(n_895),
.B(n_827),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_835),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_908),
.B(n_920),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_SL g1058 ( 
.A1(n_866),
.A2(n_875),
.B(n_881),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_908),
.B(n_895),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_887),
.B(n_910),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_908),
.A2(n_932),
.B(n_866),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_932),
.B(n_860),
.Y(n_1062)
);

AOI21xp33_ASAP7_75t_L g1063 ( 
.A1(n_884),
.A2(n_852),
.B(n_853),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_910),
.A2(n_880),
.B(n_874),
.C(n_871),
.Y(n_1064)
);

AO21x1_ASAP7_75t_L g1065 ( 
.A1(n_889),
.A2(n_932),
.B(n_853),
.Y(n_1065)
);

OR2x2_ASAP7_75t_L g1066 ( 
.A(n_857),
.B(n_888),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_852),
.B(n_853),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_926),
.B(n_808),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_948),
.A2(n_808),
.B(n_844),
.C(n_958),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_SL g1070 ( 
.A1(n_948),
.A2(n_965),
.B(n_946),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_972),
.B(n_663),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_972),
.B(n_663),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_972),
.B(n_663),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_972),
.B(n_663),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_836),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_808),
.B(n_959),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_808),
.B(n_959),
.Y(n_1077)
);

OR2x6_ASAP7_75t_L g1078 ( 
.A(n_836),
.B(n_626),
.Y(n_1078)
);

AOI221xp5_ASAP7_75t_L g1079 ( 
.A1(n_961),
.A2(n_962),
.B1(n_968),
.B2(n_764),
.C(n_948),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_809),
.Y(n_1080)
);

AO31x2_ASAP7_75t_L g1081 ( 
.A1(n_805),
.A2(n_948),
.A3(n_823),
.B(n_901),
.Y(n_1081)
);

AOI221xp5_ASAP7_75t_SL g1082 ( 
.A1(n_948),
.A2(n_977),
.B1(n_958),
.B2(n_961),
.C(n_968),
.Y(n_1082)
);

INVx5_ASAP7_75t_L g1083 ( 
.A(n_891),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_812),
.B(n_804),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_948),
.A2(n_808),
.B(n_844),
.C(n_958),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_809),
.Y(n_1086)
);

AOI21xp33_ASAP7_75t_L g1087 ( 
.A1(n_808),
.A2(n_844),
.B(n_948),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_812),
.B(n_804),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_948),
.A2(n_965),
.B(n_946),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_816),
.Y(n_1090)
);

AOI21x1_ASAP7_75t_L g1091 ( 
.A1(n_863),
.A2(n_861),
.B(n_822),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_808),
.B(n_811),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_959),
.B(n_966),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_937),
.A2(n_822),
.B(n_848),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_860),
.Y(n_1095)
);

INVx5_ASAP7_75t_L g1096 ( 
.A(n_891),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_SL g1097 ( 
.A1(n_930),
.A2(n_940),
.B(n_946),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_948),
.A2(n_808),
.B1(n_844),
.B2(n_959),
.Y(n_1098)
);

INVx2_ASAP7_75t_SL g1099 ( 
.A(n_836),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_809),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_948),
.A2(n_808),
.B(n_844),
.C(n_958),
.Y(n_1101)
);

AO21x2_ASAP7_75t_L g1102 ( 
.A1(n_948),
.A2(n_965),
.B(n_946),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_812),
.B(n_804),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_972),
.B(n_663),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_948),
.A2(n_965),
.B(n_946),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_975),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_860),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_959),
.B(n_966),
.Y(n_1108)
);

INVx3_ASAP7_75t_SL g1109 ( 
.A(n_846),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_808),
.B(n_844),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_959),
.B(n_966),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_937),
.A2(n_822),
.B(n_848),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_816),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1092),
.B(n_997),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1001),
.A2(n_1002),
.B(n_980),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_1098),
.B(n_983),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_997),
.B(n_1110),
.Y(n_1117)
);

BUFx4f_ASAP7_75t_L g1118 ( 
.A(n_1026),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_1083),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_1005),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_1028),
.B(n_983),
.Y(n_1121)
);

OR2x2_ASAP7_75t_L g1122 ( 
.A(n_1007),
.B(n_1025),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_1109),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_989),
.B(n_1071),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_1106),
.Y(n_1125)
);

INVx1_ASAP7_75t_SL g1126 ( 
.A(n_1075),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_982),
.Y(n_1127)
);

AND2x6_ASAP7_75t_L g1128 ( 
.A(n_1046),
.B(n_1051),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_1079),
.A2(n_995),
.B1(n_1098),
.B2(n_1108),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1003),
.B(n_1076),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_SL g1131 ( 
.A1(n_995),
.A2(n_1061),
.B1(n_1076),
.B2(n_1077),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_999),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1003),
.B(n_1077),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_SL g1134 ( 
.A1(n_1061),
.A2(n_1089),
.B1(n_1105),
.B2(n_987),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_1033),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_1056),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1072),
.B(n_1073),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1074),
.B(n_1104),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1036),
.B(n_1011),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_993),
.Y(n_1140)
);

CKINVDCx6p67_ASAP7_75t_R g1141 ( 
.A(n_1078),
.Y(n_1141)
);

INVx5_ASAP7_75t_L g1142 ( 
.A(n_1034),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1024),
.B(n_1035),
.Y(n_1143)
);

INVx3_ASAP7_75t_SL g1144 ( 
.A(n_1078),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1021),
.B(n_1084),
.Y(n_1145)
);

AOI222xp33_ASAP7_75t_L g1146 ( 
.A1(n_1093),
.A2(n_1111),
.B1(n_1040),
.B2(n_1008),
.C1(n_1105),
.C2(n_1089),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1069),
.A2(n_1101),
.B1(n_1085),
.B2(n_994),
.Y(n_1147)
);

BUFx12f_ASAP7_75t_L g1148 ( 
.A(n_1078),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1090),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1036),
.B(n_986),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1113),
.Y(n_1151)
);

AND2x2_ASAP7_75t_SL g1152 ( 
.A(n_1029),
.B(n_1046),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_1099),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_1056),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1087),
.B(n_1006),
.Y(n_1155)
);

CKINVDCx8_ASAP7_75t_R g1156 ( 
.A(n_1084),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_1068),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1087),
.A2(n_1000),
.B(n_1015),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1048),
.B(n_1031),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_1032),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1031),
.B(n_1060),
.Y(n_1161)
);

A2O1A1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_996),
.A2(n_1016),
.B(n_987),
.C(n_1082),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1102),
.A2(n_1058),
.B1(n_991),
.B2(n_1020),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_1068),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1027),
.Y(n_1165)
);

INVx2_ASAP7_75t_SL g1166 ( 
.A(n_1066),
.Y(n_1166)
);

NAND2xp33_ASAP7_75t_L g1167 ( 
.A(n_1050),
.B(n_1052),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1088),
.B(n_1103),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_1054),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1088),
.B(n_1103),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_1067),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_1052),
.B(n_1053),
.Y(n_1172)
);

NAND2xp33_ASAP7_75t_L g1173 ( 
.A(n_1051),
.B(n_1057),
.Y(n_1173)
);

INVxp67_ASAP7_75t_L g1174 ( 
.A(n_1023),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_1034),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_1053),
.B(n_981),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1030),
.B(n_981),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1038),
.A2(n_1082),
.B(n_1018),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1102),
.A2(n_1018),
.B1(n_1097),
.B2(n_1019),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1019),
.A2(n_1057),
.B1(n_1044),
.B2(n_1100),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1013),
.A2(n_1070),
.B(n_1022),
.Y(n_1181)
);

INVx1_ASAP7_75t_SL g1182 ( 
.A(n_1045),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_990),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_1083),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1043),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1095),
.B(n_1107),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1004),
.B(n_1086),
.Y(n_1187)
);

INVx1_ASAP7_75t_SL g1188 ( 
.A(n_1059),
.Y(n_1188)
);

AOI221x1_ASAP7_75t_L g1189 ( 
.A1(n_984),
.A2(n_1037),
.B1(n_1047),
.B2(n_1017),
.C(n_1064),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_1083),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1009),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1083),
.Y(n_1192)
);

OAI21xp33_ASAP7_75t_L g1193 ( 
.A1(n_1039),
.A2(n_1014),
.B(n_1080),
.Y(n_1193)
);

AOI21xp33_ASAP7_75t_SL g1194 ( 
.A1(n_1063),
.A2(n_1062),
.B(n_1039),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_992),
.B(n_988),
.Y(n_1195)
);

OR2x6_ASAP7_75t_SL g1196 ( 
.A(n_1042),
.B(n_1065),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1041),
.A2(n_1042),
.B1(n_1063),
.B2(n_1049),
.Y(n_1197)
);

O2A1O1Ixp33_ASAP7_75t_SL g1198 ( 
.A1(n_985),
.A2(n_1081),
.B(n_988),
.C(n_1055),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_1096),
.Y(n_1199)
);

AO31x2_ASAP7_75t_L g1200 ( 
.A1(n_985),
.A2(n_1081),
.A3(n_988),
.B(n_1010),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_1010),
.B(n_985),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1010),
.B(n_1081),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_1091),
.B(n_1012),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_998),
.B(n_1094),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_998),
.B(n_1112),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_998),
.Y(n_1206)
);

OR2x2_ASAP7_75t_L g1207 ( 
.A(n_997),
.B(n_1007),
.Y(n_1207)
);

INVx4_ASAP7_75t_L g1208 ( 
.A(n_1056),
.Y(n_1208)
);

CKINVDCx11_ASAP7_75t_R g1209 ( 
.A(n_1109),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_989),
.B(n_663),
.Y(n_1210)
);

OAI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1092),
.A2(n_808),
.B1(n_844),
.B2(n_800),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_989),
.B(n_663),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_989),
.B(n_663),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_1083),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1092),
.B(n_997),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_1021),
.B(n_1084),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_989),
.B(n_663),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_1021),
.B(n_1084),
.Y(n_1218)
);

O2A1O1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_1092),
.A2(n_948),
.B(n_808),
.C(n_844),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_982),
.Y(n_1220)
);

INVx2_ASAP7_75t_SL g1221 ( 
.A(n_1005),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_989),
.B(n_663),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_989),
.B(n_663),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_989),
.B(n_663),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_1026),
.Y(n_1225)
);

CKINVDCx9p33_ASAP7_75t_R g1226 ( 
.A(n_1092),
.Y(n_1226)
);

BUFx12f_ASAP7_75t_L g1227 ( 
.A(n_1026),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1001),
.A2(n_1002),
.B(n_980),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1092),
.A2(n_808),
.B1(n_948),
.B2(n_844),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_989),
.B(n_663),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1005),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_982),
.Y(n_1232)
);

BUFx8_ASAP7_75t_SL g1233 ( 
.A(n_1026),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_1026),
.Y(n_1234)
);

INVx2_ASAP7_75t_SL g1235 ( 
.A(n_1005),
.Y(n_1235)
);

NAND2x1p5_ASAP7_75t_L g1236 ( 
.A(n_992),
.B(n_1083),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_1083),
.Y(n_1237)
);

INVxp67_ASAP7_75t_SL g1238 ( 
.A(n_992),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_989),
.B(n_663),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_982),
.Y(n_1240)
);

CKINVDCx20_ASAP7_75t_R g1241 ( 
.A(n_1109),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1092),
.B(n_997),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1069),
.A2(n_948),
.B(n_808),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1083),
.Y(n_1244)
);

CKINVDCx16_ASAP7_75t_R g1245 ( 
.A(n_1026),
.Y(n_1245)
);

BUFx3_ASAP7_75t_L g1246 ( 
.A(n_1005),
.Y(n_1246)
);

INVx1_ASAP7_75t_SL g1247 ( 
.A(n_1075),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1001),
.A2(n_1002),
.B(n_980),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_982),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_1005),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1079),
.A2(n_808),
.B1(n_995),
.B2(n_962),
.Y(n_1251)
);

OR2x6_ASAP7_75t_L g1252 ( 
.A(n_1078),
.B(n_1057),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1092),
.B(n_997),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_1106),
.Y(n_1254)
);

OR2x6_ASAP7_75t_L g1255 ( 
.A(n_1078),
.B(n_1057),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1114),
.A2(n_1242),
.B1(n_1215),
.B2(n_1253),
.Y(n_1256)
);

INVx3_ASAP7_75t_L g1257 ( 
.A(n_1119),
.Y(n_1257)
);

OAI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1229),
.A2(n_1219),
.B(n_1243),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1127),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1132),
.Y(n_1260)
);

OAI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1251),
.A2(n_1121),
.B(n_1211),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1121),
.B(n_1152),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1211),
.A2(n_1251),
.B1(n_1129),
.B2(n_1146),
.Y(n_1263)
);

AOI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1181),
.A2(n_1228),
.B(n_1115),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1117),
.B(n_1159),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1117),
.A2(n_1174),
.B1(n_1129),
.B2(n_1139),
.Y(n_1266)
);

INVx8_ASAP7_75t_L g1267 ( 
.A(n_1142),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1149),
.Y(n_1268)
);

OA21x2_ASAP7_75t_L g1269 ( 
.A1(n_1189),
.A2(n_1158),
.B(n_1248),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1151),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1152),
.B(n_1155),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1200),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1167),
.A2(n_1155),
.B1(n_1134),
.B2(n_1131),
.Y(n_1273)
);

AND2x4_ASAP7_75t_L g1274 ( 
.A(n_1172),
.B(n_1176),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_SL g1275 ( 
.A1(n_1147),
.A2(n_1226),
.B1(n_1161),
.B2(n_1164),
.Y(n_1275)
);

OAI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1174),
.A2(n_1133),
.B1(n_1130),
.B2(n_1207),
.Y(n_1276)
);

OAI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1150),
.A2(n_1157),
.B1(n_1182),
.B2(n_1255),
.Y(n_1277)
);

AND2x4_ASAP7_75t_L g1278 ( 
.A(n_1172),
.B(n_1176),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_SL g1279 ( 
.A1(n_1226),
.A2(n_1148),
.B1(n_1177),
.B2(n_1124),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1209),
.Y(n_1280)
);

AO21x2_ASAP7_75t_L g1281 ( 
.A1(n_1178),
.A2(n_1203),
.B(n_1116),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1134),
.A2(n_1131),
.B1(n_1128),
.B2(n_1137),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1128),
.A2(n_1138),
.B1(n_1212),
.B2(n_1213),
.Y(n_1283)
);

BUFx2_ASAP7_75t_R g1284 ( 
.A(n_1233),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_SL g1285 ( 
.A1(n_1162),
.A2(n_1163),
.B(n_1217),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_1128),
.Y(n_1286)
);

BUFx3_ASAP7_75t_L g1287 ( 
.A(n_1231),
.Y(n_1287)
);

INVxp67_ASAP7_75t_SL g1288 ( 
.A(n_1125),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_SL g1289 ( 
.A1(n_1210),
.A2(n_1224),
.B1(n_1239),
.B2(n_1222),
.Y(n_1289)
);

BUFx2_ASAP7_75t_R g1290 ( 
.A(n_1233),
.Y(n_1290)
);

CKINVDCx11_ASAP7_75t_R g1291 ( 
.A(n_1227),
.Y(n_1291)
);

CKINVDCx6p67_ASAP7_75t_R g1292 ( 
.A(n_1209),
.Y(n_1292)
);

NAND2x1p5_ASAP7_75t_L g1293 ( 
.A(n_1206),
.B(n_1195),
.Y(n_1293)
);

OA21x2_ASAP7_75t_L g1294 ( 
.A1(n_1162),
.A2(n_1203),
.B(n_1163),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1128),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1220),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1232),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1240),
.Y(n_1298)
);

OAI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1252),
.A2(n_1255),
.B1(n_1166),
.B2(n_1126),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1249),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1128),
.A2(n_1223),
.B1(n_1230),
.B2(n_1173),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1183),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1191),
.Y(n_1303)
);

INVx3_ASAP7_75t_L g1304 ( 
.A(n_1199),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1252),
.A2(n_1255),
.B1(n_1188),
.B2(n_1171),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1187),
.Y(n_1306)
);

CKINVDCx11_ASAP7_75t_R g1307 ( 
.A(n_1227),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1254),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1165),
.A2(n_1185),
.B(n_1205),
.Y(n_1309)
);

BUFx12f_ASAP7_75t_L g1310 ( 
.A(n_1123),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1122),
.B(n_1143),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1231),
.Y(n_1312)
);

INVx1_ASAP7_75t_SL g1313 ( 
.A(n_1247),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1196),
.Y(n_1314)
);

AO21x2_ASAP7_75t_L g1315 ( 
.A1(n_1198),
.A2(n_1204),
.B(n_1194),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1206),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1201),
.B(n_1202),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1193),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1201),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_SL g1320 ( 
.A1(n_1169),
.A2(n_1238),
.B1(n_1118),
.B2(n_1241),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1216),
.B(n_1218),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1169),
.Y(n_1322)
);

INVx11_ASAP7_75t_L g1323 ( 
.A(n_1156),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1186),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1216),
.A2(n_1168),
.B1(n_1141),
.B2(n_1144),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1236),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1168),
.A2(n_1144),
.B1(n_1145),
.B2(n_1180),
.Y(n_1327)
);

BUFx2_ASAP7_75t_L g1328 ( 
.A(n_1184),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1184),
.Y(n_1329)
);

OA21x2_ASAP7_75t_L g1330 ( 
.A1(n_1179),
.A2(n_1197),
.B(n_1180),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1192),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1160),
.A2(n_1140),
.B1(n_1250),
.B2(n_1246),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_SL g1333 ( 
.A1(n_1238),
.A2(n_1118),
.B1(n_1241),
.B2(n_1250),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1170),
.B(n_1154),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1192),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1214),
.Y(n_1336)
);

CKINVDCx11_ASAP7_75t_R g1337 ( 
.A(n_1245),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1136),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_1120),
.Y(n_1339)
);

INVx1_ASAP7_75t_SL g1340 ( 
.A(n_1153),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_SL g1341 ( 
.A1(n_1246),
.A2(n_1235),
.B1(n_1221),
.B2(n_1135),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1208),
.A2(n_1175),
.B1(n_1190),
.B2(n_1237),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1208),
.A2(n_1175),
.B1(n_1190),
.B2(n_1244),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1225),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1234),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1128),
.Y(n_1346)
);

BUFx2_ASAP7_75t_L g1347 ( 
.A(n_1128),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1121),
.A2(n_957),
.B1(n_808),
.B2(n_844),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_SL g1349 ( 
.A1(n_1229),
.A2(n_719),
.B1(n_950),
.B2(n_800),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1121),
.A2(n_957),
.B1(n_808),
.B2(n_844),
.Y(n_1350)
);

BUFx2_ASAP7_75t_SL g1351 ( 
.A(n_1142),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1172),
.B(n_1176),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1121),
.B(n_1152),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1114),
.A2(n_1092),
.B1(n_808),
.B2(n_948),
.Y(n_1354)
);

CKINVDCx10_ASAP7_75t_R g1355 ( 
.A(n_1245),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1119),
.Y(n_1356)
);

OAI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1114),
.A2(n_719),
.B1(n_808),
.B2(n_800),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1272),
.Y(n_1358)
);

AO21x2_ASAP7_75t_L g1359 ( 
.A1(n_1258),
.A2(n_1264),
.B(n_1261),
.Y(n_1359)
);

BUFx2_ASAP7_75t_L g1360 ( 
.A(n_1293),
.Y(n_1360)
);

OAI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1348),
.A2(n_1350),
.B(n_1354),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1293),
.Y(n_1362)
);

CKINVDCx14_ASAP7_75t_R g1363 ( 
.A(n_1337),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_SL g1364 ( 
.A1(n_1266),
.A2(n_1330),
.B(n_1265),
.Y(n_1364)
);

OR2x2_ASAP7_75t_L g1365 ( 
.A(n_1293),
.B(n_1281),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1271),
.B(n_1262),
.Y(n_1366)
);

INVx1_ASAP7_75t_SL g1367 ( 
.A(n_1328),
.Y(n_1367)
);

OAI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1357),
.A2(n_1256),
.B1(n_1277),
.B2(n_1314),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1353),
.B(n_1317),
.Y(n_1369)
);

CKINVDCx20_ASAP7_75t_R g1370 ( 
.A(n_1337),
.Y(n_1370)
);

HB1xp67_ASAP7_75t_L g1371 ( 
.A(n_1288),
.Y(n_1371)
);

INVx2_ASAP7_75t_SL g1372 ( 
.A(n_1308),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1353),
.B(n_1317),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1276),
.B(n_1273),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1309),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1324),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1281),
.B(n_1294),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1324),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1309),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1329),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_1286),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1295),
.B(n_1346),
.Y(n_1382)
);

AO21x2_ASAP7_75t_L g1383 ( 
.A1(n_1281),
.A2(n_1315),
.B(n_1316),
.Y(n_1383)
);

OR2x6_ASAP7_75t_L g1384 ( 
.A(n_1295),
.B(n_1346),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1316),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1319),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1269),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1269),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1294),
.B(n_1347),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1269),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1282),
.B(n_1319),
.Y(n_1391)
);

OR2x6_ASAP7_75t_L g1392 ( 
.A(n_1330),
.B(n_1351),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1294),
.Y(n_1393)
);

AO21x1_ASAP7_75t_SL g1394 ( 
.A1(n_1263),
.A2(n_1301),
.B(n_1283),
.Y(n_1394)
);

NAND2x1p5_ASAP7_75t_L g1395 ( 
.A(n_1330),
.B(n_1318),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_1287),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1314),
.B(n_1260),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1331),
.Y(n_1398)
);

BUFx4f_ASAP7_75t_SL g1399 ( 
.A(n_1310),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1335),
.Y(n_1400)
);

INVxp67_ASAP7_75t_SL g1401 ( 
.A(n_1311),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1285),
.B(n_1297),
.Y(n_1402)
);

OA21x2_ASAP7_75t_L g1403 ( 
.A1(n_1298),
.A2(n_1300),
.B(n_1259),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1315),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1268),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1270),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1334),
.B(n_1296),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1302),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1306),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1305),
.B(n_1299),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1303),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1326),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1289),
.B(n_1352),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1287),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1336),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1338),
.Y(n_1416)
);

INVx1_ASAP7_75t_SL g1417 ( 
.A(n_1313),
.Y(n_1417)
);

INVx1_ASAP7_75t_SL g1418 ( 
.A(n_1322),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1275),
.B(n_1349),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1396),
.Y(n_1420)
);

OR2x6_ASAP7_75t_L g1421 ( 
.A(n_1392),
.B(n_1267),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1358),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1393),
.B(n_1279),
.Y(n_1423)
);

INVx2_ASAP7_75t_SL g1424 ( 
.A(n_1375),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1401),
.B(n_1327),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1360),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1361),
.A2(n_1322),
.B1(n_1352),
.B2(n_1274),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1383),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1371),
.B(n_1333),
.Y(n_1429)
);

INVxp67_ASAP7_75t_L g1430 ( 
.A(n_1380),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1387),
.B(n_1388),
.Y(n_1431)
);

BUFx2_ASAP7_75t_L g1432 ( 
.A(n_1360),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1403),
.B(n_1320),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1403),
.B(n_1257),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1403),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1403),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1361),
.A2(n_1352),
.B1(n_1274),
.B2(n_1278),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1390),
.B(n_1278),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1389),
.B(n_1312),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1390),
.B(n_1278),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1394),
.A2(n_1274),
.B1(n_1292),
.B2(n_1321),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1405),
.B(n_1356),
.Y(n_1442)
);

OA21x2_ASAP7_75t_L g1443 ( 
.A1(n_1404),
.A2(n_1325),
.B(n_1342),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1405),
.B(n_1356),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1390),
.B(n_1356),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1389),
.B(n_1312),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1379),
.Y(n_1447)
);

INVx1_ASAP7_75t_SL g1448 ( 
.A(n_1367),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1375),
.B(n_1304),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1395),
.B(n_1332),
.Y(n_1450)
);

AND2x4_ASAP7_75t_SL g1451 ( 
.A(n_1384),
.B(n_1381),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1395),
.B(n_1345),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1394),
.A2(n_1292),
.B1(n_1321),
.B2(n_1345),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1417),
.B(n_1340),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1438),
.B(n_1384),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1438),
.B(n_1384),
.Y(n_1456)
);

NAND3xp33_ASAP7_75t_L g1457 ( 
.A(n_1450),
.B(n_1419),
.C(n_1402),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1425),
.A2(n_1419),
.B1(n_1368),
.B2(n_1374),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1425),
.A2(n_1364),
.B(n_1359),
.Y(n_1459)
);

NAND3xp33_ASAP7_75t_L g1460 ( 
.A(n_1450),
.B(n_1402),
.C(n_1374),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1422),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1453),
.A2(n_1410),
.B1(n_1363),
.B2(n_1418),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1452),
.B(n_1418),
.Y(n_1463)
);

NOR3xp33_ASAP7_75t_L g1464 ( 
.A(n_1429),
.B(n_1410),
.C(n_1454),
.Y(n_1464)
);

NAND3xp33_ASAP7_75t_L g1465 ( 
.A(n_1429),
.B(n_1364),
.C(n_1341),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1448),
.B(n_1366),
.Y(n_1466)
);

AOI221xp5_ASAP7_75t_L g1467 ( 
.A1(n_1433),
.A2(n_1366),
.B1(n_1417),
.B2(n_1409),
.C(n_1397),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1427),
.A2(n_1359),
.B1(n_1391),
.B2(n_1413),
.Y(n_1468)
);

NAND3xp33_ASAP7_75t_L g1469 ( 
.A(n_1433),
.B(n_1378),
.C(n_1376),
.Y(n_1469)
);

NAND3xp33_ASAP7_75t_L g1470 ( 
.A(n_1423),
.B(n_1397),
.C(n_1365),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1441),
.A2(n_1437),
.B1(n_1370),
.B2(n_1343),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1421),
.Y(n_1472)
);

NAND3xp33_ASAP7_75t_L g1473 ( 
.A(n_1423),
.B(n_1365),
.C(n_1412),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1430),
.B(n_1439),
.Y(n_1474)
);

NAND3xp33_ASAP7_75t_L g1475 ( 
.A(n_1423),
.B(n_1412),
.C(n_1413),
.Y(n_1475)
);

NAND3xp33_ASAP7_75t_L g1476 ( 
.A(n_1443),
.B(n_1398),
.C(n_1400),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1439),
.B(n_1407),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1446),
.B(n_1372),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1438),
.B(n_1384),
.Y(n_1479)
);

OAI221xp5_ASAP7_75t_L g1480 ( 
.A1(n_1421),
.A2(n_1280),
.B1(n_1396),
.B2(n_1414),
.C(n_1362),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1440),
.B(n_1384),
.Y(n_1481)
);

OAI221xp5_ASAP7_75t_SL g1482 ( 
.A1(n_1421),
.A2(n_1377),
.B1(n_1392),
.B2(n_1391),
.C(n_1369),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1451),
.A2(n_1280),
.B1(n_1414),
.B2(n_1396),
.Y(n_1483)
);

OAI21xp33_ASAP7_75t_SL g1484 ( 
.A1(n_1442),
.A2(n_1406),
.B(n_1411),
.Y(n_1484)
);

AOI221xp5_ASAP7_75t_L g1485 ( 
.A1(n_1444),
.A2(n_1373),
.B1(n_1406),
.B2(n_1411),
.C(n_1359),
.Y(n_1485)
);

NAND4xp25_ASAP7_75t_L g1486 ( 
.A(n_1444),
.B(n_1415),
.C(n_1416),
.D(n_1408),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_SL g1487 ( 
.A(n_1420),
.B(n_1284),
.Y(n_1487)
);

OAI21xp5_ASAP7_75t_SL g1488 ( 
.A1(n_1451),
.A2(n_1344),
.B(n_1382),
.Y(n_1488)
);

NAND4xp25_ASAP7_75t_L g1489 ( 
.A(n_1434),
.B(n_1415),
.C(n_1416),
.D(n_1408),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1440),
.B(n_1382),
.Y(n_1490)
);

NAND3xp33_ASAP7_75t_L g1491 ( 
.A(n_1443),
.B(n_1385),
.C(n_1386),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1443),
.A2(n_1359),
.B1(n_1321),
.B2(n_1399),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1485),
.B(n_1484),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1472),
.Y(n_1494)
);

CKINVDCx16_ASAP7_75t_R g1495 ( 
.A(n_1487),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1474),
.B(n_1344),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1461),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1472),
.B(n_1490),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1455),
.B(n_1421),
.Y(n_1499)
);

INVx1_ASAP7_75t_SL g1500 ( 
.A(n_1478),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1490),
.B(n_1431),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1455),
.B(n_1431),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1456),
.B(n_1479),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1459),
.B(n_1422),
.Y(n_1504)
);

NOR2x1_ASAP7_75t_L g1505 ( 
.A(n_1476),
.B(n_1435),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1481),
.Y(n_1506)
);

INVxp67_ASAP7_75t_L g1507 ( 
.A(n_1463),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1491),
.B(n_1436),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1481),
.B(n_1492),
.Y(n_1509)
);

INVx3_ASAP7_75t_L g1510 ( 
.A(n_1477),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1492),
.B(n_1436),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1470),
.B(n_1440),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1473),
.B(n_1421),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1489),
.B(n_1434),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1475),
.B(n_1421),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1486),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1469),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1466),
.B(n_1428),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1468),
.B(n_1445),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1460),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1457),
.Y(n_1521)
);

INVx2_ASAP7_75t_SL g1522 ( 
.A(n_1483),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1506),
.B(n_1451),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1514),
.B(n_1482),
.Y(n_1524)
);

INVxp67_ASAP7_75t_L g1525 ( 
.A(n_1520),
.Y(n_1525)
);

INVxp67_ASAP7_75t_L g1526 ( 
.A(n_1520),
.Y(n_1526)
);

INVx3_ASAP7_75t_L g1527 ( 
.A(n_1499),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1497),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1514),
.B(n_1426),
.Y(n_1529)
);

INVx2_ASAP7_75t_SL g1530 ( 
.A(n_1494),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1508),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1508),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1497),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1514),
.B(n_1426),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1504),
.B(n_1432),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1516),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1518),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1521),
.B(n_1464),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1506),
.B(n_1488),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1499),
.B(n_1424),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1518),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1496),
.B(n_1344),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1518),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1521),
.B(n_1467),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1498),
.B(n_1499),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1501),
.Y(n_1546)
);

NOR2xp67_ASAP7_75t_L g1547 ( 
.A(n_1493),
.B(n_1465),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1493),
.B(n_1447),
.Y(n_1548)
);

INVx2_ASAP7_75t_SL g1549 ( 
.A(n_1499),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1499),
.B(n_1424),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1501),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1503),
.B(n_1449),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1501),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1508),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1528),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1531),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1528),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1547),
.A2(n_1521),
.B1(n_1522),
.B2(n_1517),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1548),
.B(n_1517),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1547),
.B(n_1538),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1545),
.B(n_1515),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1545),
.B(n_1515),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1533),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1549),
.B(n_1515),
.Y(n_1564)
);

NAND2x1_ASAP7_75t_L g1565 ( 
.A(n_1530),
.B(n_1505),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1539),
.B(n_1503),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1539),
.B(n_1503),
.Y(n_1567)
);

INVxp67_ASAP7_75t_L g1568 ( 
.A(n_1536),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1533),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1527),
.B(n_1513),
.Y(n_1570)
);

NOR2xp67_ASAP7_75t_L g1571 ( 
.A(n_1527),
.B(n_1522),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1527),
.B(n_1513),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1544),
.B(n_1516),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1549),
.B(n_1513),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1548),
.B(n_1510),
.Y(n_1575)
);

A2O1A1Ixp33_ASAP7_75t_L g1576 ( 
.A1(n_1524),
.A2(n_1505),
.B(n_1458),
.C(n_1522),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1537),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1537),
.Y(n_1578)
);

INVx1_ASAP7_75t_SL g1579 ( 
.A(n_1529),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1541),
.B(n_1510),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1525),
.B(n_1507),
.Y(n_1581)
);

AND2x4_ASAP7_75t_L g1582 ( 
.A(n_1527),
.B(n_1509),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1531),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1541),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1552),
.B(n_1509),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1543),
.Y(n_1586)
);

OR2x6_ASAP7_75t_L g1587 ( 
.A(n_1526),
.B(n_1392),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1524),
.B(n_1507),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1543),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1531),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1546),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1546),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1552),
.B(n_1509),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1523),
.B(n_1502),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1535),
.B(n_1500),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_1529),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1535),
.B(n_1500),
.Y(n_1597)
);

NOR2x1_ASAP7_75t_L g1598 ( 
.A(n_1576),
.B(n_1554),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1555),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1557),
.Y(n_1600)
);

NOR2x1_ASAP7_75t_L g1601 ( 
.A(n_1576),
.B(n_1554),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1563),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1573),
.B(n_1532),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1556),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1582),
.B(n_1532),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1569),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1577),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1560),
.A2(n_1468),
.B1(n_1458),
.B2(n_1480),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1556),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1588),
.A2(n_1462),
.B1(n_1542),
.B2(n_1519),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1568),
.Y(n_1611)
);

INVx1_ASAP7_75t_SL g1612 ( 
.A(n_1565),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1579),
.Y(n_1613)
);

INVx3_ASAP7_75t_L g1614 ( 
.A(n_1565),
.Y(n_1614)
);

INVx1_ASAP7_75t_SL g1615 ( 
.A(n_1559),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1578),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1559),
.Y(n_1617)
);

OAI21xp33_ASAP7_75t_L g1618 ( 
.A1(n_1558),
.A2(n_1511),
.B(n_1519),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1584),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1586),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1589),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1582),
.B(n_1540),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1582),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1585),
.B(n_1540),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1581),
.B(n_1551),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1595),
.B(n_1290),
.Y(n_1626)
);

INVx4_ASAP7_75t_L g1627 ( 
.A(n_1583),
.Y(n_1627)
);

INVx1_ASAP7_75t_SL g1628 ( 
.A(n_1596),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1583),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1585),
.B(n_1540),
.Y(n_1630)
);

INVx3_ASAP7_75t_L g1631 ( 
.A(n_1587),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1566),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1593),
.B(n_1540),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1628),
.B(n_1566),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1626),
.B(n_1291),
.Y(n_1635)
);

INVxp67_ASAP7_75t_L g1636 ( 
.A(n_1598),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1613),
.Y(n_1637)
);

OAI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1598),
.A2(n_1495),
.B1(n_1571),
.B2(n_1567),
.Y(n_1638)
);

NAND3xp33_ASAP7_75t_L g1639 ( 
.A(n_1601),
.B(n_1590),
.C(n_1597),
.Y(n_1639)
);

INVxp67_ASAP7_75t_L g1640 ( 
.A(n_1601),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1632),
.B(n_1567),
.Y(n_1641)
);

OAI21xp5_ASAP7_75t_SL g1642 ( 
.A1(n_1608),
.A2(n_1574),
.B(n_1564),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1613),
.Y(n_1643)
);

AOI322xp5_ASAP7_75t_L g1644 ( 
.A1(n_1618),
.A2(n_1593),
.A3(n_1519),
.B1(n_1562),
.B2(n_1561),
.C1(n_1512),
.C2(n_1553),
.Y(n_1644)
);

OAI322xp33_ASAP7_75t_L g1645 ( 
.A1(n_1611),
.A2(n_1575),
.A3(n_1580),
.B1(n_1591),
.B2(n_1592),
.C1(n_1534),
.C2(n_1590),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1632),
.B(n_1594),
.Y(n_1646)
);

AOI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1618),
.A2(n_1574),
.B1(n_1495),
.B2(n_1564),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1628),
.B(n_1594),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1623),
.B(n_1561),
.Y(n_1649)
);

INVxp67_ASAP7_75t_L g1650 ( 
.A(n_1611),
.Y(n_1650)
);

AOI222xp33_ASAP7_75t_L g1651 ( 
.A1(n_1610),
.A2(n_1511),
.B1(n_1574),
.B2(n_1564),
.C1(n_1561),
.C2(n_1562),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1615),
.B(n_1562),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1599),
.Y(n_1653)
);

OAI22xp33_ASAP7_75t_SL g1654 ( 
.A1(n_1612),
.A2(n_1587),
.B1(n_1575),
.B2(n_1580),
.Y(n_1654)
);

NOR2x1_ASAP7_75t_L g1655 ( 
.A(n_1614),
.B(n_1534),
.Y(n_1655)
);

NAND2xp33_ASAP7_75t_SL g1656 ( 
.A(n_1623),
.B(n_1530),
.Y(n_1656)
);

AOI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1622),
.A2(n_1572),
.B1(n_1570),
.B2(n_1587),
.Y(n_1657)
);

OAI21xp33_ASAP7_75t_L g1658 ( 
.A1(n_1603),
.A2(n_1572),
.B(n_1570),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1623),
.B(n_1550),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1649),
.B(n_1623),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1636),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1636),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1641),
.B(n_1622),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1637),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1640),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1643),
.B(n_1615),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1640),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_1650),
.Y(n_1668)
);

INVx1_ASAP7_75t_SL g1669 ( 
.A(n_1656),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1650),
.B(n_1617),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1634),
.B(n_1617),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1653),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1648),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1638),
.A2(n_1622),
.B1(n_1625),
.B2(n_1603),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1655),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1646),
.B(n_1605),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1635),
.B(n_1291),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1659),
.B(n_1647),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1642),
.B(n_1605),
.Y(n_1679)
);

OAI211xp5_ASAP7_75t_L g1680 ( 
.A1(n_1667),
.A2(n_1639),
.B(n_1651),
.C(n_1644),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1670),
.Y(n_1681)
);

NOR3xp33_ASAP7_75t_L g1682 ( 
.A(n_1666),
.B(n_1652),
.C(n_1645),
.Y(n_1682)
);

OAI211xp5_ASAP7_75t_L g1683 ( 
.A1(n_1669),
.A2(n_1612),
.B(n_1658),
.C(n_1657),
.Y(n_1683)
);

AOI221x1_ASAP7_75t_L g1684 ( 
.A1(n_1661),
.A2(n_1654),
.B1(n_1614),
.B2(n_1607),
.C(n_1616),
.Y(n_1684)
);

NOR3xp33_ASAP7_75t_L g1685 ( 
.A(n_1668),
.B(n_1307),
.C(n_1614),
.Y(n_1685)
);

AOI221x1_ASAP7_75t_L g1686 ( 
.A1(n_1661),
.A2(n_1614),
.B1(n_1607),
.B2(n_1616),
.C(n_1620),
.Y(n_1686)
);

OAI211xp5_ASAP7_75t_L g1687 ( 
.A1(n_1675),
.A2(n_1631),
.B(n_1627),
.C(n_1605),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1670),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1668),
.B(n_1619),
.Y(n_1689)
);

NOR3x1_ASAP7_75t_L g1690 ( 
.A(n_1679),
.B(n_1625),
.C(n_1620),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1663),
.B(n_1619),
.Y(n_1691)
);

AOI211x1_ASAP7_75t_SL g1692 ( 
.A1(n_1675),
.A2(n_1604),
.B(n_1629),
.C(n_1609),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1681),
.B(n_1673),
.Y(n_1693)
);

NOR2x1_ASAP7_75t_L g1694 ( 
.A(n_1688),
.B(n_1662),
.Y(n_1694)
);

NOR2x1_ASAP7_75t_L g1695 ( 
.A(n_1687),
.B(n_1662),
.Y(n_1695)
);

NAND4xp75_ASAP7_75t_L g1696 ( 
.A(n_1684),
.B(n_1665),
.C(n_1664),
.D(n_1678),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1682),
.B(n_1673),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1691),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1689),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1685),
.B(n_1678),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1683),
.B(n_1677),
.Y(n_1701)
);

INVx2_ASAP7_75t_SL g1702 ( 
.A(n_1686),
.Y(n_1702)
);

AOI211xp5_ASAP7_75t_L g1703 ( 
.A1(n_1680),
.A2(n_1665),
.B(n_1672),
.C(n_1671),
.Y(n_1703)
);

NAND4xp75_ASAP7_75t_L g1704 ( 
.A(n_1695),
.B(n_1690),
.C(n_1660),
.D(n_1663),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1696),
.B(n_1660),
.Y(n_1705)
);

AOI211x1_ASAP7_75t_SL g1706 ( 
.A1(n_1697),
.A2(n_1676),
.B(n_1680),
.C(n_1692),
.Y(n_1706)
);

NAND4xp25_ASAP7_75t_L g1707 ( 
.A(n_1701),
.B(n_1674),
.C(n_1631),
.D(n_1627),
.Y(n_1707)
);

AOI221xp5_ASAP7_75t_SL g1708 ( 
.A1(n_1703),
.A2(n_1621),
.B1(n_1602),
.B2(n_1606),
.C(n_1599),
.Y(n_1708)
);

OAI211xp5_ASAP7_75t_SL g1709 ( 
.A1(n_1703),
.A2(n_1307),
.B(n_1631),
.C(n_1621),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1700),
.B(n_1624),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1710),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1705),
.B(n_1694),
.Y(n_1712)
);

OAI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1704),
.A2(n_1702),
.B(n_1693),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1706),
.Y(n_1714)
);

AOI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1709),
.A2(n_1707),
.B1(n_1699),
.B2(n_1698),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1708),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1711),
.B(n_1600),
.Y(n_1717)
);

HB1xp67_ASAP7_75t_L g1718 ( 
.A(n_1712),
.Y(n_1718)
);

NAND2x1p5_ASAP7_75t_L g1719 ( 
.A(n_1715),
.B(n_1344),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1713),
.Y(n_1720)
);

NAND4xp75_ASAP7_75t_L g1721 ( 
.A(n_1714),
.B(n_1606),
.C(n_1600),
.D(n_1602),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1720),
.B(n_1716),
.Y(n_1722)
);

XNOR2x1_ASAP7_75t_L g1723 ( 
.A(n_1719),
.B(n_1339),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1721),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1722),
.Y(n_1725)
);

NAND3xp33_ASAP7_75t_L g1726 ( 
.A(n_1725),
.B(n_1718),
.C(n_1724),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1726),
.Y(n_1727)
);

AOI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1726),
.A2(n_1723),
.B(n_1722),
.Y(n_1728)
);

OAI22x1_ASAP7_75t_L g1729 ( 
.A1(n_1727),
.A2(n_1717),
.B1(n_1339),
.B2(n_1355),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1728),
.A2(n_1310),
.B1(n_1627),
.B2(n_1631),
.Y(n_1730)
);

OAI22xp5_ASAP7_75t_SL g1731 ( 
.A1(n_1729),
.A2(n_1344),
.B1(n_1627),
.B2(n_1604),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_SL g1732 ( 
.A1(n_1730),
.A2(n_1629),
.B1(n_1604),
.B2(n_1609),
.Y(n_1732)
);

OAI321xp33_ASAP7_75t_L g1733 ( 
.A1(n_1731),
.A2(n_1629),
.A3(n_1609),
.B1(n_1633),
.B2(n_1630),
.C(n_1624),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1733),
.A2(n_1732),
.B1(n_1633),
.B2(n_1630),
.Y(n_1734)
);

OAI221xp5_ASAP7_75t_R g1735 ( 
.A1(n_1734),
.A2(n_1323),
.B1(n_1267),
.B2(n_1633),
.C(n_1624),
.Y(n_1735)
);

AOI211xp5_ASAP7_75t_L g1736 ( 
.A1(n_1735),
.A2(n_1630),
.B(n_1323),
.C(n_1471),
.Y(n_1736)
);


endmodule