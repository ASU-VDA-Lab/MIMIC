module fake_jpeg_13731_n_415 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_415);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_415;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_12),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_7),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_61),
.Y(n_75)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_41),
.Y(n_106)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_18),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_44),
.Y(n_82)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_47),
.B(n_50),
.Y(n_94)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_56),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_20),
.B(n_6),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_58),
.B(n_37),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_20),
.B(n_36),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_28),
.B(n_6),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_28),
.B(n_14),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_71),
.Y(n_105)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_31),
.B(n_14),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_72),
.B(n_10),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_78),
.B(n_86),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_42),
.A2(n_31),
.B1(n_36),
.B2(n_32),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_79),
.A2(n_91),
.B1(n_109),
.B2(n_17),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_45),
.A2(n_18),
.B1(n_15),
.B2(n_23),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_83),
.B(n_82),
.C(n_106),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_46),
.B(n_32),
.Y(n_86)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_23),
.B1(n_33),
.B2(n_18),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_89),
.A2(n_23),
.B1(n_33),
.B2(n_18),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_40),
.A2(n_37),
.B1(n_29),
.B2(n_26),
.Y(n_91)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_112),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_55),
.A2(n_37),
.B1(n_29),
.B2(n_26),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_44),
.B(n_15),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_17),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_113),
.B(n_21),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_116),
.B(n_128),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_117),
.A2(n_118),
.B1(n_137),
.B2(n_74),
.Y(n_159)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_121),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_70),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_124),
.C(n_77),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_104),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_135),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_60),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_80),
.B(n_66),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_139),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_96),
.Y(n_126)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_127),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_89),
.A2(n_67),
.B1(n_65),
.B2(n_59),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_131),
.A2(n_138),
.B1(n_143),
.B2(n_73),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_132),
.B(n_123),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_75),
.B(n_25),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_133),
.B(n_144),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_104),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_136),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_25),
.B1(n_29),
.B2(n_26),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_83),
.A2(n_29),
.B1(n_26),
.B2(n_19),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_90),
.A2(n_25),
.B(n_57),
.C(n_27),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_83),
.A2(n_21),
.B1(n_1),
.B2(n_2),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_21),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_81),
.B(n_6),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_145),
.B(n_148),
.Y(n_190)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_153),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_95),
.B(n_0),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_150),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_82),
.B(n_5),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_0),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_151),
.Y(n_172)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_154),
.B(n_155),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_99),
.B(n_5),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_153),
.A2(n_101),
.B(n_88),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_157),
.A2(n_173),
.B(n_142),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_159),
.B(n_171),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_118),
.A2(n_77),
.B1(n_73),
.B2(n_100),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_160),
.B(n_175),
.Y(n_221)
);

FAx1_ASAP7_75t_SL g162 ( 
.A(n_125),
.B(n_84),
.CI(n_98),
.CON(n_162),
.SN(n_162)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_162),
.B(n_170),
.Y(n_200)
);

XNOR2x1_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_126),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_168),
.A2(n_187),
.B1(n_195),
.B2(n_127),
.Y(n_197)
);

FAx1_ASAP7_75t_SL g170 ( 
.A(n_150),
.B(n_84),
.CI(n_10),
.CON(n_170),
.SN(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_133),
.A2(n_74),
.B1(n_103),
.B2(n_85),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_134),
.A2(n_110),
.B(n_103),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_110),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_122),
.B(n_5),
.C(n_11),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_181),
.C(n_192),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_122),
.B(n_8),
.C(n_11),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_124),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_129),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_184),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_139),
.A2(n_0),
.B(n_1),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_185),
.A2(n_126),
.B(n_1),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_138),
.A2(n_8),
.B1(n_11),
.B2(n_3),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_115),
.A2(n_8),
.B1(n_11),
.B2(n_3),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_189),
.B(n_13),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_124),
.B(n_8),
.Y(n_192)
);

OA22x2_ASAP7_75t_L g193 ( 
.A1(n_143),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_160),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_L g195 ( 
.A1(n_131),
.A2(n_154),
.B1(n_152),
.B2(n_136),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_168),
.A2(n_155),
.B1(n_152),
.B2(n_149),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_196),
.A2(n_197),
.B1(n_212),
.B2(n_214),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_166),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_198),
.B(n_202),
.Y(n_266)
);

A2O1A1O1Ixp25_ASAP7_75t_L g201 ( 
.A1(n_163),
.A2(n_116),
.B(n_132),
.C(n_140),
.D(n_146),
.Y(n_201)
);

NOR2x1_ASAP7_75t_R g259 ( 
.A(n_201),
.B(n_174),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_222),
.Y(n_239)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_186),
.Y(n_204)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_204),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_165),
.B(n_163),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_206),
.Y(n_241)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_207),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_166),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_208),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_157),
.A2(n_135),
.B(n_120),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_209),
.A2(n_167),
.B(n_173),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_166),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_210),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_211),
.A2(n_219),
.B(n_185),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_162),
.A2(n_152),
.B1(n_121),
.B2(n_119),
.Y(n_212)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_174),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_213),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_187),
.A2(n_120),
.B1(n_156),
.B2(n_129),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_215),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_216),
.A2(n_217),
.B1(n_223),
.B2(n_179),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_162),
.A2(n_142),
.B1(n_141),
.B2(n_10),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_218),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_167),
.A2(n_141),
.B(n_9),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_177),
.Y(n_220)
);

OAI21xp33_ASAP7_75t_SL g248 ( 
.A1(n_220),
.A2(n_225),
.B(n_188),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_165),
.B(n_142),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_167),
.A2(n_10),
.B1(n_4),
.B2(n_9),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_175),
.B(n_4),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_232),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_178),
.B(n_9),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_227),
.B(n_183),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_180),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_228),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_180),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_229),
.Y(n_268)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_230),
.Y(n_260)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_177),
.Y(n_231)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_170),
.B(n_194),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_158),
.Y(n_233)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_233),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_161),
.Y(n_234)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_234),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_235),
.A2(n_238),
.B(n_202),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_164),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_237),
.B(n_253),
.C(n_254),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_221),
.A2(n_195),
.B1(n_176),
.B2(n_193),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_243),
.A2(n_248),
.B1(n_252),
.B2(n_223),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_246),
.B(n_200),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_225),
.A2(n_190),
.B1(n_170),
.B2(n_193),
.Y(n_252)
);

MAJx2_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_205),
.C(n_222),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_203),
.B(n_192),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_197),
.A2(n_193),
.B1(n_172),
.B2(n_181),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_255),
.A2(n_258),
.B1(n_221),
.B2(n_209),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_200),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_205),
.B(n_188),
.C(n_169),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_265),
.C(n_270),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_224),
.A2(n_158),
.B1(n_169),
.B2(n_183),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_211),
.Y(n_284)
);

OAI22x1_ASAP7_75t_L g261 ( 
.A1(n_216),
.A2(n_161),
.B1(n_201),
.B2(n_224),
.Y(n_261)
);

OA22x2_ASAP7_75t_L g298 ( 
.A1(n_261),
.A2(n_229),
.B1(n_228),
.B2(n_218),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_198),
.B(n_210),
.C(n_208),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_224),
.A2(n_196),
.B1(n_217),
.B2(n_212),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_269),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_219),
.B(n_226),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_271),
.A2(n_265),
.B1(n_261),
.B2(n_244),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_249),
.B(n_199),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_274),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g325 ( 
.A(n_275),
.Y(n_325)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_247),
.Y(n_277)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_277),
.Y(n_308)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_247),
.Y(n_278)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_278),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_251),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_281),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_199),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_280),
.B(n_292),
.Y(n_313)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_282),
.B(n_285),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_283),
.B(n_289),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_284),
.B(n_300),
.Y(n_305)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_240),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_257),
.B(n_231),
.C(n_220),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_293),
.C(n_239),
.Y(n_310)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_242),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_287),
.B(n_288),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_236),
.B(n_245),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_260),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_250),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_290),
.A2(n_296),
.B1(n_297),
.B2(n_299),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_241),
.B(n_230),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_291),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_249),
.B(n_266),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_237),
.B(n_254),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_243),
.B(n_204),
.Y(n_294)
);

MAJx2_ASAP7_75t_L g319 ( 
.A(n_294),
.B(n_264),
.C(n_213),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_268),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_295),
.Y(n_312)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_250),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_298),
.A2(n_214),
.B1(n_258),
.B2(n_235),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_270),
.B(n_207),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_302),
.A2(n_326),
.B1(n_297),
.B2(n_298),
.Y(n_328)
);

A2O1A1Ixp33_ASAP7_75t_L g303 ( 
.A1(n_291),
.A2(n_259),
.B(n_238),
.C(n_253),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_303),
.B(n_298),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_239),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_306),
.B(n_314),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_307),
.A2(n_277),
.B(n_278),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_310),
.B(n_315),
.C(n_318),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_272),
.B(n_255),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_272),
.B(n_273),
.C(n_286),
.Y(n_315)
);

XNOR2x1_ASAP7_75t_SL g316 ( 
.A(n_273),
.B(n_246),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_316),
.B(n_298),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_283),
.B(n_244),
.C(n_233),
.Y(n_318)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_319),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_276),
.A2(n_264),
.B1(n_262),
.B2(n_234),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_320),
.A2(n_285),
.B1(n_289),
.B2(n_287),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_271),
.B(n_262),
.C(n_234),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_322),
.B(n_290),
.C(n_296),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_276),
.A2(n_284),
.B1(n_300),
.B2(n_294),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_328),
.A2(n_341),
.B1(n_342),
.B2(n_343),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_295),
.Y(n_329)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_329),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_312),
.B(n_279),
.Y(n_330)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_330),
.Y(n_358)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_301),
.Y(n_331)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_331),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_321),
.B(n_288),
.Y(n_332)
);

XOR2x2_ASAP7_75t_L g354 ( 
.A(n_332),
.B(n_334),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_301),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_333),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_335),
.B(n_339),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_336),
.B(n_337),
.Y(n_353)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_321),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_311),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_340),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_302),
.A2(n_307),
.B1(n_318),
.B2(n_326),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_304),
.A2(n_322),
.B1(n_303),
.B2(n_309),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_317),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_344),
.A2(n_348),
.B(n_334),
.Y(n_364)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_317),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_345),
.B(n_319),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_325),
.B(n_308),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_347),
.A2(n_324),
.B(n_323),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_305),
.A2(n_281),
.B(n_282),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_356),
.B(n_357),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_338),
.B(n_315),
.C(n_310),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_338),
.B(n_316),
.C(n_314),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_359),
.B(n_360),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_346),
.B(n_306),
.C(n_305),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_346),
.B(n_324),
.C(n_320),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_362),
.B(n_339),
.Y(n_367)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_363),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_364),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_335),
.B(n_342),
.Y(n_365)
);

MAJx2_ASAP7_75t_L g370 ( 
.A(n_365),
.B(n_328),
.C(n_331),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_359),
.A2(n_348),
.B(n_327),
.Y(n_366)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_366),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_367),
.B(n_375),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_357),
.B(n_341),
.C(n_327),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_368),
.B(n_371),
.C(n_360),
.Y(n_386)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_370),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_362),
.B(n_344),
.C(n_345),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_355),
.B(n_358),
.Y(n_373)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_373),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_352),
.B(n_347),
.Y(n_374)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_374),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_363),
.B(n_365),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_349),
.B(n_332),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_376),
.B(n_378),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_351),
.B(n_333),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_379),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_380),
.B(n_385),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_369),
.A2(n_350),
.B1(n_353),
.B2(n_361),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_381),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_369),
.A2(n_350),
.B1(n_337),
.B2(n_343),
.Y(n_383)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_383),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_371),
.A2(n_354),
.B1(n_349),
.B2(n_364),
.Y(n_385)
);

MAJx2_ASAP7_75t_L g398 ( 
.A(n_386),
.B(n_370),
.C(n_354),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_384),
.B(n_372),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_391),
.B(n_392),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_388),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_382),
.A2(n_368),
.B(n_377),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_393),
.B(n_398),
.C(n_386),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g394 ( 
.A(n_383),
.B(n_356),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_394),
.B(n_396),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_384),
.B(n_376),
.Y(n_396)
);

BUFx24_ASAP7_75t_SL g400 ( 
.A(n_397),
.Y(n_400)
);

BUFx24_ASAP7_75t_SL g408 ( 
.A(n_400),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_401),
.B(n_385),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_399),
.B(n_389),
.C(n_388),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_403),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_395),
.B(n_387),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_405),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_406),
.B(n_398),
.C(n_390),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_407),
.A2(n_404),
.B(n_402),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_410),
.B(n_411),
.C(n_406),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_412),
.B(n_409),
.Y(n_413)
);

OAI211xp5_ASAP7_75t_L g414 ( 
.A1(n_413),
.A2(n_408),
.B(n_390),
.C(n_336),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_414),
.B(n_381),
.Y(n_415)
);


endmodule