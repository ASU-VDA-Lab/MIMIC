module real_aes_16755_n_7 (n_4, n_0, n_3, n_5, n_2, n_6, n_1, n_7);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_6;
input n_1;
output n_7;
wire n_28;
wire n_17;
wire n_22;
wire n_13;
wire n_24;
wire n_12;
wire n_19;
wire n_25;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_27;
wire n_9;
wire n_23;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_8;
wire n_10;
INVx2_ASAP7_75t_L g16 ( .A(n_0), .Y(n_16) );
INVx1_ASAP7_75t_L g20 ( .A(n_1), .Y(n_20) );
AND2x2_ASAP7_75t_L g11 ( .A(n_2), .B(n_6), .Y(n_11) );
HB1xp67_ASAP7_75t_L g12 ( .A(n_3), .Y(n_12) );
AND2x2_ASAP7_75t_L g27 ( .A(n_3), .B(n_20), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_4), .B(n_14), .Y(n_13) );
BUFx6f_ASAP7_75t_L g24 ( .A(n_5), .Y(n_24) );
AOI22xp33_ASAP7_75t_L g7 ( .A1(n_8), .A2(n_21), .B1(n_25), .B2(n_28), .Y(n_7) );
INVxp67_ASAP7_75t_SL g8 ( .A(n_9), .Y(n_8) );
AOI221xp5_ASAP7_75t_SL g9 ( .A1(n_10), .A2(n_12), .B1(n_13), .B2(n_17), .C(n_18), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_11), .Y(n_10) );
AND2x2_ASAP7_75t_L g26 ( .A(n_11), .B(n_27), .Y(n_26) );
INVx1_ASAP7_75t_L g17 ( .A(n_12), .Y(n_17) );
INVx2_ASAP7_75t_SL g14 ( .A(n_15), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_16), .Y(n_15) );
INVx1_ASAP7_75t_L g18 ( .A(n_19), .Y(n_18) );
HB1xp67_ASAP7_75t_L g19 ( .A(n_20), .Y(n_19) );
INVx1_ASAP7_75t_L g28 ( .A(n_21), .Y(n_28) );
INVx1_ASAP7_75t_L g21 ( .A(n_22), .Y(n_21) );
HB1xp67_ASAP7_75t_L g22 ( .A(n_23), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_24), .Y(n_23) );
HB1xp67_ASAP7_75t_L g25 ( .A(n_26), .Y(n_25) );
endmodule