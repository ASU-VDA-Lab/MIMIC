module fake_jpeg_3995_n_288 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_288);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_247;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_273;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_9),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_20),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_23),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_41),
.B(n_57),
.Y(n_84)
);

NAND2xp33_ASAP7_75t_SL g42 ( 
.A(n_36),
.B(n_0),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_42),
.A2(n_19),
.B(n_35),
.C(n_33),
.Y(n_86)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_49),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_36),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_48),
.Y(n_77)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_54),
.Y(n_66)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_29),
.Y(n_51)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_58),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_18),
.B(n_1),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

NOR2x1_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_37),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_59),
.B(n_25),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_48),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_60),
.B(n_61),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_56),
.A2(n_28),
.B1(n_34),
.B2(n_30),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_62),
.A2(n_21),
.B1(n_3),
.B2(n_5),
.Y(n_107)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_64),
.B(n_71),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_23),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_69),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_23),
.Y(n_69)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_22),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_72),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_34),
.B1(n_30),
.B2(n_28),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_73),
.A2(n_83),
.B1(n_91),
.B2(n_97),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_22),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_75),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_37),
.Y(n_76)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_34),
.B1(n_30),
.B2(n_33),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_78),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_110)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_86),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_25),
.Y(n_82)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_51),
.A2(n_30),
.B1(n_29),
.B2(n_20),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_93),
.Y(n_124)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_47),
.A2(n_29),
.B1(n_20),
.B2(n_24),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_43),
.B(n_24),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_96),
.Y(n_120)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_43),
.B(n_35),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_95),
.Y(n_131)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_42),
.A2(n_32),
.B(n_31),
.C(n_27),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_56),
.A2(n_24),
.B1(n_31),
.B2(n_27),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_40),
.B(n_32),
.Y(n_98)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_40),
.B(n_21),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_21),
.C(n_3),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_41),
.B(n_26),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_100),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_41),
.B(n_26),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_102),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_108),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_117),
.B1(n_125),
.B2(n_128),
.Y(n_138)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_113),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_110),
.A2(n_62),
.B1(n_84),
.B2(n_92),
.Y(n_141)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_116),
.B(n_118),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_59),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_96),
.A2(n_16),
.B1(n_7),
.B2(n_9),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_2),
.C(n_7),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_11),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_86),
.A2(n_9),
.B1(n_11),
.B2(n_13),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_66),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_133),
.B(n_60),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_79),
.A2(n_11),
.B1(n_13),
.B2(n_15),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

NAND2xp33_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_94),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_135),
.B(n_153),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_133),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_104),
.B(n_99),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_139),
.Y(n_171)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_141),
.A2(n_147),
.B1(n_151),
.B2(n_154),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_130),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_144),
.Y(n_176)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_115),
.B(n_113),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_145),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_80),
.B1(n_101),
.B2(n_94),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_152),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_SL g149 ( 
.A(n_120),
.B(n_60),
.C(n_65),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_149),
.A2(n_131),
.B(n_107),
.Y(n_183)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_112),
.A2(n_80),
.B1(n_101),
.B2(n_90),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_121),
.A2(n_64),
.B(n_70),
.C(n_67),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_121),
.A2(n_79),
.B1(n_90),
.B2(n_95),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_13),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_156),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_15),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_158),
.Y(n_191)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_114),
.A2(n_93),
.B1(n_65),
.B2(n_74),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_164),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_16),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_166),
.Y(n_170)
);

AND2x2_ASAP7_75t_SL g163 ( 
.A(n_114),
.B(n_71),
.Y(n_163)
);

A2O1A1O1Ixp25_ASAP7_75t_L g186 ( 
.A1(n_163),
.A2(n_150),
.B(n_146),
.C(n_106),
.D(n_153),
.Y(n_186)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_108),
.B(n_16),
.Y(n_166)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_159),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_169),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_140),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_173),
.B(n_174),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_178),
.B(n_179),
.Y(n_213)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_74),
.B1(n_85),
.B2(n_109),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_157),
.B1(n_152),
.B2(n_144),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_139),
.B(n_128),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_185),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_183),
.A2(n_184),
.B(n_166),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_SL g184 ( 
.A1(n_163),
.A2(n_117),
.B(n_149),
.C(n_165),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_136),
.B(n_105),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_186),
.A2(n_111),
.B(n_122),
.Y(n_214)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_187),
.B(n_194),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_105),
.Y(n_188)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_188),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_126),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_192),
.C(n_196),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_143),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_190),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_138),
.B(n_129),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_146),
.B(n_129),
.Y(n_193)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_193),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_154),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_138),
.B(n_127),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_174),
.A2(n_162),
.B1(n_165),
.B2(n_158),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_197),
.A2(n_210),
.B1(n_184),
.B2(n_173),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_198),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_176),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_199),
.B(n_212),
.Y(n_232)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_218),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_202),
.A2(n_204),
.B(n_184),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_183),
.A2(n_148),
.B(n_127),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_184),
.A2(n_142),
.B(n_103),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_207),
.A2(n_177),
.B(n_195),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_194),
.A2(n_85),
.B1(n_159),
.B2(n_88),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_184),
.A2(n_103),
.B1(n_111),
.B2(n_122),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_211),
.A2(n_175),
.B1(n_171),
.B2(n_178),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_214),
.A2(n_215),
.B(n_193),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_167),
.A2(n_88),
.B1(n_142),
.B2(n_123),
.Y(n_215)
);

MAJx2_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_132),
.C(n_89),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_189),
.C(n_196),
.Y(n_221)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_185),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_190),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_228),
.C(n_229),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_205),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_222),
.B(n_223),
.Y(n_240)
);

NAND3xp33_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_175),
.C(n_217),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_224),
.A2(n_225),
.B(n_227),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_226),
.B(n_233),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_202),
.A2(n_177),
.B(n_167),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_192),
.C(n_188),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_172),
.C(n_170),
.Y(n_229)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_182),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_214),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_235),
.B(n_238),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_172),
.C(n_170),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_200),
.C(n_216),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_237),
.A2(n_212),
.B1(n_197),
.B2(n_203),
.Y(n_249)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_206),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_225),
.A2(n_209),
.B1(n_207),
.B2(n_200),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_250),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_218),
.Y(n_245)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_245),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_227),
.C(n_230),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_221),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_252),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_236),
.A2(n_210),
.B1(n_215),
.B2(n_199),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_231),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_232),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_222),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_238),
.Y(n_254)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_257),
.C(n_261),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_229),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_260),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_241),
.A2(n_224),
.B(n_232),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_228),
.Y(n_261)
);

OA21x2_ASAP7_75t_SL g263 ( 
.A1(n_240),
.A2(n_226),
.B(n_234),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_263),
.B(n_246),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_244),
.C(n_242),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_208),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_265),
.B(n_266),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_255),
.A2(n_251),
.B1(n_258),
.B2(n_239),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_271),
.C(n_272),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_254),
.B(n_219),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_264),
.B(n_252),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_273),
.A2(n_245),
.B(n_168),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_269),
.A2(n_260),
.B(n_268),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_274),
.A2(n_277),
.B(n_243),
.Y(n_280)
);

AOI31xp67_ASAP7_75t_SL g276 ( 
.A1(n_271),
.A2(n_237),
.A3(n_250),
.B(n_247),
.Y(n_276)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_276),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_256),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_261),
.C(n_213),
.Y(n_281)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_280),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_281),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_279),
.A2(n_168),
.B(n_187),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_278),
.C(n_282),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_286),
.B(n_287),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_283),
.C(n_275),
.Y(n_287)
);


endmodule