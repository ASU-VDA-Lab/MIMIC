module real_aes_453_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_0), .B(n_504), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_1), .A2(n_506), .B(n_507), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_2), .B(n_830), .Y(n_829) );
AOI22xp5_ASAP7_75t_L g792 ( .A1(n_3), .A2(n_4), .B1(n_793), .B2(n_794), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_3), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_4), .Y(n_793) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_5), .B(n_221), .Y(n_541) );
INVx1_ASAP7_75t_L g153 ( .A(n_6), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_7), .B(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_8), .B(n_221), .Y(n_590) );
INVx1_ASAP7_75t_L g191 ( .A(n_9), .Y(n_191) );
CKINVDCx16_ASAP7_75t_R g830 ( .A(n_10), .Y(n_830) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_11), .Y(n_159) );
NAND2xp33_ASAP7_75t_L g582 ( .A(n_12), .B(n_218), .Y(n_582) );
INVx2_ASAP7_75t_L g135 ( .A(n_13), .Y(n_135) );
AOI221x1_ASAP7_75t_L g526 ( .A1(n_14), .A2(n_28), .B1(n_504), .B2(n_506), .C(n_527), .Y(n_526) );
OAI22xp5_ASAP7_75t_SL g790 ( .A1(n_15), .A2(n_791), .B1(n_792), .B2(n_795), .Y(n_790) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_15), .Y(n_795) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_16), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_17), .B(n_504), .Y(n_578) );
INVx1_ASAP7_75t_L g219 ( .A(n_18), .Y(n_219) );
AO21x2_ASAP7_75t_L g576 ( .A1(n_19), .A2(n_188), .B(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_20), .B(n_183), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_21), .A2(n_82), .B1(n_820), .B2(n_821), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_21), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_22), .B(n_221), .Y(n_515) );
AO21x1_ASAP7_75t_L g536 ( .A1(n_23), .A2(n_504), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g119 ( .A(n_24), .Y(n_119) );
INVx1_ASAP7_75t_L g216 ( .A(n_25), .Y(n_216) );
INVx1_ASAP7_75t_SL g203 ( .A(n_26), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_27), .B(n_146), .Y(n_261) );
AOI33xp33_ASAP7_75t_L g241 ( .A1(n_29), .A2(n_54), .A3(n_139), .B1(n_164), .B2(n_242), .B3(n_243), .Y(n_241) );
NAND2x1_ASAP7_75t_L g557 ( .A(n_30), .B(n_221), .Y(n_557) );
NAND2x1_ASAP7_75t_L g589 ( .A(n_31), .B(n_218), .Y(n_589) );
INVx1_ASAP7_75t_L g144 ( .A(n_32), .Y(n_144) );
OA21x2_ASAP7_75t_L g134 ( .A1(n_33), .A2(n_89), .B(n_135), .Y(n_134) );
OR2x2_ASAP7_75t_L g185 ( .A(n_33), .B(n_89), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_34), .B(n_168), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_35), .B(n_218), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_36), .B(n_221), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_37), .B(n_218), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_38), .A2(n_506), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g152 ( .A(n_39), .B(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g163 ( .A(n_39), .Y(n_163) );
AND2x2_ASAP7_75t_L g172 ( .A(n_39), .B(n_142), .Y(n_172) );
OR2x6_ASAP7_75t_L g117 ( .A(n_40), .B(n_118), .Y(n_117) );
NOR3xp33_ASAP7_75t_L g828 ( .A(n_40), .B(n_115), .C(n_829), .Y(n_828) );
CKINVDCx20_ASAP7_75t_R g154 ( .A(n_41), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_42), .B(n_504), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_43), .B(n_168), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g254 ( .A1(n_44), .A2(n_133), .B1(n_210), .B2(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_45), .B(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_46), .B(n_146), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_47), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_48), .B(n_218), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_49), .B(n_188), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_50), .B(n_146), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_51), .A2(n_506), .B(n_588), .Y(n_587) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_52), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_53), .B(n_218), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_55), .B(n_146), .Y(n_180) );
INVx1_ASAP7_75t_L g140 ( .A(n_56), .Y(n_140) );
INVx1_ASAP7_75t_L g148 ( .A(n_56), .Y(n_148) );
AND2x2_ASAP7_75t_L g182 ( .A(n_57), .B(n_183), .Y(n_182) );
AOI221xp5_ASAP7_75t_L g189 ( .A1(n_58), .A2(n_77), .B1(n_161), .B2(n_168), .C(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_59), .B(n_168), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_60), .B(n_221), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_61), .B(n_133), .Y(n_166) );
AOI21xp5_ASAP7_75t_SL g228 ( .A1(n_62), .A2(n_161), .B(n_229), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_63), .A2(n_506), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g213 ( .A(n_64), .Y(n_213) );
AO21x1_ASAP7_75t_L g538 ( .A1(n_65), .A2(n_506), .B(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_66), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g179 ( .A(n_67), .Y(n_179) );
XNOR2x1_ASAP7_75t_L g817 ( .A(n_68), .B(n_818), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_69), .A2(n_104), .B1(n_822), .B2(n_831), .Y(n_103) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_70), .B(n_504), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_71), .A2(n_161), .B(n_178), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_72), .Y(n_797) );
AND2x2_ASAP7_75t_L g551 ( .A(n_73), .B(n_184), .Y(n_551) );
INVx1_ASAP7_75t_L g142 ( .A(n_74), .Y(n_142) );
INVx1_ASAP7_75t_L g150 ( .A(n_74), .Y(n_150) );
AND2x2_ASAP7_75t_L g592 ( .A(n_75), .B(n_132), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_76), .B(n_168), .Y(n_244) );
AND2x2_ASAP7_75t_L g205 ( .A(n_78), .B(n_132), .Y(n_205) );
INVx1_ASAP7_75t_L g214 ( .A(n_79), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_80), .A2(n_161), .B(n_202), .Y(n_201) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_81), .A2(n_161), .B(n_236), .C(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g821 ( .A(n_82), .Y(n_821) );
INVx1_ASAP7_75t_L g120 ( .A(n_83), .Y(n_120) );
AND2x2_ASAP7_75t_L g501 ( .A(n_84), .B(n_132), .Y(n_501) );
AND2x2_ASAP7_75t_SL g226 ( .A(n_85), .B(n_132), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_86), .B(n_504), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_87), .A2(n_161), .B1(n_239), .B2(n_240), .Y(n_238) );
AND2x2_ASAP7_75t_L g537 ( .A(n_88), .B(n_210), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_90), .B(n_218), .Y(n_516) );
AND2x2_ASAP7_75t_L g560 ( .A(n_91), .B(n_132), .Y(n_560) );
INVx1_ASAP7_75t_L g230 ( .A(n_92), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_93), .B(n_221), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_94), .A2(n_506), .B(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_95), .B(n_218), .Y(n_528) );
AND2x2_ASAP7_75t_L g245 ( .A(n_96), .B(n_132), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_97), .B(n_221), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g136 ( .A1(n_98), .A2(n_137), .B(n_143), .C(n_151), .Y(n_136) );
BUFx2_ASAP7_75t_L g109 ( .A(n_99), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_100), .A2(n_506), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_101), .B(n_146), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_102), .B(n_112), .Y(n_111) );
AO22x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_110), .B1(n_810), .B2(n_812), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
BUFx3_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
HB1xp67_ASAP7_75t_L g811 ( .A(n_108), .Y(n_811) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_111), .B(n_121), .C(n_801), .Y(n_110) );
OAI21x1_ASAP7_75t_SL g812 ( .A1(n_111), .A2(n_813), .B(n_817), .Y(n_812) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_R g816 ( .A(n_114), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
OR2x6_ASAP7_75t_SL g492 ( .A(n_115), .B(n_116), .Y(n_492) );
AND2x6_ASAP7_75t_SL g789 ( .A(n_115), .B(n_117), .Y(n_789) );
OR2x2_ASAP7_75t_L g800 ( .A(n_115), .B(n_117), .Y(n_800) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g827 ( .A(n_119), .B(n_120), .Y(n_827) );
AOI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_790), .B(n_796), .Y(n_121) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_490), .B1(n_493), .B2(n_788), .Y(n_122) );
INVxp67_ASAP7_75t_SL g803 ( .A(n_123), .Y(n_803) );
NAND3x1_ASAP7_75t_L g123 ( .A(n_124), .B(n_369), .C(n_436), .Y(n_123) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_329), .Y(n_124) );
NOR3x1_ASAP7_75t_L g125 ( .A(n_126), .B(n_280), .C(n_309), .Y(n_125) );
OAI221xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_194), .B1(n_233), .B2(n_248), .C(n_265), .Y(n_126) );
A2O1A1Ixp33_ASAP7_75t_SL g443 ( .A1(n_127), .A2(n_207), .B(n_444), .C(n_445), .Y(n_443) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_128), .A2(n_415), .B1(n_418), .B2(n_420), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_128), .B(n_234), .Y(n_489) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_173), .Y(n_128) );
BUFx2_ASAP7_75t_L g408 ( .A(n_129), .Y(n_408) );
INVx1_ASAP7_75t_SL g421 ( .A(n_129), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_129), .B(n_276), .Y(n_463) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x4_ASAP7_75t_L g246 ( .A(n_130), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g291 ( .A(n_130), .B(n_187), .Y(n_291) );
INVx1_ASAP7_75t_L g302 ( .A(n_130), .Y(n_302) );
INVx2_ASAP7_75t_L g306 ( .A(n_130), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_130), .B(n_277), .Y(n_433) );
OR2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_156), .Y(n_130) );
OAI22xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_136), .B1(n_154), .B2(n_155), .Y(n_131) );
INVx3_ASAP7_75t_L g155 ( .A(n_132), .Y(n_155) );
INVx4_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_133), .B(n_158), .Y(n_157) );
INVx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
BUFx4f_ASAP7_75t_L g188 ( .A(n_134), .Y(n_188) );
AND2x2_ASAP7_75t_SL g184 ( .A(n_135), .B(n_185), .Y(n_184) );
AND2x4_ASAP7_75t_L g210 ( .A(n_135), .B(n_185), .Y(n_210) );
INVxp67_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
O2A1O1Ixp33_ASAP7_75t_L g178 ( .A1(n_138), .A2(n_179), .B(n_180), .C(n_181), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_SL g190 ( .A1(n_138), .A2(n_181), .B(n_191), .C(n_192), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_SL g202 ( .A1(n_138), .A2(n_181), .B(n_203), .C(n_204), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g212 ( .A1(n_138), .A2(n_145), .B1(n_213), .B2(n_214), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_138), .A2(n_181), .B(n_230), .C(n_231), .Y(n_229) );
INVx2_ASAP7_75t_L g263 ( .A(n_138), .Y(n_263) );
OR2x6_ASAP7_75t_L g138 ( .A(n_139), .B(n_141), .Y(n_138) );
AND2x2_ASAP7_75t_L g169 ( .A(n_139), .B(n_170), .Y(n_169) );
INVxp33_ASAP7_75t_L g242 ( .A(n_139), .Y(n_242) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g165 ( .A(n_140), .B(n_153), .Y(n_165) );
AND2x4_ASAP7_75t_L g221 ( .A(n_140), .B(n_149), .Y(n_221) );
INVx3_ASAP7_75t_L g164 ( .A(n_141), .Y(n_164) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x6_ASAP7_75t_L g218 ( .A(n_142), .B(n_147), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x4_ASAP7_75t_L g504 ( .A(n_146), .B(n_152), .Y(n_504) );
AND2x4_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
HB1xp67_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx5_ASAP7_75t_L g181 ( .A(n_152), .Y(n_181) );
HB1xp67_ASAP7_75t_L g170 ( .A(n_153), .Y(n_170) );
AO21x2_ASAP7_75t_L g174 ( .A1(n_155), .A2(n_175), .B(n_182), .Y(n_174) );
AO21x2_ASAP7_75t_L g277 ( .A1(n_155), .A2(n_175), .B(n_182), .Y(n_277) );
AO21x2_ASAP7_75t_L g544 ( .A1(n_155), .A2(n_545), .B(n_551), .Y(n_544) );
AO21x2_ASAP7_75t_L g553 ( .A1(n_155), .A2(n_554), .B(n_560), .Y(n_553) );
AO21x2_ASAP7_75t_L g566 ( .A1(n_155), .A2(n_554), .B(n_560), .Y(n_566) );
AO21x2_ASAP7_75t_L g569 ( .A1(n_155), .A2(n_545), .B(n_551), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_160), .B1(n_166), .B2(n_167), .Y(n_156) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVxp67_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_162), .B(n_165), .Y(n_161) );
NOR2x1p5_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
INVx1_ASAP7_75t_L g243 ( .A(n_164), .Y(n_243) );
AND2x6_ASAP7_75t_L g506 ( .A(n_165), .B(n_172), .Y(n_506) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_169), .B(n_171), .Y(n_168) );
INVx1_ASAP7_75t_L g256 ( .A(n_169), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_171), .Y(n_257) );
BUFx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AND2x2_ASAP7_75t_L g382 ( .A(n_173), .B(n_383), .Y(n_382) );
NOR2x1_ASAP7_75t_L g173 ( .A(n_174), .B(n_186), .Y(n_173) );
INVx2_ASAP7_75t_L g285 ( .A(n_174), .Y(n_285) );
AND2x2_ASAP7_75t_L g305 ( .A(n_174), .B(n_306), .Y(n_305) );
NOR2xp67_ASAP7_75t_L g430 ( .A(n_174), .B(n_306), .Y(n_430) );
AND2x2_ASAP7_75t_L g455 ( .A(n_174), .B(n_298), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_181), .B(n_210), .Y(n_222) );
INVx1_ASAP7_75t_L g239 ( .A(n_181), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_181), .A2(n_261), .B(n_262), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_181), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_181), .A2(n_515), .B(n_516), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_181), .A2(n_528), .B(n_529), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_181), .A2(n_540), .B(n_541), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_181), .A2(n_548), .B(n_549), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_181), .A2(n_557), .B(n_558), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_181), .A2(n_581), .B(n_582), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_181), .A2(n_589), .B(n_590), .Y(n_588) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_183), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_183), .A2(n_503), .B(n_505), .Y(n_502) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_183), .A2(n_526), .B(n_530), .Y(n_525) );
OA21x2_ASAP7_75t_L g596 ( .A1(n_183), .A2(n_526), .B(n_530), .Y(n_596) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g247 ( .A(n_187), .Y(n_247) );
INVx1_ASAP7_75t_L g269 ( .A(n_187), .Y(n_269) );
INVxp67_ASAP7_75t_L g308 ( .A(n_187), .Y(n_308) );
AND2x4_ASAP7_75t_L g348 ( .A(n_187), .B(n_349), .Y(n_348) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_187), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_187), .B(n_299), .Y(n_434) );
OA21x2_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_193), .Y(n_187) );
INVx2_ASAP7_75t_SL g236 ( .A(n_188), .Y(n_236) );
INVx1_ASAP7_75t_SL g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_206), .Y(n_195) );
AND2x2_ASAP7_75t_L g322 ( .A(n_196), .B(n_294), .Y(n_322) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_197), .Y(n_250) );
AND2x2_ASAP7_75t_L g278 ( .A(n_197), .B(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g289 ( .A(n_197), .Y(n_289) );
INVx1_ASAP7_75t_L g313 ( .A(n_197), .Y(n_313) );
AND2x2_ASAP7_75t_L g316 ( .A(n_197), .B(n_208), .Y(n_316) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_197), .Y(n_338) );
AO21x2_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_205), .Y(n_197) );
AO21x2_ASAP7_75t_L g585 ( .A1(n_198), .A2(n_586), .B(n_592), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
NOR2x1_ASAP7_75t_L g206 ( .A(n_207), .B(n_223), .Y(n_206) );
AND2x2_ASAP7_75t_L g303 ( .A(n_207), .B(n_225), .Y(n_303) );
NAND2x1_ASAP7_75t_L g336 ( .A(n_207), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g439 ( .A(n_207), .Y(n_439) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx3_ASAP7_75t_L g279 ( .A(n_208), .Y(n_279) );
AND2x2_ASAP7_75t_L g294 ( .A(n_208), .B(n_253), .Y(n_294) );
NOR2x1_ASAP7_75t_SL g363 ( .A(n_208), .B(n_225), .Y(n_363) );
AND2x4_ASAP7_75t_L g208 ( .A(n_209), .B(n_211), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_210), .A2(n_228), .B(n_232), .Y(n_227) );
INVx1_ASAP7_75t_SL g511 ( .A(n_210), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_210), .B(n_543), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_210), .A2(n_578), .B(n_579), .Y(n_577) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_215), .B(n_222), .Y(n_211) );
OAI22xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B1(n_219), .B2(n_220), .Y(n_215) );
INVxp67_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVxp67_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
NOR2x1_ASAP7_75t_L g400 ( .A(n_223), .B(n_387), .Y(n_400) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g325 ( .A(n_224), .B(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx4_ASAP7_75t_L g264 ( .A(n_225), .Y(n_264) );
AND2x4_ASAP7_75t_L g271 ( .A(n_225), .B(n_272), .Y(n_271) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_225), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_225), .B(n_288), .Y(n_388) );
AND2x2_ASAP7_75t_L g416 ( .A(n_225), .B(n_253), .Y(n_416) );
OR2x6_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
NAND2x1_ASAP7_75t_SL g233 ( .A(n_234), .B(n_246), .Y(n_233) );
OR2x2_ASAP7_75t_L g444 ( .A(n_234), .B(n_356), .Y(n_444) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x4_ASAP7_75t_L g284 ( .A(n_235), .B(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g349 ( .A(n_235), .Y(n_349) );
AND2x2_ASAP7_75t_L g383 ( .A(n_235), .B(n_306), .Y(n_383) );
AO21x2_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_245), .Y(n_235) );
AO21x2_ASAP7_75t_L g299 ( .A1(n_236), .A2(n_237), .B(n_245), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_238), .B(n_244), .Y(n_237) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx3_ASAP7_75t_L g356 ( .A(n_246), .Y(n_356) );
AND2x2_ASAP7_75t_L g364 ( .A(n_246), .B(n_297), .Y(n_364) );
AND2x2_ASAP7_75t_L g481 ( .A(n_246), .B(n_284), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_249), .B(n_251), .Y(n_248) );
BUFx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g435 ( .A(n_250), .B(n_376), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_250), .B(n_275), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_251), .A2(n_312), .B(n_315), .Y(n_311) );
AND2x2_ASAP7_75t_L g381 ( .A(n_251), .B(n_287), .Y(n_381) );
INVx2_ASAP7_75t_SL g468 ( .A(n_251), .Y(n_468) );
AND2x4_ASAP7_75t_SL g251 ( .A(n_252), .B(n_264), .Y(n_251) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g272 ( .A(n_253), .Y(n_272) );
INVx2_ASAP7_75t_L g319 ( .A(n_253), .Y(n_319) );
AND2x4_ASAP7_75t_L g326 ( .A(n_253), .B(n_279), .Y(n_326) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_259), .Y(n_253) );
NOR3xp33_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .C(n_258), .Y(n_255) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_264), .Y(n_282) );
AND2x4_ASAP7_75t_L g358 ( .A(n_264), .B(n_272), .Y(n_358) );
OR2x2_ASAP7_75t_L g484 ( .A(n_264), .B(n_485), .Y(n_484) );
NAND4xp25_ASAP7_75t_L g265 ( .A(n_266), .B(n_270), .C(n_273), .D(n_278), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g331 ( .A(n_267), .B(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g428 ( .A(n_267), .Y(n_428) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2x1p5_ASAP7_75t_L g328 ( .A(n_268), .B(n_276), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_268), .B(n_333), .Y(n_462) );
BUFx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_271), .B(n_287), .Y(n_340) );
INVx2_ASAP7_75t_L g442 ( .A(n_271), .Y(n_442) );
AND2x2_ASAP7_75t_SL g452 ( .A(n_271), .B(n_312), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_271), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g344 ( .A(n_275), .B(n_291), .Y(n_344) );
AND2x2_ASAP7_75t_L g412 ( .A(n_275), .B(n_348), .Y(n_412) );
INVx3_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x4_ASAP7_75t_L g297 ( .A(n_276), .B(n_298), .Y(n_297) );
INVx3_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_277), .Y(n_351) );
AND2x2_ASAP7_75t_L g402 ( .A(n_277), .B(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_277), .B(n_299), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_278), .B(n_442), .Y(n_449) );
INVx1_ASAP7_75t_SL g485 ( .A(n_278), .Y(n_485) );
INVx1_ASAP7_75t_L g314 ( .A(n_279), .Y(n_314) );
AND2x2_ASAP7_75t_L g376 ( .A(n_279), .B(n_319), .Y(n_376) );
OAI21xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_290), .B(n_292), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
AND2x2_ASAP7_75t_L g342 ( .A(n_284), .B(n_291), .Y(n_342) );
AND2x2_ASAP7_75t_L g450 ( .A(n_284), .B(n_301), .Y(n_450) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g324 ( .A(n_287), .Y(n_324) );
AND2x2_ASAP7_75t_L g357 ( .A(n_287), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g362 ( .A(n_287), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_287), .B(n_326), .Y(n_411) );
NOR3xp33_ASAP7_75t_L g461 ( .A(n_287), .B(n_462), .C(n_463), .Y(n_461) );
INVx3_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVxp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_296), .B1(n_303), .B2(n_304), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
INVx2_ASAP7_75t_L g387 ( .A(n_294), .Y(n_387) );
AND2x2_ASAP7_75t_L g321 ( .A(n_295), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g343 ( .A(n_295), .B(n_316), .Y(n_343) );
AND2x2_ASAP7_75t_SL g375 ( .A(n_295), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_300), .Y(n_296) );
INVx1_ASAP7_75t_L g354 ( .A(n_297), .Y(n_354) );
AND2x2_ASAP7_75t_L g307 ( .A(n_298), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g333 ( .A(n_298), .Y(n_333) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g396 ( .A(n_302), .B(n_348), .Y(n_396) );
INVx1_ASAP7_75t_L g454 ( .A(n_302), .Y(n_454) );
INVx1_ASAP7_75t_L g310 ( .A(n_304), .Y(n_310) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
NAND2x1p5_ASAP7_75t_L g332 ( .A(n_305), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g441 ( .A(n_305), .B(n_348), .Y(n_441) );
AND2x2_ASAP7_75t_L g407 ( .A(n_307), .B(n_408), .Y(n_407) );
NAND2x1p5_ASAP7_75t_L g475 ( .A(n_307), .B(n_476), .Y(n_475) );
OAI21xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_311), .B(n_320), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_312), .B(n_347), .Y(n_346) );
AND2x4_ASAP7_75t_L g368 ( .A(n_312), .B(n_317), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_312), .B(n_358), .Y(n_419) );
AND2x4_ASAP7_75t_SL g312 ( .A(n_313), .B(n_314), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_313), .B(n_376), .Y(n_406) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_313), .Y(n_426) );
AOI22xp5_ASAP7_75t_L g341 ( .A1(n_315), .A2(n_342), .B1(n_343), .B2(n_344), .Y(n_341) );
AND2x2_ASAP7_75t_SL g315 ( .A(n_316), .B(n_317), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_316), .B(n_358), .Y(n_377) );
INVx1_ASAP7_75t_L g478 ( .A(n_316), .Y(n_478) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OAI21xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_323), .B(n_327), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_322), .B(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g459 ( .A(n_325), .Y(n_459) );
INVx4_ASAP7_75t_L g361 ( .A(n_326), .Y(n_361) );
INVxp33_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g389 ( .A(n_328), .B(n_390), .Y(n_389) );
NOR2x1_ASAP7_75t_L g329 ( .A(n_330), .B(n_345), .Y(n_329) );
OAI21xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_334), .B(n_341), .Y(n_330) );
INVx1_ASAP7_75t_L g379 ( .A(n_332), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_335), .B(n_339), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g384 ( .A(n_336), .Y(n_384) );
INVx1_ASAP7_75t_L g417 ( .A(n_337), .Y(n_417) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_342), .A2(n_381), .B1(n_382), .B2(n_384), .Y(n_380) );
INVx1_ASAP7_75t_L g394 ( .A(n_343), .Y(n_394) );
NAND4xp25_ASAP7_75t_SL g345 ( .A(n_346), .B(n_352), .C(n_359), .D(n_365), .Y(n_345) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
INVx1_ASAP7_75t_L g367 ( .A(n_348), .Y(n_367) );
AND2x2_ASAP7_75t_L g479 ( .A(n_348), .B(n_476), .Y(n_479) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_357), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g486 ( .A(n_356), .B(n_423), .Y(n_486) );
INVx1_ASAP7_75t_L g483 ( .A(n_357), .Y(n_483) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_358), .Y(n_392) );
OAI21xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_362), .B(n_364), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_368), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_397), .Y(n_369) );
NOR3xp33_ASAP7_75t_L g370 ( .A(n_371), .B(n_385), .C(n_393), .Y(n_370) );
OAI21xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_378), .B(n_380), .Y(n_371) );
INVxp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_377), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_375), .A2(n_407), .B1(n_410), .B2(n_412), .Y(n_409) );
OAI22xp33_ASAP7_75t_L g385 ( .A1(n_378), .A2(n_386), .B1(n_389), .B2(n_391), .Y(n_385) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g390 ( .A(n_383), .Y(n_390) );
AND2x4_ASAP7_75t_L g401 ( .A(n_383), .B(n_402), .Y(n_401) );
OR2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_388), .Y(n_488) );
AOI31xp33_ASAP7_75t_L g487 ( .A1(n_391), .A2(n_464), .A3(n_488), .B(n_489), .Y(n_487) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_398), .B(n_413), .Y(n_397) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_399), .B(n_409), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B1(n_404), .B2(n_407), .Y(n_399) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_403), .Y(n_467) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_411), .B(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_414), .B(n_424), .Y(n_413) );
AND2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
AND2x2_ASAP7_75t_L g425 ( .A(n_416), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g464 ( .A(n_416), .Y(n_464) );
AOI22xp33_ASAP7_75t_SL g473 ( .A1(n_416), .A2(n_474), .B1(n_477), .B2(n_479), .Y(n_473) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_421), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_427), .B1(n_431), .B2(n_435), .Y(n_424) );
NOR2xp33_ASAP7_75t_SL g427 ( .A(n_428), .B(n_429), .Y(n_427) );
INVxp67_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
INVx2_ASAP7_75t_SL g476 ( .A(n_433), .Y(n_476) );
INVx2_ASAP7_75t_L g457 ( .A(n_434), .Y(n_457) );
AND2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_471), .Y(n_436) );
AOI211xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_443), .B(n_446), .C(n_460), .Y(n_437) );
OAI21xp33_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_440), .B(n_442), .Y(n_438) );
INVx1_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g445 ( .A(n_442), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g446 ( .A(n_447), .B(n_451), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_450), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B1(n_456), .B2(n_458), .Y(n_451) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
AND2x2_ASAP7_75t_L g456 ( .A(n_454), .B(n_457), .Y(n_456) );
AO22x1_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_464), .B1(n_465), .B2(n_469), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_468), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NOR3xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_482), .C(n_487), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_473), .B(n_480), .Y(n_472) );
INVx3_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AOI21xp33_ASAP7_75t_R g482 ( .A1(n_483), .A2(n_484), .B(n_486), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_491), .Y(n_490) );
CKINVDCx5p33_ASAP7_75t_R g804 ( .A(n_491), .Y(n_804) );
CKINVDCx11_ASAP7_75t_R g491 ( .A(n_492), .Y(n_491) );
XOR2x2_ASAP7_75t_L g818 ( .A(n_493), .B(n_819), .Y(n_818) );
INVx3_ASAP7_75t_SL g493 ( .A(n_494), .Y(n_493) );
BUFx2_ASAP7_75t_L g805 ( .A(n_494), .Y(n_805) );
NOR2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_675), .Y(n_494) );
AO211x2_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_520), .B(n_570), .C(n_643), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVxp67_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
AND3x2_ASAP7_75t_L g724 ( .A(n_498), .B(n_605), .C(n_621), .Y(n_724) );
AND2x4_ASAP7_75t_L g727 ( .A(n_498), .B(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_510), .Y(n_498) );
NAND2x1p5_ASAP7_75t_L g583 ( .A(n_499), .B(n_584), .Y(n_583) );
INVx4_ASAP7_75t_L g636 ( .A(n_499), .Y(n_636) );
AND2x2_ASAP7_75t_SL g721 ( .A(n_499), .B(n_630), .Y(n_721) );
AND2x2_ASAP7_75t_L g764 ( .A(n_499), .B(n_585), .Y(n_764) );
INVx5_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx2_ASAP7_75t_L g613 ( .A(n_500), .Y(n_613) );
AND2x2_ASAP7_75t_L g632 ( .A(n_500), .B(n_576), .Y(n_632) );
AND2x2_ASAP7_75t_L g650 ( .A(n_500), .B(n_585), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_500), .B(n_584), .Y(n_710) );
NOR2x1_ASAP7_75t_SL g737 ( .A(n_500), .B(n_510), .Y(n_737) );
OR2x6_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_510), .B(n_576), .Y(n_575) );
AO21x2_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B(n_518), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_511), .B(n_519), .Y(n_518) );
AO21x2_ASAP7_75t_L g609 ( .A1(n_511), .A2(n_512), .B(n_518), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_517), .Y(n_512) );
AO21x1_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_552), .B(n_561), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OAI22xp33_ASAP7_75t_L g618 ( .A1(n_522), .A2(n_619), .B1(n_623), .B2(n_624), .Y(n_618) );
OR2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_531), .Y(n_522) );
AND2x2_ASAP7_75t_L g679 ( .A(n_523), .B(n_567), .Y(n_679) );
BUFx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x4_ASAP7_75t_L g612 ( .A(n_524), .B(n_595), .Y(n_612) );
AND2x2_ASAP7_75t_L g684 ( .A(n_524), .B(n_569), .Y(n_684) );
AND2x2_ASAP7_75t_L g703 ( .A(n_524), .B(n_669), .Y(n_703) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g562 ( .A(n_525), .Y(n_562) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_525), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_531), .B(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g663 ( .A(n_532), .B(n_564), .Y(n_663) );
AND2x4_ASAP7_75t_L g532 ( .A(n_533), .B(n_544), .Y(n_532) );
AND2x2_ASAP7_75t_L g567 ( .A(n_533), .B(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g600 ( .A(n_533), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_SL g660 ( .A(n_533), .B(n_596), .Y(n_660) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
BUFx2_ASAP7_75t_L g753 ( .A(n_534), .Y(n_753) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g595 ( .A(n_535), .Y(n_595) );
OAI21x1_ASAP7_75t_SL g535 ( .A1(n_536), .A2(n_538), .B(n_542), .Y(n_535) );
INVx1_ASAP7_75t_L g543 ( .A(n_537), .Y(n_543) );
INVx2_ASAP7_75t_L g601 ( .A(n_544), .Y(n_601) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_544), .Y(n_701) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_546), .B(n_550), .Y(n_545) );
INVx2_ASAP7_75t_L g597 ( .A(n_552), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_552), .B(n_729), .Y(n_755) );
AND2x2_ASAP7_75t_L g774 ( .A(n_552), .B(n_764), .Y(n_774) );
BUFx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x4_ASAP7_75t_SL g642 ( .A(n_553), .B(n_601), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_559), .Y(n_554) );
AND2x2_ASAP7_75t_SL g561 ( .A(n_562), .B(n_563), .Y(n_561) );
AND2x2_ASAP7_75t_L g641 ( .A(n_562), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_562), .B(n_611), .Y(n_646) );
INVx1_ASAP7_75t_SL g773 ( .A(n_562), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_563), .B(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_567), .Y(n_563) );
INVx1_ASAP7_75t_L g599 ( .A(n_564), .Y(n_599) );
AND2x2_ASAP7_75t_L g785 ( .A(n_564), .B(n_786), .Y(n_785) );
BUFx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g661 ( .A(n_565), .B(n_568), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_565), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g715 ( .A(n_565), .B(n_569), .Y(n_715) );
AND2x2_ASAP7_75t_L g746 ( .A(n_565), .B(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g611 ( .A(n_566), .B(n_569), .Y(n_611) );
INVxp67_ASAP7_75t_L g628 ( .A(n_566), .Y(n_628) );
BUFx3_ASAP7_75t_L g669 ( .A(n_566), .Y(n_669) );
AND2x2_ASAP7_75t_L g689 ( .A(n_567), .B(n_690), .Y(n_689) );
NAND2xp33_ASAP7_75t_L g702 ( .A(n_567), .B(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_568), .B(n_595), .Y(n_658) );
AND2x2_ASAP7_75t_L g747 ( .A(n_568), .B(n_596), .Y(n_747) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g674 ( .A(n_569), .B(n_596), .Y(n_674) );
OR3x1_ASAP7_75t_L g570 ( .A(n_571), .B(n_618), .C(n_633), .Y(n_570) );
OAI321xp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_583), .A3(n_593), .B1(n_598), .B2(n_602), .C(n_610), .Y(n_571) );
INVx1_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVxp67_ASAP7_75t_SL g649 ( .A(n_575), .Y(n_649) );
INVxp67_ASAP7_75t_SL g667 ( .A(n_575), .Y(n_667) );
OR2x2_ASAP7_75t_L g671 ( .A(n_575), .B(n_583), .Y(n_671) );
BUFx3_ASAP7_75t_L g605 ( .A(n_576), .Y(n_605) );
AND2x2_ASAP7_75t_L g622 ( .A(n_576), .B(n_608), .Y(n_622) );
INVx1_ASAP7_75t_L g639 ( .A(n_576), .Y(n_639) );
INVx2_ASAP7_75t_L g655 ( .A(n_576), .Y(n_655) );
OR2x2_ASAP7_75t_L g694 ( .A(n_576), .B(n_584), .Y(n_694) );
INVx2_ASAP7_75t_L g682 ( .A(n_583), .Y(n_682) );
AND2x2_ASAP7_75t_L g606 ( .A(n_584), .B(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g621 ( .A(n_584), .Y(n_621) );
AND2x4_ASAP7_75t_L g630 ( .A(n_584), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_584), .B(n_607), .Y(n_653) );
AND2x2_ASAP7_75t_L g760 ( .A(n_584), .B(n_655), .Y(n_760) );
INVx4_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_585), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_591), .Y(n_586) );
INVx1_ASAP7_75t_L g647 ( .A(n_593), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_594), .B(n_597), .Y(n_593) );
AND2x2_ASAP7_75t_L g734 ( .A(n_594), .B(n_661), .Y(n_734) );
INVx1_ASAP7_75t_SL g751 ( .A(n_594), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_594), .B(n_727), .Y(n_780) );
AND2x4_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
OR2x2_ASAP7_75t_L g623 ( .A(n_595), .B(n_596), .Y(n_623) );
AND2x2_ASAP7_75t_L g716 ( .A(n_597), .B(n_612), .Y(n_716) );
OR2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g739 ( .A(n_601), .B(n_612), .Y(n_739) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_603), .A2(n_752), .B1(n_757), .B2(n_759), .Y(n_756) );
AND2x4_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .Y(n_603) );
AND2x2_ASAP7_75t_L g681 ( .A(n_604), .B(n_682), .Y(n_681) );
OR2x2_ASAP7_75t_L g776 ( .A(n_604), .B(n_777), .Y(n_776) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g732 ( .A(n_605), .B(n_650), .Y(n_732) );
AND2x4_ASAP7_75t_L g686 ( .A(n_606), .B(n_632), .Y(n_686) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_608), .Y(n_784) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g617 ( .A(n_609), .Y(n_617) );
INVx1_ASAP7_75t_L g631 ( .A(n_609), .Y(n_631) );
NAND4xp25_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .C(n_613), .D(n_614), .Y(n_610) );
AND2x2_ASAP7_75t_L g768 ( .A(n_611), .B(n_753), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_611), .B(n_779), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_612), .B(n_688), .Y(n_687) );
OAI322xp33_ASAP7_75t_L g695 ( .A1(n_612), .A2(n_696), .A3(n_700), .B1(n_702), .B2(n_704), .C1(n_706), .C2(n_711), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_612), .B(n_661), .Y(n_711) );
INVx1_ASAP7_75t_L g779 ( .A(n_612), .Y(n_779) );
INVx2_ASAP7_75t_L g625 ( .A(n_613), .Y(n_625) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_616), .B(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_617), .B(n_636), .Y(n_693) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_620), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
INVx1_ASAP7_75t_L g666 ( .A(n_621), .Y(n_666) );
AND2x2_ASAP7_75t_L g738 ( .A(n_621), .B(n_649), .Y(n_738) );
AOI31xp33_ASAP7_75t_L g624 ( .A1(n_622), .A2(n_625), .A3(n_626), .B(n_629), .Y(n_624) );
AND2x2_ASAP7_75t_L g635 ( .A(n_622), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g763 ( .A(n_622), .B(n_764), .Y(n_763) );
AND2x2_ASAP7_75t_SL g770 ( .A(n_622), .B(n_650), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_622), .Y(n_771) );
INVx1_ASAP7_75t_SL g729 ( .A(n_623), .Y(n_729) );
NAND3xp33_ASAP7_75t_SL g757 ( .A(n_623), .B(n_751), .C(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g657 ( .A(n_628), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
AND2x2_ASAP7_75t_L g638 ( .A(n_630), .B(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g699 ( .A(n_630), .Y(n_699) );
AOI322xp5_ASAP7_75t_L g781 ( .A1(n_630), .A2(n_660), .A3(n_663), .B1(n_782), .B2(n_783), .C1(n_785), .C2(n_787), .Y(n_781) );
AND2x2_ASAP7_75t_L g787 ( .A(n_630), .B(n_636), .Y(n_787) );
AOI21xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_637), .B(n_640), .Y(n_633) );
INVx1_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_636), .B(n_655), .Y(n_654) );
AND2x4_ASAP7_75t_L g782 ( .A(n_636), .B(n_669), .Y(n_782) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g708 ( .A(n_639), .Y(n_708) );
AND2x2_ASAP7_75t_L g736 ( .A(n_639), .B(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g783 ( .A(n_639), .B(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g688 ( .A(n_642), .Y(n_688) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
O2A1O1Ixp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_647), .B(n_648), .C(n_651), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
AND2x2_ASAP7_75t_L g705 ( .A(n_650), .B(n_655), .Y(n_705) );
OAI211xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_656), .B(n_662), .C(n_664), .Y(n_651) );
OAI221xp5_ASAP7_75t_L g677 ( .A1(n_652), .A2(n_678), .B1(n_680), .B2(n_683), .C(n_685), .Y(n_677) );
OR2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx1_ASAP7_75t_L g697 ( .A(n_654), .Y(n_697) );
OR2x2_ASAP7_75t_L g717 ( .A(n_654), .B(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .Y(n_656) );
INVx1_ASAP7_75t_L g762 ( .A(n_657), .Y(n_762) );
INVx1_ASAP7_75t_L g786 ( .A(n_658), .Y(n_786) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_660), .B(n_661), .Y(n_659) );
AND2x2_ASAP7_75t_L g668 ( .A(n_660), .B(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_660), .B(n_730), .Y(n_742) );
INVx1_ASAP7_75t_L g722 ( .A(n_661), .Y(n_722) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_668), .B1(n_670), .B2(n_672), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
INVx1_ASAP7_75t_SL g730 ( .A(n_669), .Y(n_730) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NAND4xp75_ASAP7_75t_L g675 ( .A(n_676), .B(n_712), .C(n_740), .D(n_765), .Y(n_675) );
NOR2xp67_ASAP7_75t_L g676 ( .A(n_677), .B(n_695), .Y(n_676) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_SL g752 ( .A(n_684), .B(n_753), .Y(n_752) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_687), .B1(n_689), .B2(n_691), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_688), .B(n_751), .Y(n_750) );
INVx2_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
INVx2_ASAP7_75t_L g728 ( .A(n_694), .Y(n_728) );
OR2x2_ASAP7_75t_L g743 ( .A(n_694), .B(n_744), .Y(n_743) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_697), .B(n_698), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g758 ( .A(n_703), .Y(n_758) );
INVx1_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
OAI21xp5_ASAP7_75t_SL g749 ( .A1(n_705), .A2(n_750), .B(n_752), .Y(n_749) );
INVxp67_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
NOR2x1_ASAP7_75t_L g712 ( .A(n_713), .B(n_725), .Y(n_712) );
OAI221xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_717), .B1(n_720), .B2(n_722), .C(n_723), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
OAI21xp33_ASAP7_75t_L g761 ( .A1(n_715), .A2(n_762), .B(n_763), .Y(n_761) );
INVx3_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
OAI322xp33_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_729), .A3(n_730), .B1(n_731), .B2(n_733), .C1(n_735), .C2(n_739), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
NOR2x1_ASAP7_75t_L g735 ( .A(n_736), .B(n_738), .Y(n_735) );
INVx1_ASAP7_75t_L g748 ( .A(n_736), .Y(n_748) );
INVx1_ASAP7_75t_L g744 ( .A(n_737), .Y(n_744) );
AND2x2_ASAP7_75t_L g759 ( .A(n_737), .B(n_760), .Y(n_759) );
NOR2x1_ASAP7_75t_L g740 ( .A(n_741), .B(n_754), .Y(n_740) );
OAI221xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_743), .B1(n_745), .B2(n_748), .C(n_749), .Y(n_741) );
INVx1_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
OAI211xp5_ASAP7_75t_SL g754 ( .A1(n_748), .A2(n_755), .B(n_756), .C(n_761), .Y(n_754) );
INVx2_ASAP7_75t_SL g777 ( .A(n_764), .Y(n_777) );
NOR2x1_ASAP7_75t_L g765 ( .A(n_766), .B(n_775), .Y(n_765) );
OAI22xp33_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_769), .B1(n_771), .B2(n_772), .Y(n_766) );
INVx1_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_SL g769 ( .A(n_770), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .Y(n_772) );
OAI211xp5_ASAP7_75t_SL g775 ( .A1(n_776), .A2(n_778), .B(n_780), .C(n_781), .Y(n_775) );
CKINVDCx11_ASAP7_75t_R g788 ( .A(n_789), .Y(n_788) );
CKINVDCx5p33_ASAP7_75t_R g808 ( .A(n_789), .Y(n_808) );
INVxp33_ASAP7_75t_L g809 ( .A(n_790), .Y(n_809) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g796 ( .A(n_797), .B(n_798), .Y(n_796) );
INVx1_ASAP7_75t_SL g798 ( .A(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
NAND2xp5_ASAP7_75t_SL g801 ( .A(n_802), .B(n_809), .Y(n_801) );
OAI22x1_ASAP7_75t_L g802 ( .A1(n_803), .A2(n_804), .B1(n_805), .B2(n_806), .Y(n_802) );
CKINVDCx11_ASAP7_75t_R g806 ( .A(n_807), .Y(n_806) );
INVx3_ASAP7_75t_SL g807 ( .A(n_808), .Y(n_807) );
INVx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVxp67_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
CKINVDCx5p33_ASAP7_75t_R g822 ( .A(n_823), .Y(n_822) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_824), .Y(n_823) );
CKINVDCx5p33_ASAP7_75t_R g824 ( .A(n_825), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g832 ( .A(n_825), .Y(n_832) );
INVx3_ASAP7_75t_SL g825 ( .A(n_826), .Y(n_825) );
AND2x2_ASAP7_75t_SL g826 ( .A(n_827), .B(n_828), .Y(n_826) );
INVx1_ASAP7_75t_SL g831 ( .A(n_832), .Y(n_831) );
endmodule