module fake_jpeg_18229_n_155 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_155);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_155;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_28),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_5),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_14),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_4),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_26),
.B(n_0),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx6_ASAP7_75t_SL g77 ( 
.A(n_50),
.Y(n_77)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_80),
.A2(n_83),
.B1(n_60),
.B2(n_66),
.Y(n_86)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_82),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_86),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_60),
.B1(n_48),
.B2(n_64),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_87),
.A2(n_88),
.B1(n_89),
.B2(n_94),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_66),
.B1(n_75),
.B2(n_61),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_77),
.A2(n_71),
.B1(n_83),
.B2(n_78),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_81),
.B(n_58),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_65),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_80),
.A2(n_52),
.B1(n_57),
.B2(n_54),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_97),
.B(n_103),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_101),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_88),
.A2(n_84),
.B1(n_83),
.B2(n_90),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_100),
.A2(n_82),
.B1(n_62),
.B2(n_67),
.Y(n_112)
);

NOR2xp67_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_74),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_74),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_104),
.Y(n_110)
);

OR2x2_ASAP7_75t_SL g103 ( 
.A(n_93),
.B(n_69),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_84),
.B(n_49),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_55),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_108),
.Y(n_111)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_82),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_72),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g109 ( 
.A1(n_107),
.A2(n_90),
.B1(n_79),
.B2(n_82),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_109),
.A2(n_112),
.B1(n_118),
.B2(n_119),
.Y(n_136)
);

AND2x6_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_68),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_125),
.Y(n_128)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_107),
.A2(n_73),
.B1(n_59),
.B2(n_62),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_100),
.A2(n_108),
.B1(n_73),
.B2(n_98),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_62),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_122),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_53),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_20),
.B1(n_44),
.B2(n_40),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_1),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_124),
.Y(n_130)
);

AND2x6_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_19),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_21),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_131),
.C(n_110),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_16),
.C(n_38),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_2),
.B(n_3),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_133),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_120),
.B(n_2),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_3),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_4),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_126),
.A2(n_125),
.B(n_117),
.Y(n_137)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_138),
.A2(n_139),
.B1(n_141),
.B2(n_142),
.Y(n_143)
);

NAND2x1p5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_109),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_135),
.Y(n_141)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_143),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_139),
.B1(n_144),
.B2(n_136),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_129),
.C(n_144),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_147),
.A2(n_128),
.B1(n_138),
.B2(n_127),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_130),
.B1(n_140),
.B2(n_131),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_23),
.Y(n_150)
);

AOI322xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_114),
.A3(n_24),
.B1(n_27),
.B2(n_46),
.C1(n_37),
.C2(n_35),
.Y(n_151)
);

AOI322xp5_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_12),
.A3(n_32),
.B1(n_29),
.B2(n_22),
.C1(n_15),
.C2(n_34),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_6),
.Y(n_153)
);

AOI21x1_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_7),
.B(n_8),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_8),
.Y(n_155)
);


endmodule