module fake_jpeg_22545_n_134 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_134);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx3_ASAP7_75t_SL g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx8_ASAP7_75t_SL g22 ( 
.A(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_7),
.B(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_32),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_28),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_23),
.C(n_25),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_22),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_31),
.A2(n_17),
.B(n_20),
.Y(n_55)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_5),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_27),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_44),
.Y(n_68)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_59),
.B1(n_18),
.B2(n_7),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_52),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_51),
.B(n_63),
.Y(n_74)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_18),
.B(n_21),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_31),
.A2(n_18),
.B1(n_15),
.B2(n_20),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_18),
.B1(n_8),
.B2(n_10),
.Y(n_81)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_60),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_36),
.A2(n_14),
.B1(n_26),
.B2(n_24),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_32),
.B(n_15),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_64),
.Y(n_65)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_30),
.B(n_15),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_18),
.C(n_14),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_73),
.C(n_53),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_64),
.A2(n_15),
.B1(n_27),
.B2(n_26),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_67),
.A2(n_81),
.B1(n_13),
.B2(n_83),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_SL g92 ( 
.A(n_71),
.B(n_6),
.C(n_12),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_43),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g73 ( 
.A(n_50),
.B(n_21),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_51),
.B(n_19),
.Y(n_75)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_19),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_48),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_78),
.A2(n_79),
.B(n_52),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_55),
.A2(n_21),
.B(n_18),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_57),
.A2(n_18),
.B(n_21),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_80),
.A2(n_83),
.B(n_57),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_13),
.B(n_6),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_92),
.B1(n_66),
.B2(n_79),
.Y(n_103)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_47),
.Y(n_86)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_89),
.B(n_96),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_44),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_93),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_70),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_65),
.A2(n_48),
.B1(n_54),
.B2(n_49),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_94),
.A2(n_97),
.B1(n_74),
.B2(n_76),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_61),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_67),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_12),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_98),
.A2(n_105),
.B(n_93),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_88),
.A2(n_78),
.B1(n_80),
.B2(n_81),
.Y(n_101)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_103),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_90),
.Y(n_104)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_73),
.B(n_68),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_108),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_106),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_107),
.B(n_87),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_111),
.B(n_115),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_89),
.Y(n_115)
);

NAND2x1_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_96),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_116),
.B(n_101),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_118),
.C(n_110),
.Y(n_125)
);

OAI21x1_ASAP7_75t_L g119 ( 
.A1(n_116),
.A2(n_105),
.B(n_95),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_119),
.A2(n_109),
.B(n_113),
.Y(n_124)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_120),
.B(n_121),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_102),
.B1(n_104),
.B2(n_100),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_125),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_113),
.B(n_115),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_126),
.B(n_112),
.Y(n_129)
);

OAI221xp5_ASAP7_75t_L g127 ( 
.A1(n_118),
.A2(n_99),
.B1(n_112),
.B2(n_96),
.C(n_94),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_129),
.A2(n_123),
.B(n_99),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_132),
.C(n_130),
.Y(n_133)
);

OAI21x1_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_117),
.B(n_92),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_133),
.B(n_130),
.Y(n_134)
);


endmodule