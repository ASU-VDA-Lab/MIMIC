module fake_jpeg_28808_n_53 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_53);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_53;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_7),
.B(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_19),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_24),
.C(n_20),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_2),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_26),
.B(n_30),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_25),
.B(n_4),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_21),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_36),
.B(n_21),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_27),
.Y(n_36)
);

NAND2x1_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_34),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_38),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_33),
.A2(n_20),
.B(n_21),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_9),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_40),
.A2(n_37),
.B1(n_41),
.B2(n_7),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_38),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_47),
.B(n_49),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_42),
.A2(n_10),
.B1(n_14),
.B2(n_15),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_50),
.B(n_47),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_46),
.C(n_48),
.Y(n_52)
);

O2A1O1Ixp33_ASAP7_75t_SL g53 ( 
.A1(n_52),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_53)
);


endmodule