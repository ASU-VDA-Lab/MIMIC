module real_jpeg_5337_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_233;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_205;
wire n_110;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_244;
wire n_213;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_1),
.A2(n_45),
.B1(n_48),
.B2(n_49),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_1),
.A2(n_48),
.B1(n_54),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_1),
.A2(n_48),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_2),
.B(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_2),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_2),
.A2(n_100),
.B1(n_134),
.B2(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_2),
.B(n_195),
.C(n_199),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_2),
.B(n_120),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_2),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_2),
.B(n_98),
.Y(n_240)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_4),
.A2(n_169),
.B1(n_170),
.B2(n_174),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_4),
.Y(n_174)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_6),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_6),
.Y(n_229)
);

BUFx5_ASAP7_75t_L g239 ( 
.A(n_6),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_7),
.A2(n_100),
.B1(n_104),
.B2(n_108),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_7),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_7),
.A2(n_108),
.B1(n_205),
.B2(n_208),
.Y(n_204)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_9),
.A2(n_67),
.B1(n_94),
.B2(n_96),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_9),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_9),
.A2(n_96),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_9),
.A2(n_96),
.B1(n_234),
.B2(n_237),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_10),
.A2(n_21),
.B1(n_27),
.B2(n_28),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_11),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g166 ( 
.A(n_11),
.Y(n_166)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_12),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_12),
.Y(n_82)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_12),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_12),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_180),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_178),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_142),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_16),
.B(n_142),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_73),
.C(n_109),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_17),
.B(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_52),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_18),
.B(n_52),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_32),
.B(n_35),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_20),
.A2(n_36),
.B1(n_168),
.B2(n_175),
.Y(n_167)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx4_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_26),
.Y(n_210)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_31),
.Y(n_201)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_35),
.A2(n_233),
.B(n_239),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_44),
.Y(n_35)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_36),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_36),
.A2(n_213),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_39),
.Y(n_176)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_43),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_43),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_44),
.B(n_213),
.Y(n_212)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_47),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g227 ( 
.A(n_47),
.Y(n_227)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_50),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AOI32xp33_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_57),
.A3(n_59),
.B1(n_63),
.B2(n_66),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_55),
.A2(n_139),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_58),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

INVxp33_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp33_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_70),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_69),
.Y(n_151)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_69),
.Y(n_188)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_72),
.A2(n_114),
.B1(n_115),
.B2(n_118),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_73),
.A2(n_109),
.B1(n_110),
.B2(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_73),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_93),
.B1(n_97),
.B2(n_99),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_74),
.A2(n_99),
.B(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_74),
.A2(n_146),
.B(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_75),
.B(n_147),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_85),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_79),
.B1(n_81),
.B2(n_83),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_80),
.Y(n_198)
);

INVx4_ASAP7_75t_SL g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_85),
.A2(n_93),
.B(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_98),
.B(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

INVx5_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_130),
.B(n_136),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_120),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

AO22x2_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_124),
.B1(n_126),
.B2(n_128),
.Y(n_120)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_134),
.B(n_135),
.Y(n_130)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_162),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_134),
.A2(n_211),
.B(n_212),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_141),
.Y(n_136)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

INVx4_ASAP7_75t_SL g138 ( 
.A(n_139),
.Y(n_138)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_141),
.A2(n_155),
.B(n_158),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_153),
.B2(n_177),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_152),
.Y(n_144)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_160),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_167),
.Y(n_160)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI21x1_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_250),
.B(n_255),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_221),
.B(n_249),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_202),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_183),
.B(n_202),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_189),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_184),
.A2(n_189),
.B1(n_190),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_184),
.Y(n_247)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_215),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_203),
.B(n_216),
.C(n_220),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_211),
.B(n_212),
.Y(n_203)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_204),
.Y(n_245)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_242),
.B(n_248),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_231),
.B(n_241),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_230),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_228),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_240),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_240),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_233),
.Y(n_244)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_246),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_252),
.Y(n_255)
);


endmodule