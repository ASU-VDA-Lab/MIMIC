module fake_jpeg_27824_n_140 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_140);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx14_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NOR3xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_30),
.C(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_21),
.B1(n_19),
.B2(n_14),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_17),
.B1(n_25),
.B2(n_23),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_2),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_18),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_24),
.B1(n_21),
.B2(n_18),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_39),
.A2(n_16),
.B1(n_27),
.B2(n_20),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_48),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_21),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_47),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_35),
.A2(n_24),
.B1(n_36),
.B2(n_26),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_46),
.B1(n_25),
.B2(n_23),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_28),
.A2(n_26),
.B1(n_22),
.B2(n_17),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_49),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_55),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_48),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_SL g55 ( 
.A(n_45),
.B(n_18),
.C(n_32),
.Y(n_55)
);

OA21x2_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_63),
.B(n_38),
.Y(n_82)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_61),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_29),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_27),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_60),
.B(n_16),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_50),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_3),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_4),
.B(n_6),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_65),
.A2(n_44),
.B1(n_41),
.B2(n_7),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_20),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_12),
.Y(n_74)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_38),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_37),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_68),
.B(n_75),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_70),
.B(n_74),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_71),
.Y(n_96)
);

OAI32xp33_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_44),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_10),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_76),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_52),
.A2(n_38),
.B1(n_6),
.B2(n_7),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_59),
.B(n_10),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_83),
.B(n_64),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_54),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_83)
);

XNOR2x2_ASAP7_75t_SL g85 ( 
.A(n_73),
.B(n_55),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_75),
.B(n_54),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_87),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_73),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_93),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_71),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_81),
.A2(n_54),
.B(n_56),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_95),
.A2(n_97),
.B(n_81),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_68),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_98),
.B(n_100),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_99),
.B(n_101),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_87),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_81),
.C(n_82),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_107),
.C(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_105),
.A2(n_88),
.B1(n_85),
.B2(n_91),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_82),
.C(n_80),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_77),
.B1(n_79),
.B2(n_53),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_109),
.A2(n_96),
.B1(n_86),
.B2(n_79),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_115),
.C(n_118),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_102),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_95),
.C(n_93),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_109),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_70),
.C(n_83),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_120),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_107),
.C(n_99),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_122),
.B(n_123),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_104),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_123),
.A2(n_114),
.B1(n_110),
.B2(n_62),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_125),
.A2(n_67),
.B1(n_62),
.B2(n_51),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_121),
.B(n_89),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_127),
.B(n_128),
.Y(n_131)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_9),
.Y(n_135)
);

AOI211xp5_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_113),
.B(n_100),
.C(n_84),
.Y(n_132)
);

AOI322xp5_ASAP7_75t_L g134 ( 
.A1(n_132),
.A2(n_125),
.A3(n_98),
.B1(n_64),
.B2(n_9),
.C1(n_8),
.C2(n_57),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_133),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_133),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_135),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

AOI221xp5_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_136),
.B1(n_132),
.B2(n_138),
.C(n_131),
.Y(n_140)
);


endmodule