module fake_aes_971_n_42 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_42);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_42;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
NAND2xp5_ASAP7_75t_L g11 ( .A(n_9), .B(n_2), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_0), .Y(n_13) );
BUFx2_ASAP7_75t_L g14 ( .A(n_8), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_4), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_1), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_0), .Y(n_17) );
NOR3xp33_ASAP7_75t_SL g18 ( .A(n_15), .B(n_1), .C(n_2), .Y(n_18) );
BUFx6f_ASAP7_75t_L g19 ( .A(n_12), .Y(n_19) );
INVx6_ASAP7_75t_L g20 ( .A(n_14), .Y(n_20) );
BUFx2_ASAP7_75t_L g21 ( .A(n_15), .Y(n_21) );
NOR2xp33_ASAP7_75t_R g22 ( .A(n_14), .B(n_6), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_21), .Y(n_23) );
AOI22xp33_ASAP7_75t_L g24 ( .A1(n_20), .A2(n_17), .B1(n_16), .B2(n_13), .Y(n_24) );
AOI22xp33_ASAP7_75t_L g25 ( .A1(n_20), .A2(n_11), .B1(n_5), .B2(n_3), .Y(n_25) );
INVxp67_ASAP7_75t_L g26 ( .A(n_19), .Y(n_26) );
BUFx2_ASAP7_75t_SL g27 ( .A(n_23), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_26), .Y(n_28) );
HB1xp67_ASAP7_75t_L g29 ( .A(n_25), .Y(n_29) );
AND2x2_ASAP7_75t_L g30 ( .A(n_27), .B(n_24), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
NAND2x1p5_ASAP7_75t_L g32 ( .A(n_30), .B(n_27), .Y(n_32) );
NOR3xp33_ASAP7_75t_SL g33 ( .A(n_31), .B(n_18), .C(n_28), .Y(n_33) );
NAND2xp5_ASAP7_75t_L g34 ( .A(n_30), .B(n_29), .Y(n_34) );
NOR4xp25_ASAP7_75t_L g35 ( .A(n_34), .B(n_31), .C(n_18), .D(n_26), .Y(n_35) );
AND2x2_ASAP7_75t_L g36 ( .A(n_32), .B(n_22), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_33), .Y(n_37) );
HB1xp67_ASAP7_75t_L g38 ( .A(n_37), .Y(n_38) );
CKINVDCx5p33_ASAP7_75t_R g39 ( .A(n_37), .Y(n_39) );
AOI22xp33_ASAP7_75t_SL g40 ( .A1(n_38), .A2(n_36), .B1(n_19), .B2(n_35), .Y(n_40) );
AOI22xp5_ASAP7_75t_L g41 ( .A1(n_39), .A2(n_36), .B1(n_19), .B2(n_5), .Y(n_41) );
AOI222xp33_ASAP7_75t_L g42 ( .A1(n_40), .A2(n_3), .B1(n_7), .B2(n_10), .C1(n_38), .C2(n_41), .Y(n_42) );
endmodule