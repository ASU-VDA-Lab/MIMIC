module fake_jpeg_15125_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

INVx5_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVxp33_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_5),
.B(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_0),
.Y(n_18)
);

FAx1_ASAP7_75t_SL g33 ( 
.A(n_18),
.B(n_21),
.CI(n_1),
.CON(n_33),
.SN(n_33)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_12),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_22),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_17),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_6),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_15),
.B1(n_11),
.B2(n_10),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_16),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_27),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_13),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_32),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_23),
.B1(n_7),
.B2(n_14),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_14),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_41),
.B1(n_7),
.B2(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_40),
.Y(n_44)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_14),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_28),
.B(n_26),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_SL g49 ( 
.A(n_43),
.B(n_37),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_42),
.B1(n_38),
.B2(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_50),
.B(n_51),
.Y(n_53)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_38),
.B(n_49),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_55),
.C(n_33),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_44),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_33),
.B(n_45),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_19),
.C(n_29),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_19),
.Y(n_59)
);


endmodule