module fake_jpeg_568_n_226 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_226);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_25),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_28),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_10),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_6),
.B(n_33),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_3),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

BUFx10_ASAP7_75t_L g76 ( 
.A(n_3),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_84),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_65),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_59),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_65),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_80),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_83),
.Y(n_110)
);

BUFx12_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_92),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_67),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_93),
.B(n_59),
.Y(n_106)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_75),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_98),
.B(n_105),
.Y(n_124)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_84),
.B1(n_65),
.B2(n_67),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_102),
.A2(n_104),
.B1(n_66),
.B2(n_54),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_87),
.A2(n_54),
.B1(n_66),
.B2(n_73),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_87),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_106),
.B(n_107),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_93),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_90),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_58),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_85),
.B(n_71),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_109),
.B(n_112),
.Y(n_134)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_92),
.A2(n_91),
.B1(n_94),
.B2(n_95),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_78),
.B1(n_77),
.B2(n_96),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_86),
.Y(n_112)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_56),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_61),
.C(n_56),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_98),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_130),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_119),
.Y(n_151)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_126),
.A2(n_131),
.B1(n_135),
.B2(n_101),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_113),
.A2(n_97),
.B1(n_88),
.B2(n_64),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_128),
.A2(n_101),
.B1(n_68),
.B2(n_63),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_129),
.B(n_72),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_107),
.A2(n_62),
.B(n_61),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_88),
.B1(n_64),
.B2(n_55),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_100),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_138),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_55),
.B1(n_70),
.B2(n_68),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_69),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_140),
.B(n_152),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_99),
.C(n_103),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_150),
.C(n_128),
.Y(n_167)
);

AOI32xp33_ASAP7_75t_L g145 ( 
.A1(n_122),
.A2(n_60),
.A3(n_76),
.B1(n_66),
.B2(n_54),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_155),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_158),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_99),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_134),
.B(n_0),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_70),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_156),
.Y(n_168)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_127),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_157),
.A2(n_131),
.B1(n_127),
.B2(n_120),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_135),
.A2(n_76),
.B1(n_2),
.B2(n_4),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_118),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_160),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_1),
.Y(n_160)
);

AO21x1_ASAP7_75t_L g161 ( 
.A1(n_121),
.A2(n_76),
.B(n_26),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_161),
.A2(n_29),
.B(n_47),
.Y(n_175)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_169),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_172),
.B1(n_9),
.B2(n_11),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_148),
.Y(n_187)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_23),
.C(n_50),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_177),
.C(n_179),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_SL g171 ( 
.A1(n_143),
.A2(n_52),
.B(n_21),
.C(n_27),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_174),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_172)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_181),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_5),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_8),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_154),
.A2(n_161),
.B(n_144),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_7),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_178),
.B(n_180),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_20),
.C(n_43),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_141),
.B(n_7),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_155),
.A2(n_30),
.B(n_42),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_166),
.A2(n_148),
.B1(n_9),
.B2(n_10),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_183),
.A2(n_172),
.B1(n_179),
.B2(n_171),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_188),
.C(n_190),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_48),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_41),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_8),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_193),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_194),
.A2(n_171),
.B1(n_174),
.B2(n_13),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_173),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_196),
.B(n_197),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_195),
.A2(n_163),
.B(n_175),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_170),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_199),
.B(n_201),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_187),
.B(n_166),
.Y(n_200)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_200),
.Y(n_206)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_202),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_SL g204 ( 
.A1(n_186),
.A2(n_171),
.B(n_12),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_184),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_31),
.C(n_39),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_40),
.C(n_38),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_208),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_200),
.A2(n_189),
.B1(n_185),
.B2(n_15),
.Y(n_209)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_209),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_198),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_215),
.C(n_210),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_203),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_217),
.A2(n_218),
.B(n_206),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_216),
.B(n_207),
.Y(n_218)
);

OAI211xp5_ASAP7_75t_L g220 ( 
.A1(n_219),
.A2(n_211),
.B(n_214),
.C(n_212),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_36),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_221),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_222),
.A2(n_34),
.B(n_32),
.Y(n_223)
);

AOI311xp33_ASAP7_75t_L g224 ( 
.A1(n_223),
.A2(n_19),
.A3(n_13),
.B(n_15),
.C(n_16),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_224),
.A2(n_11),
.B1(n_17),
.B2(n_18),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_17),
.Y(n_226)
);


endmodule