module fake_jpeg_7042_n_256 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_256);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_25),
.Y(n_26)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_12),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_27),
.B(n_34),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx5_ASAP7_75t_SL g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_13),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_27),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_20),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_16),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_26),
.A2(n_20),
.B1(n_23),
.B2(n_16),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_20),
.B1(n_13),
.B2(n_17),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_26),
.A2(n_20),
.B1(n_13),
.B2(n_17),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_13),
.B1(n_17),
.B2(n_16),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_32),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_59),
.B1(n_36),
.B2(n_43),
.Y(n_72)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_51),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_52),
.A2(n_58),
.B(n_36),
.Y(n_67)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_53),
.B(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_32),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_32),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_36),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_57),
.A2(n_60),
.B1(n_38),
.B2(n_37),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_20),
.B1(n_33),
.B2(n_30),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_30),
.B1(n_33),
.B2(n_31),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_35),
.A2(n_33),
.B1(n_38),
.B2(n_40),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_42),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_61),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_78),
.B1(n_60),
.B2(n_59),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_56),
.Y(n_80)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_73),
.Y(n_83)
);

BUFx4f_ASAP7_75t_SL g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_74),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_53),
.B1(n_54),
.B2(n_59),
.Y(n_84)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

AO22x1_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_37),
.B1(n_40),
.B2(n_43),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_50),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_84),
.B1(n_86),
.B2(n_90),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_65),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_85),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_63),
.B(n_64),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_76),
.B(n_55),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_92),
.Y(n_102)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_68),
.Y(n_105)
);

NAND3xp33_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_61),
.C(n_52),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_54),
.B1(n_56),
.B2(n_55),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_78),
.A2(n_52),
.B1(n_58),
.B2(n_48),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_91),
.A2(n_94),
.B1(n_62),
.B2(n_38),
.Y(n_104)
);

MAJx2_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_58),
.C(n_52),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_69),
.A2(n_48),
.B1(n_47),
.B2(n_38),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_96),
.Y(n_110)
);

MAJx2_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_41),
.C(n_28),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_48),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

AO21x1_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_78),
.B(n_73),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_86),
.B(n_80),
.Y(n_117)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_108),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_101),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_106),
.B1(n_112),
.B2(n_35),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_105),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_70),
.B1(n_71),
.B2(n_74),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_93),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_77),
.B1(n_75),
.B2(n_67),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_23),
.B1(n_14),
.B2(n_29),
.Y(n_131)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_115),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_91),
.A2(n_63),
.B1(n_35),
.B2(n_41),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_39),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_90),
.Y(n_118)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_65),
.Y(n_116)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_117),
.A2(n_106),
.B(n_98),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_0),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_95),
.Y(n_119)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_80),
.Y(n_120)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_34),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_107),
.A2(n_96),
.B1(n_92),
.B2(n_35),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_127),
.B1(n_131),
.B2(n_34),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_102),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_130),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_100),
.B1(n_108),
.B2(n_115),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_107),
.A2(n_92),
.B1(n_70),
.B2(n_33),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_70),
.B1(n_23),
.B2(n_14),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_128),
.A2(n_103),
.B1(n_99),
.B2(n_22),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_17),
.Y(n_129)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_28),
.C(n_31),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_112),
.C(n_106),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_135),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_105),
.A2(n_23),
.B(n_25),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_123),
.B(n_100),
.Y(n_137)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_106),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_139),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_116),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_153),
.Y(n_166)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_113),
.B1(n_98),
.B2(n_103),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_142),
.A2(n_150),
.B1(n_128),
.B2(n_134),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_148),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_123),
.B(n_11),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_151),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_28),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_0),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_129),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_127),
.B(n_28),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_157),
.C(n_136),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_132),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_156),
.Y(n_163)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

XNOR2x1_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_133),
.Y(n_158)
);

MAJx2_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_176),
.C(n_28),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_130),
.C(n_133),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_159),
.B(n_161),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_119),
.C(n_120),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_134),
.C(n_118),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_169),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_164),
.A2(n_22),
.B1(n_19),
.B2(n_18),
.Y(n_192)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_131),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_155),
.C(n_146),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_171),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_135),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_124),
.C(n_121),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_173),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_139),
.A2(n_121),
.B1(n_22),
.B2(n_19),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_153),
.B(n_28),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_154),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_178),
.A2(n_186),
.B(n_188),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_160),
.B(n_152),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_179),
.B(n_195),
.Y(n_197)
);

AOI322xp5_ASAP7_75t_L g181 ( 
.A1(n_177),
.A2(n_147),
.A3(n_148),
.B1(n_34),
.B2(n_31),
.C1(n_29),
.C2(n_22),
.Y(n_181)
);

BUFx24_ASAP7_75t_SL g204 ( 
.A(n_181),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_163),
.Y(n_182)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

BUFx24_ASAP7_75t_SL g183 ( 
.A(n_166),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_183),
.B(n_21),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_12),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_11),
.Y(n_189)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_192),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_170),
.A2(n_34),
.B1(n_31),
.B2(n_29),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_194),
.A2(n_29),
.B1(n_22),
.B2(n_19),
.Y(n_202)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_161),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_196),
.B(n_0),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_159),
.C(n_174),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_203),
.C(n_185),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_190),
.A2(n_176),
.B(n_1),
.Y(n_200)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_200),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_11),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_206),
.B(n_1),
.Y(n_222)
);

NAND2xp33_ASAP7_75t_SL g207 ( 
.A(n_186),
.B(n_0),
.Y(n_207)
);

FAx1_ASAP7_75t_SL g225 ( 
.A(n_207),
.B(n_200),
.CI(n_202),
.CON(n_225),
.SN(n_225)
);

OAI322xp33_ASAP7_75t_L g208 ( 
.A1(n_191),
.A2(n_21),
.A3(n_15),
.B1(n_19),
.B2(n_18),
.C1(n_4),
.C2(n_5),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_208),
.A2(n_21),
.B1(n_15),
.B2(n_3),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_1),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_211),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_185),
.C(n_187),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_191),
.C(n_193),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_216),
.B(n_225),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_212),
.A2(n_184),
.B1(n_192),
.B2(n_3),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_220),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_198),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_197),
.A2(n_19),
.B1(n_18),
.B2(n_4),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_5),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_223),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_210),
.B(n_2),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_2),
.Y(n_231)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_203),
.C(n_201),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_213),
.C(n_215),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_232),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_204),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_233),
.B(n_234),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_18),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_218),
.A2(n_18),
.B1(n_6),
.B2(n_7),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_235),
.Y(n_241)
);

AOI31xp67_ASAP7_75t_SL g236 ( 
.A1(n_225),
.A2(n_5),
.A3(n_7),
.B(n_8),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_236),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_217),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_238),
.A2(n_240),
.B(n_228),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_229),
.B(n_218),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_243),
.B(n_242),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_250),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_249),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_238),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_246),
.A2(n_247),
.B(n_248),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_241),
.A2(n_227),
.B(n_9),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_239),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_8),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_10),
.C(n_15),
.Y(n_250)
);

AOI321xp33_ASAP7_75t_L g254 ( 
.A1(n_253),
.A2(n_10),
.A3(n_15),
.B1(n_21),
.B2(n_252),
.C(n_251),
.Y(n_254)
);

AO21x1_ASAP7_75t_L g255 ( 
.A1(n_254),
.A2(n_15),
.B(n_21),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_21),
.Y(n_256)
);


endmodule