module fake_jpeg_29030_n_546 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_546);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_546;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_434;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_3),
.B(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_56),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_8),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_58),
.B(n_74),
.Y(n_115)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_8),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_62),
.B(n_73),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_65),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_66),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_69),
.Y(n_138)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_70),
.Y(n_146)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_71),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_8),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_85),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_22),
.B(n_9),
.Y(n_73)
);

NOR3xp33_ASAP7_75t_L g74 ( 
.A(n_22),
.B(n_9),
.C(n_14),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_76),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_77),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_78),
.Y(n_177)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_81),
.Y(n_178)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_82),
.Y(n_140)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_83),
.Y(n_155)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_19),
.B(n_9),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_86),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_19),
.B(n_9),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_87),
.B(n_106),
.Y(n_172)
);

OR2x2_ASAP7_75t_SL g88 ( 
.A(n_43),
.B(n_7),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_89),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_39),
.B(n_12),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_91),
.Y(n_167)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_92),
.Y(n_175)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_96),
.Y(n_147)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_98),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_18),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_101),
.Y(n_158)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_104),
.Y(n_174)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_105),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_25),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_29),
.B(n_12),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_46),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_41),
.Y(n_108)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_44),
.Y(n_109)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_44),
.Y(n_110)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_110),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_104),
.A2(n_53),
.B1(n_36),
.B2(n_44),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_111),
.A2(n_143),
.B1(n_152),
.B2(n_53),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_72),
.A2(n_34),
.B1(n_52),
.B2(n_29),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_116),
.A2(n_134),
.B1(n_37),
.B2(n_17),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_73),
.A2(n_25),
.B1(n_43),
.B2(n_35),
.Y(n_122)
);

AO22x1_ASAP7_75t_L g215 ( 
.A1(n_122),
.A2(n_1),
.B1(n_2),
.B2(n_6),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_130),
.B(n_151),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_105),
.A2(n_44),
.B1(n_54),
.B2(n_47),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_55),
.Y(n_135)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_135),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_92),
.A2(n_53),
.B1(n_36),
.B2(n_54),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_58),
.B(n_25),
.C(n_40),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_150),
.B(n_37),
.C(n_17),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_87),
.B(n_34),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_74),
.A2(n_53),
.B1(n_54),
.B2(n_35),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_106),
.B(n_50),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_154),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_56),
.B(n_50),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_89),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_157),
.B(n_173),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_59),
.A2(n_38),
.B1(n_52),
.B2(n_46),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_39),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_71),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_63),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_65),
.A2(n_54),
.B1(n_53),
.B2(n_35),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_171),
.A2(n_2),
.B1(n_165),
.B2(n_170),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_66),
.B(n_38),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_179),
.B(n_181),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_183),
.A2(n_210),
.B1(n_213),
.B2(n_142),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_157),
.A2(n_108),
.B1(n_98),
.B2(n_95),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_185),
.A2(n_192),
.B1(n_201),
.B2(n_215),
.Y(n_235)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_186),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_31),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_187),
.B(n_194),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_121),
.A2(n_31),
.B1(n_51),
.B2(n_45),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_188),
.A2(n_189),
.B1(n_191),
.B2(n_195),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_123),
.A2(n_28),
.B1(n_51),
.B2(n_45),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_126),
.A2(n_40),
.B1(n_28),
.B2(n_132),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_124),
.A2(n_90),
.B1(n_81),
.B2(n_78),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_149),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_193),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_128),
.B(n_119),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_164),
.A2(n_77),
.B1(n_25),
.B2(n_47),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_196),
.B(n_203),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_173),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_197),
.B(n_200),
.Y(n_236)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_129),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_198),
.Y(n_240)
);

O2A1O1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_122),
.A2(n_49),
.B(n_32),
.C(n_16),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_199),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_117),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_178),
.A2(n_134),
.B1(n_122),
.B2(n_136),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_115),
.B(n_49),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_127),
.Y(n_204)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_204),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_120),
.A2(n_32),
.B1(n_16),
.B2(n_5),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_205),
.A2(n_221),
.B1(n_135),
.B2(n_131),
.Y(n_245)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_118),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_207),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_129),
.Y(n_208)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_208),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_167),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_209),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_152),
.A2(n_111),
.B1(n_143),
.B2(n_112),
.Y(n_210)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_211),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_114),
.B(n_16),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_212),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_156),
.A2(n_12),
.B1(n_14),
.B2(n_5),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_117),
.B(n_5),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_224),
.Y(n_238)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_147),
.Y(n_216)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_158),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_217),
.Y(n_265)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_174),
.Y(n_218)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_218),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_120),
.A2(n_6),
.B1(n_13),
.B2(n_15),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_219),
.A2(n_230),
.B1(n_177),
.B2(n_137),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_168),
.B(n_146),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_220),
.B(n_225),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_136),
.A2(n_2),
.B1(n_6),
.B2(n_165),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_118),
.Y(n_222)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_139),
.Y(n_223)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_223),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_170),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_133),
.B(n_138),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_166),
.Y(n_226)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_226),
.Y(n_257)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_140),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_228),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_113),
.B(n_6),
.Y(n_228)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_163),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_231),
.Y(n_250)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_163),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_141),
.B(n_176),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_233),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_125),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_207),
.Y(n_242)
);

INVx11_ASAP7_75t_L g277 ( 
.A(n_242),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_244),
.A2(n_212),
.B1(n_214),
.B2(n_194),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_245),
.A2(n_190),
.B1(n_211),
.B2(n_231),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_246),
.B(n_271),
.Y(n_283)
);

INVx13_ASAP7_75t_L g249 ( 
.A(n_182),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_249),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_253),
.A2(n_258),
.B1(n_262),
.B2(n_273),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_184),
.B(n_125),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_255),
.B(n_269),
.Y(n_290)
);

CKINVDCx12_ASAP7_75t_R g256 ( 
.A(n_233),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_256),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_215),
.A2(n_177),
.B1(n_137),
.B2(n_145),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_215),
.A2(n_145),
.B1(n_161),
.B2(n_169),
.Y(n_262)
);

INVx13_ASAP7_75t_L g267 ( 
.A(n_182),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_267),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_184),
.B(n_197),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_180),
.B(n_171),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_210),
.A2(n_169),
.B1(n_161),
.B2(n_155),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_266),
.A2(n_181),
.B(n_199),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_275),
.A2(n_279),
.B(n_264),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_266),
.A2(n_179),
.B1(n_181),
.B2(n_206),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_276),
.A2(n_302),
.B1(n_279),
.B2(n_281),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_265),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_278),
.B(n_288),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_244),
.A2(n_212),
.B(n_206),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_271),
.A2(n_230),
.B1(n_225),
.B2(n_208),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_280),
.A2(n_284),
.B1(n_295),
.B2(n_235),
.Y(n_316)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_265),
.Y(n_282)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_282),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_272),
.A2(n_208),
.B1(n_204),
.B2(n_198),
.Y(n_284)
);

BUFx24_ASAP7_75t_SL g285 ( 
.A(n_269),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_285),
.Y(n_312)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_239),
.Y(n_286)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_286),
.Y(n_311)
);

AND2x4_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_232),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_287),
.B(n_247),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_265),
.Y(n_288)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_239),
.Y(n_291)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_291),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_237),
.A2(n_203),
.B(n_228),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_292),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_236),
.B(n_180),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_294),
.B(n_297),
.Y(n_314)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_259),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_296),
.Y(n_331)
);

AO22x1_ASAP7_75t_SL g297 ( 
.A1(n_237),
.A2(n_223),
.B1(n_227),
.B2(n_186),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_237),
.A2(n_216),
.B1(n_217),
.B2(n_224),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_298),
.A2(n_303),
.B1(n_274),
.B2(n_242),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_236),
.B(n_196),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_299),
.B(n_247),
.Y(n_322)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_241),
.Y(n_300)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_300),
.Y(n_325)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_259),
.Y(n_301)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_301),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_237),
.A2(n_213),
.B1(n_198),
.B2(n_222),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_256),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_305),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_255),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_264),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_234),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_308),
.B(n_287),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_309),
.A2(n_316),
.B1(n_321),
.B2(n_326),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_283),
.A2(n_238),
.B(n_243),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_313),
.A2(n_328),
.B(n_333),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_290),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_315),
.B(n_322),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_247),
.C(n_251),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_318),
.B(n_287),
.C(n_304),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_302),
.A2(n_251),
.B1(n_238),
.B2(n_243),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_324),
.B(n_332),
.Y(n_354)
);

OAI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_275),
.A2(n_270),
.B1(n_241),
.B2(n_240),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_327),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_275),
.B(n_250),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_286),
.Y(n_330)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_330),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_307),
.B(n_234),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_283),
.A2(n_247),
.B(n_248),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_305),
.B(n_248),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_334),
.B(n_335),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_290),
.B(n_250),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_336),
.A2(n_295),
.B1(n_298),
.B2(n_280),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_293),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_337),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_338),
.B(n_350),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_322),
.B(n_292),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_339),
.B(n_313),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_334),
.B(n_287),
.Y(n_343)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_343),
.Y(n_371)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_323),
.Y(n_344)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_344),
.Y(n_393)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_311),
.Y(n_348)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_348),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_328),
.A2(n_276),
.B(n_303),
.Y(n_349)
);

AO21x1_ASAP7_75t_L g369 ( 
.A1(n_349),
.A2(n_357),
.B(n_359),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_336),
.A2(n_295),
.B1(n_298),
.B2(n_294),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_352),
.B(n_353),
.C(n_327),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_318),
.B(n_287),
.C(n_289),
.Y(n_353)
);

FAx1_ASAP7_75t_L g396 ( 
.A(n_355),
.B(n_300),
.CI(n_281),
.CON(n_396),
.SN(n_396)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_311),
.Y(n_356)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_356),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_328),
.A2(n_284),
.B(n_287),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_320),
.Y(n_358)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_358),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_328),
.A2(n_309),
.B(n_314),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_320),
.Y(n_360)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_360),
.Y(n_375)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_325),
.Y(n_361)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_361),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_314),
.A2(n_306),
.B(n_297),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_362),
.A2(n_327),
.B(n_326),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_315),
.B(n_297),
.Y(n_363)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_363),
.Y(n_387)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_325),
.Y(n_364)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_364),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_321),
.B(n_257),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_365),
.B(n_362),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_323),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_366),
.B(n_337),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_354),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_370),
.B(n_384),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_373),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_374),
.B(n_381),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_353),
.B(n_318),
.C(n_327),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_376),
.B(n_386),
.C(n_389),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_340),
.B(n_354),
.Y(n_377)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_377),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_340),
.B(n_335),
.Y(n_378)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_378),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_352),
.B(n_308),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_379),
.B(n_380),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_339),
.B(n_333),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_342),
.A2(n_310),
.B1(n_316),
.B2(n_324),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_383),
.A2(n_338),
.B1(n_342),
.B2(n_361),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_346),
.A2(n_319),
.B(n_317),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_385),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_355),
.B(n_310),
.C(n_319),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_345),
.B(n_317),
.C(n_332),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_390),
.B(n_347),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_341),
.B(n_330),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_391),
.B(n_396),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_363),
.B(n_297),
.Y(n_392)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_392),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_351),
.B(n_291),
.Y(n_394)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_394),
.Y(n_407)
);

BUFx12f_ASAP7_75t_L g397 ( 
.A(n_393),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_397),
.B(n_402),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_377),
.B(n_351),
.Y(n_401)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_401),
.Y(n_446)
);

BUFx12_ASAP7_75t_L g402 ( 
.A(n_384),
.Y(n_402)
);

MAJx2_ASAP7_75t_L g403 ( 
.A(n_374),
.B(n_359),
.C(n_343),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_403),
.B(n_426),
.Y(n_438)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_394),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_408),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_389),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_409),
.B(n_416),
.Y(n_433)
);

NOR3xp33_ASAP7_75t_L g410 ( 
.A(n_386),
.B(n_349),
.C(n_346),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_410),
.B(n_422),
.Y(n_436)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_375),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_411),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_376),
.B(n_357),
.C(n_350),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_413),
.B(n_380),
.C(n_368),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_378),
.B(n_312),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_417),
.A2(n_368),
.B1(n_387),
.B2(n_392),
.Y(n_431)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_375),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_418),
.B(n_420),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_419),
.B(n_421),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_393),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_382),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_391),
.B(n_257),
.Y(n_422)
);

OR2x4_ASAP7_75t_L g423 ( 
.A(n_371),
.B(n_387),
.Y(n_423)
);

AO21x1_ASAP7_75t_L g442 ( 
.A1(n_423),
.A2(n_369),
.B(n_388),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_381),
.B(n_356),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_424),
.A2(n_404),
.B1(n_423),
.B2(n_414),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_379),
.B(n_358),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_428),
.B(n_445),
.Y(n_465)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_401),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_429),
.B(n_444),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_400),
.B(n_398),
.C(n_413),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_430),
.B(n_434),
.C(n_439),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_431),
.A2(n_425),
.B1(n_402),
.B2(n_412),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_400),
.B(n_373),
.C(n_371),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_398),
.B(n_383),
.C(n_396),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_426),
.B(n_396),
.C(n_382),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_441),
.B(n_450),
.C(n_331),
.Y(n_460)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_442),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_414),
.A2(n_399),
.B1(n_407),
.B2(n_405),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_443),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_403),
.B(n_369),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_417),
.A2(n_388),
.B1(n_395),
.B2(n_372),
.Y(n_447)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_447),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_415),
.A2(n_367),
.B1(n_360),
.B2(n_364),
.Y(n_448)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_448),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_425),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_449),
.B(n_288),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_412),
.B(n_347),
.C(n_348),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_433),
.A2(n_415),
.B1(n_406),
.B2(n_420),
.Y(n_452)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_452),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_457),
.A2(n_443),
.B1(n_444),
.B2(n_438),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g458 ( 
.A1(n_440),
.A2(n_397),
.B1(n_366),
.B2(n_344),
.Y(n_458)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_458),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_427),
.B(n_402),
.Y(n_459)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_459),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_460),
.B(n_463),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_446),
.A2(n_397),
.B(n_366),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_461),
.A2(n_261),
.B(n_252),
.Y(n_488)
);

INVx1_ASAP7_75t_SL g462 ( 
.A(n_446),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_462),
.B(n_466),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_430),
.B(n_329),
.C(n_278),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_464),
.B(n_470),
.C(n_434),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_435),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_440),
.A2(n_331),
.B1(n_329),
.B2(n_323),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_468),
.B(n_469),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_428),
.B(n_254),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_450),
.B(n_282),
.C(n_296),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_437),
.B(n_301),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_471),
.A2(n_293),
.B1(n_254),
.B2(n_268),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_472),
.B(n_464),
.Y(n_490)
);

MAJx2_ASAP7_75t_L g473 ( 
.A(n_454),
.B(n_439),
.C(n_441),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_473),
.B(n_475),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_456),
.A2(n_431),
.B1(n_436),
.B2(n_442),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_476),
.A2(n_486),
.B1(n_455),
.B2(n_468),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_459),
.A2(n_436),
.B(n_438),
.Y(n_477)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_477),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_451),
.A2(n_432),
.B1(n_242),
.B2(n_277),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_480),
.B(n_487),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_465),
.B(n_261),
.C(n_270),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_482),
.B(n_485),
.C(n_470),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_465),
.B(n_261),
.C(n_270),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_453),
.A2(n_240),
.B1(n_293),
.B2(n_260),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_488),
.B(n_457),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_454),
.A2(n_268),
.B(n_252),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_489),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_490),
.B(n_494),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_484),
.B(n_461),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_495),
.B(n_496),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_481),
.B(n_459),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_498),
.B(n_499),
.Y(n_514)
);

CKINVDCx14_ASAP7_75t_R g499 ( 
.A(n_478),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_480),
.B(n_462),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_500),
.B(n_502),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_472),
.B(n_469),
.C(n_460),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_501),
.B(n_240),
.C(n_190),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_481),
.B(n_467),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_503),
.B(n_505),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_474),
.A2(n_455),
.B(n_268),
.Y(n_504)
);

AOI21x1_ASAP7_75t_L g506 ( 
.A1(n_504),
.A2(n_488),
.B(n_479),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_476),
.B(n_277),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_506),
.B(n_495),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_493),
.A2(n_475),
.B1(n_483),
.B2(n_473),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_507),
.B(n_518),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_501),
.A2(n_494),
.B(n_491),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_510),
.B(n_511),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_492),
.A2(n_486),
.B1(n_485),
.B2(n_482),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_500),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_512),
.B(n_517),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_504),
.A2(n_483),
.B(n_277),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_515),
.B(n_263),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_490),
.B(n_260),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_497),
.B(n_260),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_519),
.B(n_263),
.C(n_202),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_519),
.B(n_497),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_521),
.B(n_522),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_R g525 ( 
.A1(n_512),
.A2(n_502),
.B(n_498),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_525),
.A2(n_529),
.B1(n_513),
.B2(n_515),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_514),
.B(n_202),
.C(n_263),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_526),
.B(n_527),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_508),
.B(n_218),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_SL g532 ( 
.A(n_528),
.B(n_509),
.Y(n_532)
);

INVxp67_ASAP7_75t_SL g531 ( 
.A(n_523),
.Y(n_531)
);

OAI21x1_ASAP7_75t_L g536 ( 
.A1(n_531),
.A2(n_532),
.B(n_534),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_533),
.B(n_522),
.C(n_524),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g534 ( 
.A(n_520),
.B(n_516),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_537),
.B(n_538),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_535),
.A2(n_527),
.B(n_529),
.Y(n_538)
);

AOI21xp33_ASAP7_75t_L g539 ( 
.A1(n_530),
.A2(n_267),
.B(n_249),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_539),
.B(n_209),
.C(n_193),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_540),
.B(n_222),
.C(n_536),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g543 ( 
.A1(n_542),
.A2(n_541),
.B(n_229),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_543),
.A2(n_148),
.B(n_249),
.Y(n_544)
);

BUFx24_ASAP7_75t_SL g545 ( 
.A(n_544),
.Y(n_545)
);

FAx1_ASAP7_75t_SL g546 ( 
.A(n_545),
.B(n_267),
.CI(n_2),
.CON(n_546),
.SN(n_546)
);


endmodule