module real_jpeg_26713_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_139;
wire n_33;
wire n_188;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_244;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_0),
.A2(n_39),
.B1(n_76),
.B2(n_77),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_0),
.A2(n_39),
.B1(n_57),
.B2(n_59),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_0),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_1),
.B(n_27),
.Y(n_26)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_1),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_2),
.A2(n_43),
.B1(n_44),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_2),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_52),
.Y(n_98)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_4),
.A2(n_76),
.B1(n_77),
.B2(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_4),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_4),
.A2(n_57),
.B1(n_59),
.B2(n_138),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_4),
.A2(n_43),
.B1(n_44),
.B2(n_138),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_138),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_6),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_6),
.B(n_79),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_6),
.B(n_59),
.Y(n_181)
);

AOI21xp33_ASAP7_75t_L g185 ( 
.A1(n_6),
.A2(n_59),
.B(n_181),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_6),
.A2(n_43),
.B1(n_44),
.B2(n_126),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_6),
.A2(n_11),
.B(n_28),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_6),
.B(n_60),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_6),
.A2(n_35),
.B1(n_88),
.B2(n_230),
.Y(n_232)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_8),
.A2(n_43),
.B1(n_44),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_8),
.A2(n_50),
.B1(n_57),
.B2(n_59),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_50),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_9),
.A2(n_76),
.B1(n_77),
.B2(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_9),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_9),
.A2(n_57),
.B1(n_59),
.B2(n_81),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_9),
.A2(n_43),
.B1(n_44),
.B2(n_81),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_81),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_10),
.A2(n_76),
.B1(n_77),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_10),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_10),
.A2(n_57),
.B1(n_59),
.B2(n_112),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_10),
.A2(n_43),
.B1(n_44),
.B2(n_112),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_112),
.Y(n_222)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_12),
.A2(n_32),
.B1(n_57),
.B2(n_59),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_12),
.A2(n_32),
.B1(n_43),
.B2(n_44),
.Y(n_92)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_15),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_141),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_139),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_114),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_19),
.B(n_114),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_95),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_84),
.B2(n_85),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_53),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_40),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_24),
.B(n_40),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_33),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_25),
.A2(n_128),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_26),
.A2(n_38),
.B(n_100),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_26),
.A2(n_34),
.B1(n_221),
.B2(n_223),
.Y(n_220)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_27),
.A2(n_28),
.B1(n_46),
.B2(n_47),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_27),
.B(n_234),
.Y(n_233)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_31),
.B(n_37),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_33),
.A2(n_88),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_38),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_35),
.A2(n_88),
.B(n_89),
.Y(n_87)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_SL g129 ( 
.A(n_36),
.Y(n_129)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_37),
.A2(n_88),
.B1(n_222),
.B2(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_37),
.B(n_126),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_41),
.A2(n_51),
.B(n_91),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_41),
.A2(n_91),
.B(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_41),
.A2(n_48),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_41),
.A2(n_189),
.B(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_41),
.A2(n_48),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_41),
.A2(n_48),
.B1(n_188),
.B2(n_207),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_48),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_44),
.B1(n_62),
.B2(n_64),
.Y(n_61)
);

AOI32xp33_ASAP7_75t_L g179 ( 
.A1(n_43),
.A2(n_57),
.A3(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_179)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp33_ASAP7_75t_SL g182 ( 
.A(n_44),
.B(n_69),
.Y(n_182)
);

A2O1A1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_44),
.A2(n_47),
.B(n_126),
.C(n_209),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_48),
.A2(n_49),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_48),
.B(n_126),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_70),
.B2(n_71),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_60),
.B(n_65),
.Y(n_55)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_59),
.B1(n_63),
.B2(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_59),
.B1(n_74),
.B2(n_75),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_57),
.A2(n_78),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_59),
.B(n_74),
.Y(n_124)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_61),
.B(n_66),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_61),
.B(n_107),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_61),
.A2(n_67),
.B1(n_132),
.B2(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_61),
.A2(n_67),
.B1(n_153),
.B2(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_61),
.A2(n_67),
.B1(n_166),
.B2(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_69),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_80),
.B(n_82),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_72),
.A2(n_80),
.B1(n_111),
.B2(n_113),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_72),
.A2(n_111),
.B1(n_113),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_73),
.A2(n_79),
.B1(n_125),
.B2(n_137),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_76),
.B(n_78),
.C(n_79),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_76),
.Y(n_78)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

HAxp5_ASAP7_75t_SL g125 ( 
.A(n_76),
.B(n_126),
.CON(n_125),
.SN(n_125)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_79),
.B(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_90),
.B2(n_94),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_88),
.A2(n_98),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_90),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_92),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_93),
.B(n_150),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_104),
.C(n_109),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_101),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_97),
.B(n_101),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_104),
.A2(n_109),
.B1(n_110),
.B2(n_117),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_104),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B(n_108),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_131),
.B(n_133),
.Y(n_130)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.C(n_120),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_115),
.A2(n_118),
.B1(n_119),
.B2(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_115),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_120),
.A2(n_121),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_130),
.C(n_134),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_122),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_123),
.B(n_127),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_130),
.A2(n_134),
.B1(n_135),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_130),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_171),
.B(n_253),
.C(n_259),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_158),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_143),
.B(n_158),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_155),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_145),
.B(n_146),
.C(n_155),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.C(n_154),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_147),
.A2(n_148),
.B1(n_151),
.B2(n_152),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_154),
.B(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.C(n_164),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_159),
.A2(n_160),
.B1(n_248),
.B2(n_250),
.Y(n_247)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_164),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.C(n_169),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_169),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_252),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_245),
.B(n_251),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_200),
.B(n_244),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_190),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_175),
.B(n_190),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_183),
.C(n_186),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_176),
.A2(n_177),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_179),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_183),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_195),
.B2(n_196),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_191),
.B(n_197),
.C(n_198),
.Y(n_246)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_238),
.B(n_243),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_218),
.B(n_237),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_210),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_203),
.B(n_210),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_208),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_204),
.A2(n_205),
.B1(n_208),
.B2(n_225),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_208),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_216),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_215),
.C(n_216),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_217),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_226),
.B(n_236),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_224),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_220),
.B(n_224),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_231),
.B(n_235),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_228),
.B(n_229),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_239),
.B(n_240),
.Y(n_243)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_246),
.B(n_247),
.Y(n_251)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_248),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_254),
.B(n_255),
.Y(n_259)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);


endmodule