module fake_jpeg_2692_n_69 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_69);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_69;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_32;
wire n_66;

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_21),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_5),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_20),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_30),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_19),
.B1(n_18),
.B2(n_16),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_26),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_24),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_33),
.B(n_25),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_34),
.B(n_38),
.Y(n_43)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_26),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_27),
.B1(n_23),
.B2(n_22),
.Y(n_44)
);

NOR2x1_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_27),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_29),
.C(n_23),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_25),
.C(n_24),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_22),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_48),
.B(n_49),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_47),
.A2(n_40),
.B(n_37),
.Y(n_49)
);

AND2x6_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_13),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_50),
.B(n_11),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_52),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_54),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_1),
.B(n_2),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_58),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_51),
.A2(n_42),
.B1(n_43),
.B2(n_41),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_52),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_55),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_61),
.A2(n_56),
.B1(n_59),
.B2(n_6),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_9),
.C(n_4),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_55),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_65),
.C(n_62),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_64),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_3),
.C(n_5),
.Y(n_68)
);

AOI311xp33_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_6),
.A3(n_7),
.B(n_8),
.C(n_50),
.Y(n_69)
);


endmodule