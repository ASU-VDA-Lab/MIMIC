module real_jpeg_24768_n_23 (n_17, n_108, n_8, n_116, n_0, n_21, n_111, n_2, n_10, n_114, n_9, n_12, n_6, n_11, n_14, n_110, n_112, n_7, n_22, n_18, n_3, n_117, n_5, n_4, n_109, n_115, n_1, n_20, n_19, n_16, n_15, n_13, n_113, n_23);

input n_17;
input n_108;
input n_8;
input n_116;
input n_0;
input n_21;
input n_111;
input n_2;
input n_10;
input n_114;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_110;
input n_112;
input n_7;
input n_22;
input n_18;
input n_3;
input n_117;
input n_5;
input n_4;
input n_109;
input n_115;
input n_1;
input n_20;
input n_19;
input n_16;
input n_15;
input n_13;
input n_113;

output n_23;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_87;
wire n_105;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_30;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_1),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_3),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_4),
.B(n_36),
.C(n_89),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_5),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_6),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_7),
.B(n_42),
.C(n_63),
.Y(n_41)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_8),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_9),
.B(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_11),
.B(n_34),
.C(n_99),
.Y(n_33)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_12),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_13),
.B(n_44),
.C(n_55),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_38),
.C(n_78),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_15),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_16),
.Y(n_101)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_32),
.C(n_105),
.Y(n_31)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_20),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_40),
.C(n_71),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_22),
.A2(n_25),
.B1(n_26),
.B2(n_30),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_31),
.Y(n_23)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_28),
.B(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_28),
.B(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_28),
.B(n_106),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_29),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_29),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_101),
.C(n_102),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_92),
.C(n_93),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_82),
.C(n_83),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_74),
.C(n_75),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_65),
.C(n_66),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_58),
.C(n_59),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_50),
.C(n_51),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_49),
.Y(n_62)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_108),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_109),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_110),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_111),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_112),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_113),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_114),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_115),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_116),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_117),
.Y(n_85)
);


endmodule