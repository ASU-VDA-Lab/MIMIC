module fake_jpeg_2556_n_47 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_43;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_SL g7 ( 
.A(n_6),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_4),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_6),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_16),
.B(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_1),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_11),
.B(n_2),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_16),
.Y(n_30)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_13),
.A2(n_5),
.B1(n_2),
.B2(n_3),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_11),
.A2(n_2),
.B1(n_5),
.B2(n_13),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_23),
.B(n_14),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_26),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_L g27 ( 
.A1(n_23),
.A2(n_10),
.B1(n_15),
.B2(n_12),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_30),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_21),
.A2(n_5),
.B1(n_12),
.B2(n_17),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_23),
.B(n_22),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g32 ( 
.A(n_25),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_32),
.A2(n_34),
.B1(n_21),
.B2(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_30),
.C(n_19),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_35),
.A2(n_24),
.B1(n_28),
.B2(n_26),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_38),
.C(n_39),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_31),
.C(n_36),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_31),
.C(n_37),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_43),
.C(n_35),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_34),
.B(n_29),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_29),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_45),
.A2(n_20),
.B(n_32),
.Y(n_46)
);

BUFx24_ASAP7_75t_SL g47 ( 
.A(n_46),
.Y(n_47)
);


endmodule