module fake_jpeg_884_n_618 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_618);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_618;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_387;
wire n_270;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_15),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_8),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_20),
.B(n_17),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_60),
.B(n_63),
.Y(n_119)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_62),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_28),
.B(n_56),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_64),
.Y(n_139)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_65),
.Y(n_174)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_66),
.Y(n_188)
);

BUFx4f_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_67),
.Y(n_175)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_68),
.Y(n_183)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_69),
.Y(n_180)
);

BUFx4f_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_72),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_28),
.B(n_17),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_73),
.B(n_85),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx4f_ASAP7_75t_SL g179 ( 
.A(n_74),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_21),
.Y(n_75)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_75),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_28),
.B(n_16),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_76),
.B(n_84),
.Y(n_123)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_77),
.Y(n_172)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_80),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_81),
.Y(n_155)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_82),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_83),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_30),
.B(n_14),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_21),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_54),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_86),
.B(n_87),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_50),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_18),
.Y(n_91)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_51),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_92),
.B(n_104),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_41),
.B(n_14),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_94),
.B(n_13),
.Y(n_170)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_97),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_98),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

BUFx2_ASAP7_75t_R g143 ( 
.A(n_100),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_101),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

INVx6_ASAP7_75t_SL g104 ( 
.A(n_20),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_105),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_20),
.B(n_14),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_106),
.B(n_108),
.Y(n_186)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_107),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_40),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_19),
.Y(n_109)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

BUFx10_ASAP7_75t_L g110 ( 
.A(n_32),
.Y(n_110)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_110),
.Y(n_178)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_19),
.Y(n_112)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_112),
.Y(n_182)
);

BUFx16f_ASAP7_75t_L g113 ( 
.A(n_32),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_113),
.Y(n_138)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_32),
.Y(n_114)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_114),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_19),
.Y(n_115)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_115),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_62),
.A2(n_30),
.B1(n_53),
.B2(n_47),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_121),
.A2(n_130),
.B1(n_152),
.B2(n_160),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_72),
.A2(n_55),
.B1(n_52),
.B2(n_46),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_122),
.A2(n_146),
.B1(n_26),
.B2(n_55),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_109),
.A2(n_49),
.B1(n_56),
.B2(n_47),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_126),
.A2(n_127),
.B1(n_131),
.B2(n_133),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_112),
.A2(n_49),
.B1(n_56),
.B2(n_47),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_65),
.A2(n_53),
.B1(n_44),
.B2(n_42),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_91),
.A2(n_53),
.B1(n_44),
.B2(n_42),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_66),
.A2(n_44),
.B1(n_42),
.B2(n_30),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_68),
.B(n_37),
.C(n_24),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_137),
.B(n_83),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_103),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_140),
.B(n_147),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_106),
.A2(n_23),
.B1(n_52),
.B2(n_46),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_105),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_74),
.A2(n_23),
.B1(n_52),
.B2(n_46),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_75),
.B(n_22),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_158),
.B(n_168),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_100),
.A2(n_22),
.B1(n_38),
.B2(n_31),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_159),
.A2(n_161),
.B1(n_48),
.B2(n_178),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_79),
.A2(n_57),
.B1(n_93),
.B2(n_88),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_78),
.A2(n_22),
.B1(n_38),
.B2(n_31),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_89),
.A2(n_23),
.B1(n_38),
.B2(n_31),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_166),
.A2(n_26),
.B1(n_48),
.B2(n_43),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_67),
.B(n_55),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_170),
.B(n_13),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_113),
.B(n_36),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_173),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_113),
.B(n_36),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_184),
.B(n_83),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_175),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_190),
.Y(n_308)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_142),
.Y(n_191)
);

INVx3_ASAP7_75t_SL g264 ( 
.A(n_191),
.Y(n_264)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_192),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_123),
.B(n_70),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_193),
.B(n_197),
.Y(n_262)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_187),
.Y(n_194)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_194),
.Y(n_258)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_118),
.Y(n_195)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_195),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_176),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_196),
.B(n_199),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_137),
.B(n_70),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_198),
.A2(n_214),
.B1(n_223),
.B2(n_232),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_143),
.Y(n_199)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_142),
.Y(n_201)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_201),
.Y(n_261)
);

NAND2xp33_ASAP7_75t_SL g202 ( 
.A(n_143),
.B(n_173),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_202),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_203),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_150),
.Y(n_204)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_204),
.Y(n_270)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_206),
.Y(n_277)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_164),
.Y(n_207)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_207),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_165),
.B(n_67),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_208),
.B(n_246),
.Y(n_273)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_124),
.Y(n_210)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_210),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_211),
.Y(n_318)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_124),
.Y(n_213)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_213),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_186),
.A2(n_58),
.B1(n_64),
.B2(n_71),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_215),
.B(n_222),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_153),
.A2(n_26),
.B1(n_115),
.B2(n_98),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_216),
.A2(n_220),
.B1(n_241),
.B2(n_171),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_217),
.B(n_230),
.Y(n_297)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_162),
.Y(n_218)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_218),
.Y(n_287)
);

INVx4_ASAP7_75t_SL g219 ( 
.A(n_184),
.Y(n_219)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_219),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_153),
.A2(n_61),
.B1(n_29),
.B2(n_43),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_162),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_221),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_119),
.A2(n_69),
.B1(n_81),
.B2(n_95),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_177),
.B(n_90),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_224),
.Y(n_265)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_132),
.Y(n_225)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_225),
.Y(n_294)
);

INVx6_ASAP7_75t_SL g226 ( 
.A(n_138),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_226),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_164),
.B(n_29),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_228),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_134),
.B(n_99),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_183),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_229),
.Y(n_301)
);

AO22x1_ASAP7_75t_L g230 ( 
.A1(n_121),
.A2(n_130),
.B1(n_163),
.B2(n_116),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_141),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_231),
.B(n_237),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_117),
.A2(n_101),
.B1(n_102),
.B2(n_24),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_129),
.Y(n_233)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_233),
.Y(n_314)
);

AND2x4_ASAP7_75t_SL g234 ( 
.A(n_116),
.B(n_36),
.Y(n_234)
);

AND2x2_ASAP7_75t_SL g312 ( 
.A(n_234),
.B(n_249),
.Y(n_312)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_163),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_235),
.B(n_247),
.Y(n_302)
);

O2A1O1Ixp33_ASAP7_75t_L g236 ( 
.A1(n_135),
.A2(n_39),
.B(n_29),
.C(n_33),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_236),
.B(n_179),
.Y(n_266)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_129),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_117),
.A2(n_39),
.B1(n_33),
.B2(n_37),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_238),
.A2(n_240),
.B1(n_151),
.B2(n_157),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_172),
.B(n_39),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_244),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_132),
.A2(n_110),
.B1(n_43),
.B2(n_48),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_179),
.A2(n_37),
.B1(n_33),
.B2(n_24),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_242),
.A2(n_199),
.B1(n_219),
.B2(n_190),
.Y(n_299)
);

BUFx8_ASAP7_75t_L g243 ( 
.A(n_183),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_243),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_125),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_125),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_251),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_144),
.B(n_0),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_144),
.Y(n_247)
);

NAND2x1_ASAP7_75t_SL g248 ( 
.A(n_178),
.B(n_145),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_248),
.B(n_250),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_188),
.B(n_111),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_148),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_148),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_181),
.B(n_107),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_254),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_167),
.B(n_1),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_253),
.B(n_1),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_174),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_185),
.A2(n_110),
.B1(n_35),
.B2(n_3),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_255),
.B(n_2),
.Y(n_319)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_139),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_257),
.Y(n_279)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_139),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_189),
.A2(n_180),
.B1(n_174),
.B2(n_136),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_263),
.A2(n_275),
.B1(n_286),
.B2(n_291),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_266),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_189),
.A2(n_180),
.B1(n_136),
.B2(n_156),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_197),
.B(n_149),
.C(n_155),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_280),
.B(n_298),
.C(n_315),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_212),
.B(n_149),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_281),
.B(n_284),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_193),
.B(n_188),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_200),
.A2(n_156),
.B1(n_154),
.B2(n_169),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_212),
.B(n_120),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_289),
.B(n_307),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_217),
.A2(n_154),
.B1(n_169),
.B2(n_157),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_230),
.A2(n_179),
.B1(n_151),
.B2(n_171),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_293),
.A2(n_305),
.B1(n_309),
.B2(n_255),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_296),
.B(n_304),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_217),
.B(n_155),
.C(n_120),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_299),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_230),
.A2(n_223),
.B1(n_227),
.B2(n_219),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_203),
.A2(n_253),
.B1(n_246),
.B2(n_205),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_306),
.A2(n_273),
.B1(n_307),
.B2(n_284),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_208),
.B(n_145),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_234),
.A2(n_135),
.B1(n_128),
.B2(n_118),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_310),
.B(n_6),
.Y(n_373)
);

O2A1O1Ixp33_ASAP7_75t_SL g311 ( 
.A1(n_234),
.A2(n_128),
.B(n_118),
.C(n_35),
.Y(n_311)
);

A2O1A1O1Ixp25_ASAP7_75t_L g338 ( 
.A1(n_311),
.A2(n_234),
.B(n_243),
.C(n_248),
.D(n_249),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_206),
.B(n_35),
.C(n_2),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_209),
.B(n_231),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_316),
.B(n_317),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_247),
.B(n_1),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_319),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_196),
.B(n_2),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_320),
.B(n_190),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_266),
.A2(n_202),
.B(n_226),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_321),
.A2(n_329),
.B(n_338),
.Y(n_389)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_274),
.Y(n_324)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_324),
.Y(n_377)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_274),
.Y(n_326)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_326),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_262),
.B(n_207),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_327),
.B(n_328),
.C(n_341),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_262),
.B(n_280),
.C(n_298),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_290),
.A2(n_236),
.B(n_248),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_330),
.A2(n_367),
.B1(n_303),
.B2(n_311),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_265),
.B(n_251),
.Y(n_331)
);

OAI21xp33_ASAP7_75t_L g405 ( 
.A1(n_331),
.A2(n_347),
.B(n_349),
.Y(n_405)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_308),
.Y(n_333)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_333),
.Y(n_395)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_308),
.Y(n_334)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_334),
.Y(n_401)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_308),
.Y(n_337)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_337),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_313),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_339),
.B(n_348),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_297),
.A2(n_254),
.B1(n_244),
.B2(n_235),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_340),
.A2(n_352),
.B1(n_369),
.B2(n_370),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_273),
.B(n_250),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_344),
.B(n_282),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_263),
.A2(n_194),
.B1(n_233),
.B2(n_237),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_345),
.A2(n_346),
.B1(n_354),
.B2(n_357),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_275),
.A2(n_213),
.B1(n_210),
.B2(n_225),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_313),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_292),
.B(n_316),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_313),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_350),
.B(n_359),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_310),
.B(n_201),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_351),
.B(n_366),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_297),
.A2(n_249),
.B1(n_245),
.B2(n_191),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_258),
.Y(n_353)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_353),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_297),
.A2(n_245),
.B1(n_256),
.B2(n_257),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_289),
.B(n_221),
.C(n_204),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_355),
.B(n_356),
.C(n_312),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_297),
.B(n_243),
.C(n_211),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_300),
.A2(n_211),
.B1(n_192),
.B2(n_243),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_258),
.Y(n_358)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_358),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_302),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_300),
.A2(n_218),
.B1(n_195),
.B2(n_5),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_360),
.Y(n_379)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_302),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_361),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_290),
.A2(n_299),
.B(n_288),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_362),
.A2(n_303),
.B(n_279),
.Y(n_417)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_302),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_363),
.Y(n_414)
);

INVx5_ASAP7_75t_L g364 ( 
.A(n_269),
.Y(n_364)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_364),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_313),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_365),
.Y(n_383)
);

O2A1O1Ixp33_ASAP7_75t_L g366 ( 
.A1(n_288),
.A2(n_311),
.B(n_304),
.C(n_306),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_264),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_272),
.B(n_3),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_368),
.B(n_373),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_305),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_278),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_278),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_371),
.A2(n_293),
.B1(n_296),
.B2(n_277),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_292),
.B(n_6),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_374),
.B(n_320),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_381),
.B(n_404),
.C(n_408),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_331),
.Y(n_382)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_382),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_384),
.A2(n_386),
.B1(n_399),
.B2(n_407),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_330),
.A2(n_319),
.B1(n_286),
.B2(n_268),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_385),
.A2(n_390),
.B1(n_403),
.B2(n_416),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_344),
.A2(n_335),
.B1(n_323),
.B2(n_371),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_347),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_387),
.B(n_393),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_335),
.A2(n_268),
.B1(n_272),
.B2(n_276),
.Y(n_390)
);

OAI21xp33_ASAP7_75t_SL g452 ( 
.A1(n_391),
.A2(n_357),
.B(n_322),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_342),
.A2(n_276),
.B1(n_281),
.B2(n_267),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_396),
.A2(n_417),
.B(n_338),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_364),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_397),
.B(n_398),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_364),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_335),
.A2(n_312),
.B1(n_309),
.B2(n_317),
.Y(n_399)
);

OAI32xp33_ASAP7_75t_L g402 ( 
.A1(n_372),
.A2(n_271),
.A3(n_267),
.B1(n_277),
.B2(n_302),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_402),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_370),
.A2(n_291),
.B1(n_271),
.B2(n_312),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_328),
.B(n_312),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_406),
.B(n_368),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_323),
.A2(n_366),
.B1(n_332),
.B2(n_343),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_341),
.B(n_279),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g409 ( 
.A(n_327),
.B(n_315),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_409),
.B(n_412),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g412 ( 
.A(n_332),
.B(n_295),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_324),
.B(n_295),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_413),
.B(n_420),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_366),
.A2(n_362),
.B1(n_326),
.B2(n_340),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_359),
.B(n_282),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_423),
.A2(n_430),
.B(n_399),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_379),
.A2(n_339),
.B1(n_348),
.B2(n_372),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_424),
.A2(n_439),
.B1(n_443),
.B2(n_448),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_377),
.B(n_351),
.Y(n_426)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_426),
.Y(n_462)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_415),
.Y(n_428)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_428),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_389),
.A2(n_321),
.B(n_338),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_390),
.B(n_349),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_431),
.B(n_441),
.Y(n_467)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_413),
.Y(n_433)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_433),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_378),
.B(n_325),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_436),
.B(n_360),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_377),
.B(n_361),
.Y(n_437)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_437),
.Y(n_474)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_415),
.Y(n_438)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_438),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_388),
.A2(n_325),
.B1(n_336),
.B2(n_363),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_418),
.Y(n_440)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_440),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_405),
.B(n_374),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_378),
.B(n_356),
.C(n_355),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_442),
.B(n_449),
.C(n_458),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_388),
.A2(n_336),
.B1(n_329),
.B2(n_345),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_394),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_444),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_420),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_445),
.B(n_446),
.Y(n_461)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_418),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_394),
.B(n_322),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_447),
.B(n_450),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_386),
.A2(n_369),
.B1(n_352),
.B2(n_354),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_404),
.B(n_353),
.C(n_358),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_382),
.B(n_301),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_451),
.B(n_454),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_452),
.A2(n_417),
.B1(n_379),
.B2(n_419),
.Y(n_478)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_395),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_453),
.B(n_455),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_392),
.B(n_393),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_387),
.B(n_373),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_392),
.B(n_337),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_456),
.B(n_410),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_408),
.B(n_314),
.C(n_259),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_407),
.A2(n_346),
.B1(n_334),
.B2(n_333),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_459),
.A2(n_376),
.B1(n_411),
.B2(n_383),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_381),
.B(n_314),
.C(n_260),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_460),
.B(n_409),
.C(n_383),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_434),
.A2(n_416),
.B1(n_385),
.B2(n_406),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_466),
.A2(n_470),
.B1(n_469),
.B2(n_485),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_434),
.A2(n_376),
.B1(n_403),
.B2(n_389),
.Y(n_470)
);

FAx1_ASAP7_75t_SL g471 ( 
.A(n_430),
.B(n_412),
.CI(n_375),
.CON(n_471),
.SN(n_471)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_471),
.B(n_435),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_472),
.B(n_475),
.C(n_481),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_429),
.B(n_375),
.C(n_414),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_476),
.A2(n_485),
.B1(n_489),
.B2(n_494),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_478),
.A2(n_482),
.B(n_427),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_435),
.B(n_402),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g513 ( 
.A(n_479),
.B(n_449),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_429),
.B(n_380),
.C(n_396),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_421),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_484),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_422),
.A2(n_411),
.B1(n_384),
.B2(n_397),
.Y(n_485)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_486),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_487),
.B(n_490),
.C(n_423),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_436),
.B(n_401),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_488),
.B(n_491),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_422),
.A2(n_398),
.B1(n_401),
.B2(n_395),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_460),
.B(n_260),
.C(n_410),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_439),
.B(n_261),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_425),
.B(n_400),
.Y(n_493)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_493),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_432),
.A2(n_445),
.B1(n_443),
.B2(n_433),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_432),
.A2(n_400),
.B1(n_367),
.B2(n_287),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_495),
.A2(n_453),
.B1(n_446),
.B2(n_440),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_497),
.A2(n_510),
.B1(n_512),
.B2(n_489),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g528 ( 
.A(n_499),
.B(n_524),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_503),
.B(n_504),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_465),
.B(n_442),
.Y(n_504)
);

INVxp67_ASAP7_75t_SL g505 ( 
.A(n_473),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_505),
.A2(n_506),
.B1(n_514),
.B2(n_515),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_494),
.A2(n_425),
.B1(n_448),
.B2(n_457),
.Y(n_506)
);

CKINVDCx16_ASAP7_75t_R g507 ( 
.A(n_493),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_507),
.B(n_483),
.Y(n_539)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_486),
.Y(n_508)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_508),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_478),
.A2(n_447),
.B(n_424),
.Y(n_509)
);

O2A1O1Ixp33_ASAP7_75t_L g541 ( 
.A1(n_509),
.A2(n_462),
.B(n_468),
.C(n_480),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_466),
.A2(n_457),
.B1(n_437),
.B2(n_459),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_511),
.A2(n_495),
.B(n_502),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_470),
.A2(n_455),
.B1(n_426),
.B2(n_427),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_513),
.B(n_517),
.Y(n_540)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_483),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_463),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_488),
.B(n_458),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_490),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_518),
.B(n_482),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_474),
.A2(n_456),
.B1(n_421),
.B2(n_438),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_519),
.A2(n_521),
.B1(n_522),
.B2(n_477),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_465),
.B(n_450),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_520),
.B(n_523),
.C(n_472),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_474),
.A2(n_428),
.B1(n_269),
.B2(n_318),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_475),
.B(n_287),
.C(n_270),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_491),
.B(n_261),
.Y(n_524)
);

A2O1A1O1Ixp25_ASAP7_75t_L g525 ( 
.A1(n_509),
.A2(n_471),
.B(n_479),
.C(n_484),
.D(n_467),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_525),
.B(n_529),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_526),
.A2(n_542),
.B1(n_547),
.B2(n_548),
.Y(n_558)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_527),
.Y(n_549)
);

A2O1A1O1Ixp25_ASAP7_75t_L g529 ( 
.A1(n_512),
.A2(n_471),
.B(n_514),
.C(n_500),
.D(n_508),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_532),
.B(n_531),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_504),
.B(n_481),
.C(n_487),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_533),
.B(n_535),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_506),
.A2(n_464),
.B1(n_462),
.B2(n_461),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_534),
.A2(n_545),
.B1(n_515),
.B2(n_522),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_518),
.B(n_464),
.C(n_461),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_536),
.B(n_539),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_537),
.Y(n_567)
);

A2O1A1Ixp33_ASAP7_75t_L g551 ( 
.A1(n_541),
.A2(n_511),
.B(n_519),
.C(n_510),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_SL g542 ( 
.A(n_500),
.B(n_468),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_523),
.B(n_463),
.C(n_477),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_543),
.B(n_546),
.C(n_531),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_501),
.B(n_492),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_544),
.B(n_496),
.Y(n_561)
);

OAI321xp33_ASAP7_75t_L g545 ( 
.A1(n_502),
.A2(n_492),
.A3(n_480),
.B1(n_294),
.B2(n_285),
.C(n_283),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_498),
.B(n_270),
.C(n_294),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g547 ( 
.A(n_501),
.B(n_285),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_497),
.A2(n_269),
.B1(n_318),
.B2(n_283),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_543),
.Y(n_550)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_550),
.Y(n_572)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_551),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_552),
.B(n_525),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_532),
.B(n_498),
.C(n_520),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_553),
.B(n_556),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_530),
.A2(n_515),
.B1(n_516),
.B2(n_513),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_557),
.A2(n_538),
.B1(n_548),
.B2(n_542),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_546),
.B(n_517),
.C(n_503),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_559),
.B(n_563),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_561),
.A2(n_529),
.B1(n_9),
.B2(n_10),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_536),
.B(n_496),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_562),
.B(n_568),
.Y(n_571)
);

A2O1A1O1Ixp25_ASAP7_75t_L g564 ( 
.A1(n_541),
.A2(n_264),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g575 ( 
.A1(n_564),
.A2(n_547),
.B(n_544),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_533),
.B(n_264),
.C(n_7),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_565),
.B(n_566),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_540),
.B(n_535),
.C(n_537),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_SL g568 ( 
.A(n_540),
.B(n_6),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_552),
.B(n_526),
.C(n_527),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_570),
.B(n_573),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_553),
.B(n_538),
.C(n_534),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_560),
.B(n_528),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_574),
.B(n_577),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_575),
.B(n_580),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_555),
.B(n_528),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_578),
.B(n_568),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_SL g589 ( 
.A(n_579),
.B(n_565),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_562),
.B(n_7),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_581),
.B(n_582),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_559),
.B(n_554),
.C(n_566),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_561),
.B(n_9),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_585),
.B(n_9),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_570),
.B(n_549),
.C(n_567),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_586),
.B(n_592),
.Y(n_603)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_583),
.A2(n_567),
.B(n_555),
.Y(n_587)
);

OAI21x1_ASAP7_75t_SL g606 ( 
.A1(n_587),
.A2(n_597),
.B(n_584),
.Y(n_606)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_588),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_589),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_SL g592 ( 
.A1(n_569),
.A2(n_558),
.B(n_551),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_SL g601 ( 
.A(n_593),
.B(n_596),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_582),
.B(n_564),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_572),
.A2(n_11),
.B(n_12),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_573),
.B(n_11),
.C(n_12),
.Y(n_598)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_598),
.B(n_581),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_599),
.B(n_600),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_594),
.A2(n_579),
.B1(n_580),
.B2(n_576),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_SL g602 ( 
.A1(n_587),
.A2(n_586),
.B(n_590),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_L g608 ( 
.A1(n_602),
.A2(n_590),
.B1(n_591),
.B2(n_595),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_SL g610 ( 
.A1(n_606),
.A2(n_597),
.B1(n_598),
.B2(n_585),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_608),
.A2(n_610),
.B(n_602),
.Y(n_611)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_603),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_609),
.B(n_601),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_611),
.A2(n_612),
.B(n_613),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_609),
.B(n_605),
.C(n_604),
.Y(n_612)
);

O2A1O1Ixp33_ASAP7_75t_L g615 ( 
.A1(n_612),
.A2(n_607),
.B(n_599),
.C(n_571),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_615),
.B(n_571),
.C(n_11),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_L g617 ( 
.A(n_616),
.B(n_614),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_617),
.B(n_11),
.Y(n_618)
);


endmodule