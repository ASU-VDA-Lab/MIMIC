module fake_jpeg_517_n_510 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_510);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_510;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_29),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_55),
.B(n_61),
.Y(n_133)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_56),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_58),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_59),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_17),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_60),
.B(n_94),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_17),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_62),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_63),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_49),
.B(n_16),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_66),
.B(n_70),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_67),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_69),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_35),
.B(n_16),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_22),
.B(n_0),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_71),
.B(n_76),
.Y(n_127)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_72),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_73),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_75),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_22),
.B(n_2),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx4_ASAP7_75t_SL g128 ( 
.A(n_78),
.Y(n_128)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_79),
.Y(n_186)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_80),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_81),
.Y(n_176)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_83),
.Y(n_173)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_84),
.Y(n_151)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_85),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_25),
.B(n_3),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_86),
.B(n_88),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g182 ( 
.A(n_87),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_25),
.B(n_3),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_37),
.B(n_4),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_101),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_90),
.Y(n_181)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_93),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_37),
.B(n_4),
.Y(n_94)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_95),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_96),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_27),
.B(n_15),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_97),
.B(n_105),
.Y(n_184)
);

BUFx12_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_99),
.Y(n_202)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_46),
.Y(n_100)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_100),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_41),
.B(n_44),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_102),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_103),
.Y(n_177)
);

INVx4_ASAP7_75t_SL g104 ( 
.A(n_36),
.Y(n_104)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_27),
.B(n_15),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g106 ( 
.A(n_30),
.Y(n_106)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_106),
.Y(n_162)
);

BUFx4f_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_107),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_108),
.Y(n_170)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_109),
.Y(n_172)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_36),
.Y(n_110)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_110),
.Y(n_175)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_46),
.Y(n_111)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_111),
.Y(n_179)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_44),
.Y(n_112)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_112),
.Y(n_185)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_36),
.Y(n_113)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_113),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_114),
.Y(n_189)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_115),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_36),
.Y(n_116)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_116),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_47),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_117),
.A2(n_113),
.B1(n_116),
.B2(n_118),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_47),
.Y(n_118)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_118),
.Y(n_201)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_23),
.Y(n_119)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_119),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_50),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_4),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_75),
.A2(n_19),
.B1(n_45),
.B2(n_43),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_123),
.A2(n_125),
.B1(n_150),
.B2(n_160),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_57),
.A2(n_19),
.B1(n_45),
.B2(n_43),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_88),
.B(n_18),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_136),
.B(n_144),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_64),
.A2(n_52),
.B1(n_50),
.B2(n_18),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_141),
.A2(n_142),
.B1(n_145),
.B2(n_148),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_104),
.A2(n_52),
.B1(n_26),
.B2(n_21),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_62),
.B(n_26),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_65),
.A2(n_21),
.B1(n_30),
.B2(n_32),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_147),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_119),
.A2(n_32),
.B1(n_24),
.B2(n_23),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_77),
.A2(n_24),
.B1(n_23),
.B2(n_7),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_149),
.A2(n_194),
.B1(n_148),
.B2(n_161),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_69),
.A2(n_24),
.B1(n_6),
.B2(n_7),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_87),
.B(n_15),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_155),
.B(n_163),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_73),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_156),
.A2(n_161),
.B1(n_178),
.B2(n_180),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_83),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_107),
.A2(n_10),
.B1(n_12),
.B2(n_15),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_87),
.B(n_59),
.Y(n_163)
);

AO22x1_ASAP7_75t_L g164 ( 
.A1(n_100),
.A2(n_10),
.B1(n_12),
.B2(n_95),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_164),
.A2(n_188),
.B1(n_125),
.B2(n_147),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_90),
.A2(n_10),
.B1(n_103),
.B2(n_102),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_167),
.A2(n_168),
.B1(n_131),
.B2(n_143),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_80),
.B(n_85),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_169),
.B(n_193),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_82),
.A2(n_10),
.B1(n_84),
.B2(n_110),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_96),
.A2(n_99),
.B1(n_108),
.B2(n_114),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_120),
.B(n_78),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_117),
.A2(n_98),
.B1(n_106),
.B2(n_94),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_98),
.B(n_106),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_196),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_94),
.B(n_66),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_197),
.B(n_133),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_55),
.B(n_66),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_199),
.B(n_135),
.Y(n_267)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_146),
.Y(n_206)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_206),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_196),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_208),
.B(n_212),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_130),
.A2(n_165),
.B1(n_124),
.B2(n_137),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_209),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_210),
.A2(n_211),
.B1(n_214),
.B2(n_219),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_201),
.A2(n_172),
.B1(n_185),
.B2(n_170),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_203),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_213),
.B(n_223),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_122),
.A2(n_159),
.B1(n_154),
.B2(n_129),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_215),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_216),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_127),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_217),
.B(n_221),
.Y(n_279)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_166),
.Y(n_218)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_218),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_179),
.A2(n_190),
.B1(n_186),
.B2(n_168),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_195),
.Y(n_220)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_220),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_140),
.B(n_134),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_164),
.B(n_121),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_222),
.B(n_246),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_128),
.Y(n_223)
);

INVx3_ASAP7_75t_SL g224 ( 
.A(n_146),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_224),
.Y(n_324)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_225),
.Y(n_282)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_171),
.Y(n_226)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_226),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_137),
.A2(n_139),
.B1(n_132),
.B2(n_198),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_227),
.A2(n_256),
.B1(n_269),
.B2(n_272),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_158),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_228),
.B(n_234),
.Y(n_284)
);

INVx4_ASAP7_75t_SL g230 ( 
.A(n_128),
.Y(n_230)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_230),
.Y(n_314)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_126),
.Y(n_231)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_231),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_158),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_175),
.Y(n_235)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_235),
.Y(n_313)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_174),
.Y(n_236)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_236),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_198),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_237),
.B(n_242),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_131),
.Y(n_238)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_238),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_239),
.A2(n_264),
.B1(n_273),
.B2(n_255),
.Y(n_296)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_143),
.Y(n_240)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_240),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_241),
.B(n_248),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_153),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_126),
.Y(n_243)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_243),
.Y(n_320)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_183),
.Y(n_244)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_244),
.Y(n_297)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_151),
.Y(n_245)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_245),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_142),
.B(n_187),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_174),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_247),
.B(n_249),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_203),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_176),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_171),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_250),
.B(n_251),
.Y(n_292)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_202),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_202),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_252),
.B(n_254),
.Y(n_304)
);

AND2x2_ASAP7_75t_SL g253 ( 
.A(n_151),
.B(n_191),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_253),
.Y(n_318)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_191),
.Y(n_254)
);

INVx8_ASAP7_75t_L g256 ( 
.A(n_152),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_152),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_257),
.B(n_267),
.Y(n_295)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_153),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_258),
.B(n_263),
.Y(n_311)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_200),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_259),
.B(n_261),
.Y(n_291)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_200),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_132),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_268),
.Y(n_293)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_173),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_145),
.A2(n_178),
.B1(n_181),
.B2(n_192),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_173),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_265),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_182),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_266),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_182),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_139),
.A2(n_135),
.B1(n_176),
.B2(n_162),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_181),
.A2(n_192),
.B1(n_162),
.B2(n_157),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_207),
.B(n_264),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_182),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_271),
.B(n_223),
.Y(n_308)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_157),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_138),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_230),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_210),
.A2(n_138),
.B1(n_177),
.B2(n_232),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_275),
.A2(n_290),
.B1(n_317),
.B2(n_216),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_283),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_232),
.A2(n_177),
.B1(n_222),
.B2(n_246),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_296),
.A2(n_305),
.B1(n_247),
.B2(n_224),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_301),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_239),
.A2(n_205),
.B1(n_229),
.B2(n_233),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_205),
.B(n_217),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_307),
.B(n_319),
.C(n_321),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_308),
.B(n_322),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_253),
.B(n_221),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_309),
.B(n_261),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_270),
.A2(n_253),
.B1(n_251),
.B2(n_252),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_235),
.B(n_244),
.C(n_215),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_260),
.B(n_220),
.Y(n_321)
);

AOI32xp33_ASAP7_75t_L g322 ( 
.A1(n_225),
.A2(n_254),
.A3(n_236),
.B1(n_250),
.B2(n_226),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_284),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_325),
.B(n_328),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_326),
.A2(n_299),
.B1(n_280),
.B2(n_282),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_327),
.B(n_360),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_311),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_306),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_329),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_288),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_330),
.B(n_352),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_296),
.A2(n_265),
.B1(n_263),
.B2(n_240),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_331),
.A2(n_332),
.B1(n_344),
.B2(n_346),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_286),
.A2(n_238),
.B1(n_272),
.B2(n_256),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_313),
.Y(n_333)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_333),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_279),
.B(n_245),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_334),
.B(n_335),
.Y(n_363)
);

OAI32xp33_ASAP7_75t_L g335 ( 
.A1(n_286),
.A2(n_218),
.A3(n_262),
.B1(n_259),
.B2(n_242),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_279),
.B(n_206),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_337),
.B(n_354),
.Y(n_364)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_292),
.Y(n_340)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_340),
.Y(n_372)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_313),
.Y(n_341)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_341),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_309),
.A2(n_228),
.B(n_234),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_342),
.A2(n_345),
.B(n_351),
.Y(n_366)
);

XNOR2x1_ASAP7_75t_SL g343 ( 
.A(n_321),
.B(n_307),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_343),
.A2(n_323),
.B(n_320),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_281),
.A2(n_274),
.B(n_249),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_312),
.A2(n_290),
.B1(n_305),
.B2(n_283),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_298),
.Y(n_347)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_347),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_295),
.B(n_315),
.Y(n_348)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_348),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_275),
.A2(n_312),
.B1(n_318),
.B2(n_281),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_349),
.A2(n_344),
.B1(n_346),
.B2(n_332),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_312),
.A2(n_302),
.B1(n_317),
.B2(n_278),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_285),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_291),
.A2(n_301),
.B1(n_293),
.B2(n_287),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_353),
.A2(n_356),
.B(n_349),
.Y(n_386)
);

OAI32xp33_ASAP7_75t_L g354 ( 
.A1(n_291),
.A2(n_293),
.A3(n_319),
.B1(n_304),
.B2(n_276),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_314),
.B(n_323),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_355),
.B(n_359),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_316),
.A2(n_310),
.B1(n_306),
.B2(n_297),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_298),
.Y(n_357)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_357),
.Y(n_392)
);

INVx4_ASAP7_75t_L g358 ( 
.A(n_303),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_276),
.B(n_297),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_300),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_324),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_L g378 ( 
.A1(n_361),
.A2(n_362),
.B1(n_280),
.B2(n_289),
.Y(n_378)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_300),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_343),
.B(n_320),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_367),
.B(n_381),
.C(n_382),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_329),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_370),
.B(n_371),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_329),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_373),
.B(n_389),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_336),
.A2(n_277),
.B1(n_303),
.B2(n_324),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_375),
.Y(n_399)
);

A2O1A1Ixp33_ASAP7_75t_SL g376 ( 
.A1(n_336),
.A2(n_294),
.B(n_277),
.C(n_289),
.Y(n_376)
);

AO22x1_ASAP7_75t_SL g415 ( 
.A1(n_376),
.A2(n_333),
.B1(n_341),
.B2(n_358),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_378),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_379),
.A2(n_388),
.B1(n_357),
.B2(n_362),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_338),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_380),
.B(n_334),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_343),
.B(n_282),
.C(n_299),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_350),
.B(n_294),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_386),
.B(n_358),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_350),
.B(n_327),
.C(n_342),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_331),
.A2(n_339),
.B1(n_338),
.B2(n_337),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_391),
.A2(n_356),
.B1(n_359),
.B2(n_347),
.Y(n_410)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_393),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_368),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_394),
.B(n_398),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_380),
.B(n_354),
.Y(n_395)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_395),
.Y(n_421)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_387),
.Y(n_396)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_396),
.Y(n_432)
);

CKINVDCx14_ASAP7_75t_R g398 ( 
.A(n_390),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_365),
.B(n_353),
.Y(n_400)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_400),
.Y(n_436)
);

CKINVDCx14_ASAP7_75t_R g402 ( 
.A(n_366),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_402),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_366),
.A2(n_345),
.B(n_339),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_403),
.A2(n_404),
.B(n_405),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_384),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_363),
.A2(n_335),
.B(n_351),
.Y(n_405)
);

FAx1_ASAP7_75t_SL g406 ( 
.A(n_389),
.B(n_326),
.CI(n_328),
.CON(n_406),
.SN(n_406)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_406),
.B(n_400),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_365),
.B(n_340),
.Y(n_407)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_407),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_382),
.B(n_355),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_408),
.B(n_381),
.C(n_373),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_410),
.A2(n_379),
.B1(n_376),
.B2(n_386),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_411),
.A2(n_412),
.B1(n_413),
.B2(n_414),
.Y(n_441)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_387),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_392),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_388),
.A2(n_391),
.B1(n_364),
.B2(n_374),
.Y(n_414)
);

AOI22x1_ASAP7_75t_L g438 ( 
.A1(n_415),
.A2(n_376),
.B1(n_412),
.B2(n_413),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_417),
.A2(n_418),
.B1(n_376),
.B2(n_371),
.Y(n_434)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_392),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_364),
.A2(n_348),
.B1(n_360),
.B2(n_361),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_419),
.A2(n_363),
.B1(n_374),
.B2(n_372),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_408),
.B(n_367),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_420),
.B(n_424),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_426),
.A2(n_439),
.B1(n_393),
.B2(n_411),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_428),
.A2(n_429),
.B1(n_434),
.B2(n_401),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_410),
.A2(n_414),
.B1(n_405),
.B2(n_419),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_409),
.B(n_372),
.C(n_383),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_431),
.B(n_433),
.C(n_435),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_409),
.B(n_375),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_397),
.B(n_369),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g437 ( 
.A(n_397),
.B(n_376),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_437),
.B(n_417),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_438),
.A2(n_415),
.B1(n_396),
.B2(n_385),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_395),
.A2(n_370),
.B1(n_369),
.B2(n_377),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_440),
.B(n_404),
.Y(n_450)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_442),
.Y(n_463)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_422),
.Y(n_443)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_443),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_441),
.A2(n_417),
.B1(n_402),
.B2(n_403),
.Y(n_445)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_445),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_447),
.B(n_437),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_426),
.A2(n_417),
.B1(n_407),
.B2(n_398),
.Y(n_448)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_448),
.Y(n_466)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_422),
.Y(n_449)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_449),
.Y(n_467)
);

CKINVDCx14_ASAP7_75t_R g468 ( 
.A(n_450),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g451 ( 
.A(n_439),
.Y(n_451)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_451),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_421),
.A2(n_417),
.B1(n_399),
.B2(n_394),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_452),
.B(n_454),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_435),
.B(n_406),
.C(n_418),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_453),
.B(n_431),
.C(n_425),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_430),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_455),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_421),
.A2(n_406),
.B1(n_401),
.B2(n_416),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_456),
.B(n_457),
.Y(n_460)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_430),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_458),
.B(n_427),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_461),
.B(n_453),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_469),
.B(n_455),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_470),
.B(n_433),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_472),
.B(n_474),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_468),
.A2(n_458),
.B1(n_436),
.B2(n_454),
.Y(n_473)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_473),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_460),
.B(n_444),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_475),
.B(n_476),
.C(n_478),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_470),
.B(n_446),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_463),
.A2(n_442),
.B1(n_429),
.B2(n_457),
.Y(n_477)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_477),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_459),
.B(n_446),
.C(n_444),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_463),
.A2(n_456),
.B1(n_448),
.B2(n_449),
.Y(n_479)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_479),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_480),
.B(n_481),
.C(n_482),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_471),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_462),
.B(n_425),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_478),
.B(n_459),
.C(n_460),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_487),
.B(n_491),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_481),
.A2(n_464),
.B(n_423),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_489),
.A2(n_466),
.B(n_452),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_480),
.B(n_471),
.C(n_464),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_485),
.A2(n_484),
.B1(n_486),
.B2(n_488),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_492),
.B(n_490),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_493),
.A2(n_494),
.B(n_495),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_483),
.B(n_469),
.Y(n_494)
);

NOR2xp67_ASAP7_75t_L g495 ( 
.A(n_490),
.B(n_474),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_487),
.A2(n_438),
.B1(n_466),
.B2(n_428),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_496),
.B(n_438),
.C(n_434),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_498),
.A2(n_499),
.B(n_500),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_497),
.B(n_475),
.Y(n_500)
);

A2O1A1Ixp33_ASAP7_75t_L g503 ( 
.A1(n_501),
.A2(n_443),
.B(n_467),
.C(n_465),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_503),
.Y(n_505)
);

NOR3xp33_ASAP7_75t_SL g504 ( 
.A(n_502),
.B(n_432),
.C(n_492),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_504),
.B(n_377),
.C(n_385),
.Y(n_506)
);

OAI21xp33_ASAP7_75t_L g507 ( 
.A1(n_506),
.A2(n_505),
.B(n_445),
.Y(n_507)
);

NOR3xp33_ASAP7_75t_L g508 ( 
.A(n_507),
.B(n_424),
.C(n_406),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_508),
.B(n_461),
.C(n_447),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_509),
.A2(n_420),
.B(n_415),
.Y(n_510)
);


endmodule