module fake_netlist_1_12488_n_513 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_513);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_513;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g76 ( .A(n_15), .Y(n_76) );
BUFx5_ASAP7_75t_L g77 ( .A(n_60), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_42), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_4), .Y(n_79) );
NOR2xp67_ASAP7_75t_L g80 ( .A(n_67), .B(n_61), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_28), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_30), .Y(n_82) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_2), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_20), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_65), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_23), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_9), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_23), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_53), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_71), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_11), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_40), .Y(n_92) );
INVx2_ASAP7_75t_SL g93 ( .A(n_68), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_8), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_51), .Y(n_95) );
INVxp33_ASAP7_75t_L g96 ( .A(n_38), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_63), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_22), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_21), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_27), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_54), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_8), .Y(n_102) );
INVxp33_ASAP7_75t_SL g103 ( .A(n_15), .Y(n_103) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_58), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_75), .Y(n_105) );
INVxp67_ASAP7_75t_SL g106 ( .A(n_45), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_57), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_48), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_25), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_20), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_35), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_34), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_3), .Y(n_113) );
INVxp67_ASAP7_75t_SL g114 ( .A(n_16), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_44), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_36), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_112), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_76), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_93), .B(n_0), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_93), .B(n_0), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_78), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_78), .Y(n_122) );
INVx4_ASAP7_75t_L g123 ( .A(n_104), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_79), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_81), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_77), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_96), .B(n_1), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_94), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_103), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_77), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_104), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_77), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_115), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_76), .B(n_1), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_88), .B(n_2), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_81), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_85), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_83), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_126), .Y(n_139) );
NAND2xp33_ASAP7_75t_L g140 ( .A(n_126), .B(n_77), .Y(n_140) );
INVx4_ASAP7_75t_L g141 ( .A(n_135), .Y(n_141) );
INVxp67_ASAP7_75t_L g142 ( .A(n_118), .Y(n_142) );
INVx4_ASAP7_75t_L g143 ( .A(n_135), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_121), .B(n_82), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_123), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_131), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_126), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_121), .B(n_122), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_122), .B(n_82), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_131), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_135), .B(n_88), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_126), .Y(n_152) );
INVxp67_ASAP7_75t_L g153 ( .A(n_118), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_123), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_134), .B(n_84), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_130), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_131), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_125), .B(n_100), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_135), .B(n_84), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_130), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_130), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_130), .Y(n_162) );
INVx4_ASAP7_75t_L g163 ( .A(n_135), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_142), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_141), .Y(n_165) );
INVx1_ASAP7_75t_SL g166 ( .A(n_155), .Y(n_166) );
HB1xp67_ASAP7_75t_L g167 ( .A(n_142), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_153), .B(n_133), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_153), .B(n_133), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_155), .B(n_125), .Y(n_170) );
NOR3xp33_ASAP7_75t_SL g171 ( .A(n_144), .B(n_117), .C(n_138), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_141), .Y(n_172) );
HB1xp67_ASAP7_75t_L g173 ( .A(n_155), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_141), .Y(n_174) );
BUFx5_ASAP7_75t_L g175 ( .A(n_139), .Y(n_175) );
NOR2xp33_ASAP7_75t_R g176 ( .A(n_140), .B(n_117), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_141), .Y(n_177) );
NOR2x1p5_ASAP7_75t_L g178 ( .A(n_141), .B(n_129), .Y(n_178) );
BUFx2_ASAP7_75t_L g179 ( .A(n_143), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_143), .Y(n_180) );
BUFx2_ASAP7_75t_L g181 ( .A(n_143), .Y(n_181) );
OAI22xp5_ASAP7_75t_L g182 ( .A1(n_143), .A2(n_124), .B1(n_128), .B2(n_137), .Y(n_182) );
INVxp67_ASAP7_75t_L g183 ( .A(n_148), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_143), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_148), .B(n_136), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_163), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_163), .B(n_136), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_163), .B(n_134), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g189 ( .A1(n_144), .A2(n_137), .B(n_134), .C(n_119), .Y(n_189) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_159), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_163), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_163), .Y(n_192) );
INVxp67_ASAP7_75t_SL g193 ( .A(n_139), .Y(n_193) );
BUFx4f_ASAP7_75t_L g194 ( .A(n_159), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_147), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_147), .Y(n_196) );
AOI21xp33_ASAP7_75t_L g197 ( .A1(n_164), .A2(n_128), .B(n_124), .Y(n_197) );
CKINVDCx8_ASAP7_75t_R g198 ( .A(n_190), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_183), .A2(n_159), .B1(n_151), .B2(n_158), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_195), .Y(n_200) );
BUFx10_ASAP7_75t_L g201 ( .A(n_167), .Y(n_201) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_189), .A2(n_159), .B(n_151), .C(n_158), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_188), .A2(n_159), .B1(n_151), .B2(n_149), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_188), .A2(n_151), .B1(n_149), .B2(n_140), .Y(n_204) );
NAND3xp33_ASAP7_75t_L g205 ( .A(n_168), .B(n_127), .C(n_161), .Y(n_205) );
INVx8_ASAP7_75t_L g206 ( .A(n_194), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_187), .A2(n_162), .B(n_161), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_175), .Y(n_208) );
BUFx12f_ASAP7_75t_L g209 ( .A(n_178), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_176), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_166), .B(n_151), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_169), .B(n_127), .Y(n_212) );
BUFx8_ASAP7_75t_SL g213 ( .A(n_194), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g214 ( .A1(n_194), .A2(n_119), .B1(n_120), .B2(n_156), .Y(n_214) );
OAI22xp5_ASAP7_75t_L g215 ( .A1(n_193), .A2(n_113), .B1(n_120), .B2(n_162), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_175), .B(n_152), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_179), .Y(n_217) );
BUFx12f_ASAP7_75t_L g218 ( .A(n_178), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_173), .B(n_114), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_179), .A2(n_160), .B1(n_156), .B2(n_152), .Y(n_220) );
CKINVDCx11_ASAP7_75t_R g221 ( .A(n_175), .Y(n_221) );
AND2x2_ASAP7_75t_L g222 ( .A(n_170), .B(n_160), .Y(n_222) );
AOI21x1_ASAP7_75t_L g223 ( .A1(n_195), .A2(n_132), .B(n_150), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_185), .B(n_132), .Y(n_224) );
INVxp67_ASAP7_75t_SL g225 ( .A(n_175), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_181), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_175), .B(n_145), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_175), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_196), .B(n_132), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_200), .Y(n_230) );
OR2x6_ASAP7_75t_L g231 ( .A(n_206), .B(n_181), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_221), .A2(n_215), .B1(n_197), .B2(n_206), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_199), .A2(n_182), .B1(n_196), .B2(n_175), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_222), .A2(n_175), .B1(n_171), .B2(n_186), .Y(n_234) );
BUFx8_ASAP7_75t_L g235 ( .A(n_209), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_222), .B(n_175), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_200), .Y(n_237) );
INVx3_ASAP7_75t_L g238 ( .A(n_208), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_206), .A2(n_192), .B1(n_191), .B2(n_186), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_214), .B(n_165), .Y(n_240) );
OAI21x1_ASAP7_75t_L g241 ( .A1(n_223), .A2(n_85), .B(n_105), .Y(n_241) );
AOI21xp33_ASAP7_75t_L g242 ( .A1(n_202), .A2(n_97), .B(n_105), .Y(n_242) );
OR2x2_ASAP7_75t_L g243 ( .A(n_211), .B(n_165), .Y(n_243) );
AOI22xp33_ASAP7_75t_SL g244 ( .A1(n_210), .A2(n_99), .B1(n_86), .B2(n_87), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_206), .A2(n_192), .B1(n_191), .B2(n_184), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_223), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_206), .A2(n_184), .B1(n_180), .B2(n_177), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_229), .Y(n_248) );
BUFx12f_ASAP7_75t_L g249 ( .A(n_201), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_219), .A2(n_180), .B1(n_177), .B2(n_174), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_214), .B(n_174), .Y(n_251) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_208), .Y(n_252) );
NAND2x1p5_ASAP7_75t_L g253 ( .A(n_228), .B(n_172), .Y(n_253) );
NAND3xp33_ASAP7_75t_SL g254 ( .A(n_210), .B(n_98), .C(n_91), .Y(n_254) );
AO22x1_ASAP7_75t_L g255 ( .A1(n_225), .A2(n_106), .B1(n_107), .B2(n_111), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_224), .B(n_172), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_228), .Y(n_257) );
AOI221xp5_ASAP7_75t_L g258 ( .A1(n_242), .A2(n_212), .B1(n_205), .B2(n_91), .C(n_110), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_232), .A2(n_218), .B1(n_209), .B2(n_213), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g260 ( .A1(n_254), .A2(n_218), .B1(n_217), .B2(n_226), .Y(n_260) );
AOI22xp5_ASAP7_75t_L g261 ( .A1(n_236), .A2(n_233), .B1(n_234), .B2(n_251), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_246), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_248), .B(n_224), .Y(n_263) );
CKINVDCx20_ASAP7_75t_R g264 ( .A(n_235), .Y(n_264) );
OAI221xp5_ASAP7_75t_L g265 ( .A1(n_244), .A2(n_203), .B1(n_198), .B2(n_204), .C(n_220), .Y(n_265) );
BUFx6f_ASAP7_75t_SL g266 ( .A(n_231), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_242), .A2(n_204), .B(n_203), .C(n_207), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_248), .A2(n_226), .B1(n_217), .B2(n_201), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_234), .A2(n_226), .B1(n_217), .B2(n_201), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_249), .A2(n_226), .B1(n_217), .B2(n_229), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_230), .B(n_217), .Y(n_271) );
AOI22xp33_ASAP7_75t_SL g272 ( .A1(n_249), .A2(n_226), .B1(n_198), .B2(n_87), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_230), .A2(n_227), .B1(n_216), .B2(n_86), .Y(n_273) );
OR2x6_ASAP7_75t_L g274 ( .A(n_231), .B(n_89), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_237), .B(n_132), .Y(n_275) );
AOI221xp5_ASAP7_75t_L g276 ( .A1(n_250), .A2(n_99), .B1(n_102), .B2(n_109), .C(n_110), .Y(n_276) );
OA21x2_ASAP7_75t_L g277 ( .A1(n_241), .A2(n_90), .B(n_92), .Y(n_277) );
OAI22xp5_ASAP7_75t_L g278 ( .A1(n_233), .A2(n_109), .B1(n_102), .B2(n_90), .Y(n_278) );
AO21x2_ASAP7_75t_L g279 ( .A1(n_246), .A2(n_108), .B(n_116), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g280 ( .A1(n_237), .A2(n_108), .B1(n_89), .B2(n_92), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_256), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_265), .A2(n_231), .B1(n_240), .B2(n_243), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_264), .Y(n_283) );
OAI211xp5_ASAP7_75t_L g284 ( .A1(n_272), .A2(n_80), .B(n_239), .C(n_245), .Y(n_284) );
NAND4xp25_ASAP7_75t_L g285 ( .A(n_276), .B(n_95), .C(n_101), .D(n_116), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_281), .B(n_255), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_262), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_274), .A2(n_231), .B1(n_255), .B2(n_243), .Y(n_288) );
AOI211xp5_ASAP7_75t_L g289 ( .A1(n_265), .A2(n_101), .B(n_95), .C(n_100), .Y(n_289) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_274), .Y(n_290) );
NOR2xp33_ASAP7_75t_R g291 ( .A(n_266), .B(n_235), .Y(n_291) );
NAND2xp33_ASAP7_75t_R g292 ( .A(n_274), .B(n_231), .Y(n_292) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_274), .Y(n_293) );
AND2x4_ASAP7_75t_L g294 ( .A(n_271), .B(n_238), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_274), .B(n_257), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_262), .Y(n_296) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_271), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_262), .Y(n_298) );
INVxp67_ASAP7_75t_SL g299 ( .A(n_281), .Y(n_299) );
AOI32xp33_ASAP7_75t_L g300 ( .A1(n_278), .A2(n_241), .A3(n_257), .B1(n_123), .B2(n_6), .Y(n_300) );
NAND2xp33_ASAP7_75t_SL g301 ( .A(n_266), .B(n_235), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_263), .B(n_235), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_263), .B(n_238), .Y(n_303) );
AOI22xp5_ASAP7_75t_L g304 ( .A1(n_266), .A2(n_247), .B1(n_238), .B2(n_253), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_297), .B(n_261), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_296), .B(n_261), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_296), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_298), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_298), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_287), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_282), .A2(n_266), .B1(n_278), .B2(n_258), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_287), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_299), .Y(n_313) );
OR2x2_ASAP7_75t_L g314 ( .A(n_295), .B(n_279), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_286), .B(n_258), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_295), .Y(n_316) );
OR2x2_ASAP7_75t_L g317 ( .A(n_290), .B(n_279), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_293), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_303), .B(n_279), .Y(n_319) );
NAND2x1_ASAP7_75t_SL g320 ( .A(n_288), .B(n_277), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_294), .Y(n_321) );
INVxp67_ASAP7_75t_SL g322 ( .A(n_292), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_301), .A2(n_259), .B1(n_276), .B2(n_260), .Y(n_323) );
OAI33xp33_ASAP7_75t_L g324 ( .A1(n_285), .A2(n_3), .A3(n_4), .B1(n_5), .B2(n_6), .B3(n_7), .Y(n_324) );
OAI31xp33_ASAP7_75t_L g325 ( .A1(n_284), .A2(n_267), .A3(n_302), .B(n_303), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_294), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_294), .B(n_277), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_294), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_288), .B(n_277), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_304), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_289), .B(n_277), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_291), .A2(n_280), .B1(n_269), .B2(n_270), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_304), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_312), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_329), .B(n_104), .Y(n_335) );
NAND3xp33_ASAP7_75t_L g336 ( .A(n_325), .B(n_300), .C(n_104), .Y(n_336) );
NAND3xp33_ASAP7_75t_L g337 ( .A(n_325), .B(n_313), .C(n_300), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_307), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_307), .B(n_275), .Y(n_339) );
AOI221xp5_ASAP7_75t_SL g340 ( .A1(n_323), .A2(n_104), .B1(n_268), .B2(n_273), .C(n_131), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_308), .Y(n_341) );
NOR2xp33_ASAP7_75t_R g342 ( .A(n_313), .B(n_283), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_309), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_312), .Y(n_344) );
AND2x4_ASAP7_75t_L g345 ( .A(n_321), .B(n_131), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_329), .B(n_77), .Y(n_346) );
AND2x4_ASAP7_75t_L g347 ( .A(n_321), .B(n_131), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_312), .Y(n_348) );
OAI22xp5_ASAP7_75t_SL g349 ( .A1(n_322), .A2(n_283), .B1(n_253), .B2(n_252), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_329), .B(n_77), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_309), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_316), .B(n_5), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_321), .B(n_77), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_310), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_316), .B(n_7), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_326), .B(n_77), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_326), .B(n_77), .Y(n_357) );
NAND2xp33_ASAP7_75t_R g358 ( .A(n_331), .B(n_9), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_310), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_306), .B(n_10), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_326), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_327), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_327), .B(n_131), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_327), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_305), .B(n_10), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_311), .A2(n_252), .B1(n_123), .B2(n_13), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_319), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_306), .B(n_11), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_305), .B(n_12), .Y(n_369) );
NAND2xp5_ASAP7_75t_SL g370 ( .A(n_322), .B(n_252), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_328), .Y(n_371) );
INVx3_ASAP7_75t_L g372 ( .A(n_328), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_306), .B(n_131), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_365), .B(n_324), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_367), .B(n_314), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_346), .B(n_319), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_363), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_338), .Y(n_378) );
INVxp67_ASAP7_75t_L g379 ( .A(n_358), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_365), .B(n_315), .Y(n_380) );
AOI22xp33_ASAP7_75t_SL g381 ( .A1(n_342), .A2(n_331), .B1(n_318), .B2(n_333), .Y(n_381) );
AOI221x1_ASAP7_75t_L g382 ( .A1(n_336), .A2(n_315), .B1(n_330), .B2(n_333), .C(n_319), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_362), .B(n_318), .Y(n_383) );
AOI321xp33_ASAP7_75t_L g384 ( .A1(n_366), .A2(n_323), .A3(n_330), .B1(n_332), .B2(n_305), .C(n_317), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_346), .B(n_318), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_337), .A2(n_332), .B1(n_317), .B2(n_314), .Y(n_386) );
O2A1O1Ixp33_ASAP7_75t_L g387 ( .A1(n_366), .A2(n_317), .B(n_314), .C(n_320), .Y(n_387) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_349), .B(n_320), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_334), .Y(n_389) );
NOR2x1_ASAP7_75t_L g390 ( .A(n_352), .B(n_123), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_334), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_341), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_346), .B(n_12), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_343), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_351), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_351), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_354), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_367), .B(n_13), .Y(n_398) );
INVx1_ASAP7_75t_SL g399 ( .A(n_363), .Y(n_399) );
AOI322xp5_ASAP7_75t_L g400 ( .A1(n_350), .A2(n_14), .A3(n_16), .B1(n_17), .B2(n_18), .C1(n_19), .C2(n_21), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_334), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_344), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_362), .B(n_14), .Y(n_403) );
OAI332xp33_ASAP7_75t_L g404 ( .A1(n_369), .A2(n_17), .A3(n_18), .B1(n_19), .B2(n_22), .B3(n_24), .C1(n_25), .C2(n_26), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_354), .Y(n_405) );
OAI22xp33_ASAP7_75t_SL g406 ( .A1(n_352), .A2(n_24), .B1(n_26), .B2(n_29), .Y(n_406) );
AND2x4_ASAP7_75t_L g407 ( .A(n_362), .B(n_31), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_344), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_344), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_371), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_371), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_364), .B(n_32), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_350), .B(n_252), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_355), .A2(n_33), .B1(n_37), .B2(n_39), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_355), .Y(n_415) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_350), .A2(n_157), .B1(n_150), .B2(n_146), .C(n_154), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_359), .Y(n_417) );
INVx1_ASAP7_75t_SL g418 ( .A(n_399), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_415), .B(n_335), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_381), .B(n_340), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_380), .B(n_335), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_378), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_379), .A2(n_360), .B1(n_368), .B2(n_340), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_383), .B(n_364), .Y(n_424) );
INVxp67_ASAP7_75t_L g425 ( .A(n_377), .Y(n_425) );
INVx1_ASAP7_75t_SL g426 ( .A(n_403), .Y(n_426) );
NOR3xp33_ASAP7_75t_SL g427 ( .A(n_374), .B(n_370), .C(n_339), .Y(n_427) );
NOR4xp25_ASAP7_75t_SL g428 ( .A(n_388), .B(n_361), .C(n_363), .D(n_373), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_386), .B(n_373), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_410), .Y(n_430) );
BUFx2_ASAP7_75t_L g431 ( .A(n_383), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_375), .B(n_359), .Y(n_432) );
NAND2xp33_ASAP7_75t_SL g433 ( .A(n_388), .B(n_353), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_375), .B(n_372), .Y(n_434) );
INVxp67_ASAP7_75t_L g435 ( .A(n_390), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_411), .B(n_376), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_404), .B(n_373), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_392), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_394), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_395), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_387), .B(n_384), .Y(n_441) );
XNOR2x1_ASAP7_75t_L g442 ( .A(n_403), .B(n_357), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_396), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_417), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_389), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_389), .B(n_372), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_397), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_391), .B(n_372), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_405), .Y(n_449) );
OAI32xp33_ASAP7_75t_L g450 ( .A1(n_398), .A2(n_372), .A3(n_357), .B1(n_356), .B2(n_353), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_385), .B(n_356), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_391), .B(n_401), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_401), .Y(n_453) );
AO22x2_ASAP7_75t_L g454 ( .A1(n_441), .A2(n_382), .B1(n_402), .B2(n_408), .Y(n_454) );
NOR3xp33_ASAP7_75t_L g455 ( .A(n_441), .B(n_406), .C(n_414), .Y(n_455) );
NAND3xp33_ASAP7_75t_L g456 ( .A(n_420), .B(n_400), .C(n_393), .Y(n_456) );
O2A1O1Ixp5_ASAP7_75t_L g457 ( .A1(n_433), .A2(n_407), .B(n_408), .C(n_409), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_433), .A2(n_407), .B1(n_412), .B2(n_413), .Y(n_458) );
NAND2xp33_ASAP7_75t_SL g459 ( .A(n_428), .B(n_407), .Y(n_459) );
OAI21xp5_ASAP7_75t_SL g460 ( .A1(n_420), .A2(n_412), .B(n_416), .Y(n_460) );
NAND3xp33_ASAP7_75t_L g461 ( .A(n_427), .B(n_409), .C(n_402), .Y(n_461) );
AOI221xp5_ASAP7_75t_L g462 ( .A1(n_437), .A2(n_347), .B1(n_345), .B2(n_348), .C(n_157), .Y(n_462) );
XOR2xp5_ASAP7_75t_L g463 ( .A(n_442), .B(n_347), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_429), .B(n_347), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_444), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_445), .Y(n_466) );
NOR2x1_ASAP7_75t_L g467 ( .A(n_431), .B(n_345), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_445), .Y(n_468) );
OAI21xp5_ASAP7_75t_SL g469 ( .A1(n_423), .A2(n_345), .B(n_41), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_453), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_418), .B(n_431), .Y(n_471) );
INVxp67_ASAP7_75t_L g472 ( .A(n_430), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_438), .Y(n_473) );
NOR2x1_ASAP7_75t_L g474 ( .A(n_442), .B(n_43), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_424), .B(n_46), .Y(n_475) );
NOR2x1_ASAP7_75t_L g476 ( .A(n_474), .B(n_422), .Y(n_476) );
AOI221xp5_ASAP7_75t_L g477 ( .A1(n_456), .A2(n_425), .B1(n_436), .B2(n_450), .C(n_435), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_463), .A2(n_426), .B1(n_421), .B2(n_419), .Y(n_478) );
INVxp67_ASAP7_75t_L g479 ( .A(n_471), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_467), .A2(n_424), .B1(n_451), .B2(n_432), .Y(n_480) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_465), .Y(n_481) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_455), .A2(n_450), .B(n_434), .C(n_447), .Y(n_482) );
AOI211xp5_ASAP7_75t_L g483 ( .A1(n_455), .A2(n_434), .B(n_439), .C(n_440), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_472), .Y(n_484) );
XNOR2xp5_ASAP7_75t_L g485 ( .A(n_454), .B(n_449), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_460), .A2(n_443), .B1(n_448), .B2(n_446), .Y(n_486) );
OAI222xp33_ASAP7_75t_L g487 ( .A1(n_458), .A2(n_452), .B1(n_49), .B2(n_50), .C1(n_52), .C2(n_55), .Y(n_487) );
NAND4xp25_ASAP7_75t_L g488 ( .A(n_462), .B(n_47), .C(n_56), .D(n_59), .Y(n_488) );
XNOR2x1_ASAP7_75t_L g489 ( .A(n_454), .B(n_62), .Y(n_489) );
AOI211xp5_ASAP7_75t_L g490 ( .A1(n_469), .A2(n_64), .B(n_66), .C(n_69), .Y(n_490) );
AND2x4_ASAP7_75t_L g491 ( .A(n_461), .B(n_70), .Y(n_491) );
OAI221xp5_ASAP7_75t_L g492 ( .A1(n_459), .A2(n_72), .B1(n_73), .B2(n_74), .C(n_145), .Y(n_492) );
NAND3xp33_ASAP7_75t_SL g493 ( .A(n_459), .B(n_145), .C(n_154), .Y(n_493) );
AOI322xp5_ASAP7_75t_L g494 ( .A1(n_464), .A2(n_473), .A3(n_454), .B1(n_470), .B2(n_466), .C1(n_468), .C2(n_475), .Y(n_494) );
OAI211xp5_ASAP7_75t_L g495 ( .A1(n_466), .A2(n_468), .B(n_470), .C(n_457), .Y(n_495) );
XNOR2xp5_ASAP7_75t_L g496 ( .A(n_457), .B(n_463), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_455), .A2(n_441), .B1(n_456), .B2(n_379), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_455), .A2(n_474), .B(n_459), .C(n_433), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_481), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g500 ( .A(n_497), .Y(n_500) );
BUFx2_ASAP7_75t_L g501 ( .A(n_498), .Y(n_501) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_484), .Y(n_502) );
O2A1O1Ixp33_ASAP7_75t_L g503 ( .A1(n_493), .A2(n_482), .B(n_492), .C(n_483), .Y(n_503) );
NAND3xp33_ASAP7_75t_SL g504 ( .A(n_490), .B(n_477), .C(n_494), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_500), .A2(n_496), .B1(n_489), .B2(n_485), .Y(n_505) );
OAI21x1_ASAP7_75t_L g506 ( .A1(n_502), .A2(n_476), .B(n_480), .Y(n_506) );
NOR3xp33_ASAP7_75t_L g507 ( .A(n_501), .B(n_487), .C(n_488), .Y(n_507) );
INVx1_ASAP7_75t_SL g508 ( .A(n_505), .Y(n_508) );
XNOR2xp5_ASAP7_75t_L g509 ( .A(n_507), .B(n_504), .Y(n_509) );
OAI22xp33_ASAP7_75t_L g510 ( .A1(n_508), .A2(n_502), .B1(n_499), .B2(n_486), .Y(n_510) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_509), .Y(n_511) );
AOI222xp33_ASAP7_75t_L g512 ( .A1(n_511), .A2(n_509), .B1(n_506), .B2(n_479), .C1(n_495), .C2(n_491), .Y(n_512) );
AOI221xp5_ASAP7_75t_L g513 ( .A1(n_512), .A2(n_510), .B1(n_503), .B2(n_478), .C(n_491), .Y(n_513) );
endmodule