module fake_netlist_1_8344_n_22 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_22);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_22;
wire n_20;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
wire n_7;
HB1xp67_ASAP7_75t_L g7 ( .A(n_1), .Y(n_7) );
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_5), .Y(n_8) );
CKINVDCx20_ASAP7_75t_R g9 ( .A(n_2), .Y(n_9) );
INVx2_ASAP7_75t_SL g10 ( .A(n_0), .Y(n_10) );
BUFx2_ASAP7_75t_L g11 ( .A(n_7), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_7), .B(n_6), .Y(n_12) );
INVx3_ASAP7_75t_L g13 ( .A(n_10), .Y(n_13) );
OR2x2_ASAP7_75t_L g14 ( .A(n_10), .B(n_0), .Y(n_14) );
BUFx6f_ASAP7_75t_L g15 ( .A(n_13), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_11), .B(n_8), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_16), .B(n_12), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
AOI221xp5_ASAP7_75t_SL g19 ( .A1(n_18), .A2(n_15), .B1(n_14), .B2(n_9), .C(n_13), .Y(n_19) );
BUFx3_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
OAI22xp5_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_22) );
endmodule