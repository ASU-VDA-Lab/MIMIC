module fake_jpeg_12025_n_140 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_140);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_140;

wire n_117;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_3),
.B(n_0),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_28),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g29 ( 
.A(n_12),
.B(n_3),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_29),
.B(n_40),
.Y(n_58)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_30),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_24),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_31),
.B(n_33),
.Y(n_65)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_32),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_5),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_10),
.B(n_5),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_43),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_11),
.B(n_5),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_47),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_45),
.Y(n_70)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_24),
.B(n_23),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_11),
.B(n_6),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_50),
.A2(n_56),
.B1(n_9),
.B2(n_32),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_10),
.B(n_6),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_17),
.B(n_7),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_53),
.A2(n_55),
.B1(n_19),
.B2(n_26),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_17),
.B(n_7),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_54),
.B(n_53),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_29),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_74),
.Y(n_95)
);

AOI32xp33_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_19),
.A3(n_23),
.B1(n_15),
.B2(n_14),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_73),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_27),
.A2(n_9),
.B1(n_52),
.B2(n_36),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_79),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_28),
.A2(n_38),
.B1(n_39),
.B2(n_51),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_48),
.A2(n_40),
.B1(n_27),
.B2(n_46),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_50),
.B(n_56),
.C(n_45),
.Y(n_89)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_90),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_89),
.A2(n_95),
.B1(n_75),
.B2(n_67),
.Y(n_108)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_94),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_65),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_93),
.B(n_96),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_77),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_58),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_62),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_62),
.B(n_66),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_106),
.B(n_69),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_101),
.B(n_98),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_95),
.B(n_89),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_57),
.C(n_70),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_70),
.C(n_77),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_83),
.A2(n_88),
.B(n_98),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_87),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_111),
.B(n_113),
.Y(n_123)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_118),
.Y(n_124)
);

AND2x6_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_64),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_106),
.A2(n_69),
.B1(n_67),
.B2(n_81),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_108),
.B1(n_103),
.B2(n_67),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_117),
.A2(n_119),
.B(n_99),
.Y(n_121)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_SL g129 ( 
.A1(n_121),
.A2(n_122),
.B(n_115),
.C(n_107),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_104),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_125),
.A2(n_105),
.B(n_96),
.Y(n_127)
);

OAI321xp33_ASAP7_75t_L g126 ( 
.A1(n_123),
.A2(n_102),
.A3(n_113),
.B1(n_117),
.B2(n_119),
.C(n_101),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_127),
.Y(n_131)
);

AO221x1_ASAP7_75t_L g128 ( 
.A1(n_120),
.A2(n_115),
.B1(n_60),
.B2(n_78),
.C(n_80),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_128),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_116),
.C(n_120),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_75),
.C(n_78),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_131),
.A2(n_124),
.B1(n_86),
.B2(n_84),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_133),
.A2(n_135),
.B1(n_132),
.B2(n_75),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_132),
.A2(n_90),
.B(n_60),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_71),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_136),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_137),
.B(n_72),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_72),
.Y(n_140)
);


endmodule