module fake_netlist_5_690_n_73 (n_16, n_0, n_12, n_9, n_18, n_22, n_1, n_8, n_10, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_20, n_5, n_14, n_2, n_13, n_3, n_6, n_73);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_22;
input n_1;
input n_8;
input n_10;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_20;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_73;

wire n_54;
wire n_29;
wire n_43;
wire n_47;
wire n_58;
wire n_67;
wire n_69;
wire n_36;
wire n_25;
wire n_53;
wire n_27;
wire n_42;
wire n_64;
wire n_45;
wire n_24;
wire n_46;
wire n_28;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_70;
wire n_38;
wire n_71;
wire n_61;
wire n_68;
wire n_72;
wire n_32;
wire n_35;
wire n_41;
wire n_65;
wire n_56;
wire n_51;
wire n_63;
wire n_57;
wire n_37;
wire n_59;
wire n_26;
wire n_30;
wire n_55;
wire n_33;
wire n_48;
wire n_31;
wire n_23;
wire n_50;
wire n_66;
wire n_52;
wire n_49;
wire n_60;
wire n_39;

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_8),
.B(n_15),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_1),
.A2(n_7),
.B1(n_3),
.B2(n_6),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_19),
.A2(n_3),
.B1(n_6),
.B2(n_10),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_2),
.B(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_0),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_29),
.A2(n_0),
.B1(n_5),
.B2(n_14),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

AOI221xp5_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_5),
.B1(n_18),
.B2(n_23),
.C(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_37),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_35),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_25),
.B(n_32),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_24),
.B(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_47),
.B(n_25),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_25),
.B(n_30),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_50),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_44),
.B(n_39),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_26),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_26),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_40),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_42),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_40),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_58),
.B(n_62),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_64),
.B1(n_66),
.B2(n_65),
.Y(n_68)
);

NOR2xp67_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_53),
.Y(n_69)
);

NOR3xp33_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_33),
.C(n_41),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_25),
.B(n_43),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_28),
.B(n_34),
.Y(n_72)
);

OR2x6_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_28),
.Y(n_73)
);


endmodule