module fake_jpeg_17980_n_115 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_115);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_115;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_3),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_57),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_51),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_1),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_1),
.Y(n_63)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_64),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_68),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_49),
.B(n_45),
.C(n_43),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_53),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_71),
.Y(n_80)
);

CKINVDCx12_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_52),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_50),
.Y(n_71)
);

INVx2_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_73),
.A2(n_52),
.B1(n_40),
.B2(n_41),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_75),
.A2(n_6),
.B1(n_11),
.B2(n_12),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_67),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_76),
.B(n_81),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_40),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_84),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_2),
.Y(n_84)
);

INVxp33_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_65),
.B1(n_44),
.B2(n_4),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_86),
.A2(n_88),
.B1(n_82),
.B2(n_79),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_88)
);

AOI32xp33_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_44),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_80),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_92),
.A2(n_75),
.B1(n_6),
.B2(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_95),
.Y(n_102)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_93),
.Y(n_99)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_89),
.C(n_14),
.Y(n_100)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_13),
.B(n_16),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_17),
.B(n_18),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_103),
.A2(n_21),
.B(n_23),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_104),
.B(n_102),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_107),
.C(n_105),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_24),
.C(n_25),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_86),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_78),
.Y(n_111)
);

OAI21x1_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_27),
.B(n_28),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_112),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_30),
.B(n_32),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_34),
.B(n_35),
.Y(n_115)
);


endmodule