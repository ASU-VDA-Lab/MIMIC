module fake_jpeg_8364_n_53 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_53);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_53;

wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_32;

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

AOI32xp33_ASAP7_75t_L g30 ( 
.A1(n_24),
.A2(n_10),
.A3(n_21),
.B1(n_20),
.B2(n_4),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_15),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_27),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_31)
);

AOI22x1_ASAP7_75t_SL g37 ( 
.A1(n_31),
.A2(n_5),
.B1(n_9),
.B2(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_13),
.Y(n_40)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_2),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_36),
.B(n_37),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_33),
.B(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_28),
.A2(n_23),
.B1(n_6),
.B2(n_8),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_41),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_16),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_29),
.A2(n_18),
.B(n_22),
.Y(n_43)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_38),
.C(n_39),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_50),
.B(n_47),
.Y(n_51)
);

NOR3xp33_ASAP7_75t_SL g52 ( 
.A(n_51),
.B(n_43),
.C(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_49),
.Y(n_53)
);


endmodule