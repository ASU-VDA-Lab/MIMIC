module real_aes_3819_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_963, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_963;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_792;
wire n_673;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_952;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_260;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_955;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_958;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_961;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_960;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_925;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_936;
wire n_610;
wire n_581;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_142;
wire n_947;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_957;
wire n_296;
wire n_702;
wire n_954;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_193;
wire n_293;
wire n_162;
wire n_397;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_928;
wire n_155;
wire n_637;
wire n_243;
wire n_899;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_922;
wire n_149;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_959;
wire n_715;
wire n_134;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_949;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
NAND2xp5_ASAP7_75t_L g597 ( .A(n_0), .B(n_172), .Y(n_597) );
CKINVDCx5p33_ASAP7_75t_R g611 ( .A(n_1), .Y(n_611) );
INVx1_ASAP7_75t_L g271 ( .A(n_2), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_SL g668 ( .A1(n_3), .A2(n_140), .B(n_669), .C(n_670), .Y(n_668) );
OAI22xp33_ASAP7_75t_L g602 ( .A1(n_4), .A2(n_84), .B1(n_122), .B2(n_131), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_5), .B(n_121), .Y(n_247) );
INVxp67_ASAP7_75t_L g540 ( .A(n_6), .Y(n_540) );
INVx1_ASAP7_75t_L g569 ( .A(n_6), .Y(n_569) );
INVx1_ASAP7_75t_L g573 ( .A(n_6), .Y(n_573) );
BUFx2_ASAP7_75t_L g959 ( .A(n_6), .Y(n_959) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_7), .B(n_249), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_8), .A2(n_37), .B1(n_120), .B2(n_233), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_9), .A2(n_97), .B1(n_425), .B2(n_426), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_9), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_9), .A2(n_425), .B1(n_426), .B2(n_549), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_10), .A2(n_43), .B1(n_155), .B2(n_182), .Y(n_181) );
AOI22xp5_ASAP7_75t_L g300 ( .A1(n_11), .A2(n_66), .B1(n_190), .B2(n_293), .Y(n_300) );
INVx1_ASAP7_75t_L g265 ( .A(n_12), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g629 ( .A(n_13), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_14), .A2(n_73), .B1(n_131), .B2(n_184), .Y(n_660) );
CKINVDCx5p33_ASAP7_75t_R g699 ( .A(n_15), .Y(n_699) );
INVx1_ASAP7_75t_L g269 ( .A(n_16), .Y(n_269) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_17), .A2(n_64), .B1(n_122), .B2(n_136), .Y(n_659) );
CKINVDCx5p33_ASAP7_75t_R g945 ( .A(n_18), .Y(n_945) );
OA21x2_ASAP7_75t_L g145 ( .A1(n_19), .A2(n_72), .B(n_146), .Y(n_145) );
OA21x2_ASAP7_75t_L g195 ( .A1(n_19), .A2(n_72), .B(n_146), .Y(n_195) );
OAI21xp5_ASAP7_75t_L g105 ( .A1(n_20), .A2(n_106), .B(n_546), .Y(n_105) );
INVx1_ASAP7_75t_L g553 ( .A(n_20), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g292 ( .A1(n_21), .A2(n_69), .B1(n_190), .B2(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g262 ( .A(n_22), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g624 ( .A(n_23), .Y(n_624) );
BUFx8_ASAP7_75t_SL g560 ( .A(n_24), .Y(n_560) );
BUFx3_ASAP7_75t_L g942 ( .A(n_24), .Y(n_942) );
O2A1O1Ixp33_ASAP7_75t_L g674 ( .A1(n_25), .A2(n_299), .B(n_675), .C(n_676), .Y(n_674) );
OAI22xp33_ASAP7_75t_SL g600 ( .A1(n_26), .A2(n_49), .B1(n_122), .B2(n_157), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_27), .A2(n_35), .B1(n_157), .B2(n_245), .Y(n_589) );
AO22x1_ASAP7_75t_L g242 ( .A1(n_28), .A2(n_80), .B1(n_138), .B2(n_243), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_29), .Y(n_125) );
AND2x2_ASAP7_75t_L g154 ( .A(n_30), .B(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_31), .B(n_138), .Y(n_137) );
O2A1O1Ixp5_ASAP7_75t_L g640 ( .A1(n_32), .A2(n_140), .B(n_641), .C(n_642), .Y(n_640) );
INVx1_ASAP7_75t_L g545 ( .A(n_33), .Y(n_545) );
AOI22x1_ASAP7_75t_L g188 ( .A1(n_34), .A2(n_96), .B1(n_189), .B2(n_190), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_36), .B(n_193), .Y(n_235) );
AND2x2_ASAP7_75t_L g957 ( .A(n_38), .B(n_958), .Y(n_957) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_39), .B(n_593), .Y(n_592) );
CKINVDCx5p33_ASAP7_75t_R g643 ( .A(n_40), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_41), .B(n_166), .Y(n_165) );
OAI22xp5_ASAP7_75t_L g924 ( .A1(n_42), .A2(n_925), .B1(n_926), .B2(n_929), .Y(n_924) );
CKINVDCx5p33_ASAP7_75t_R g929 ( .A(n_42), .Y(n_929) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_44), .Y(n_559) );
CKINVDCx5p33_ASAP7_75t_R g672 ( .A(n_45), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_46), .B(n_214), .Y(n_213) );
AOI22xp5_ASAP7_75t_SL g926 ( .A1(n_47), .A2(n_74), .B1(n_927), .B2(n_928), .Y(n_926) );
INVx1_ASAP7_75t_L g928 ( .A(n_47), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_48), .B(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g146 ( .A(n_50), .Y(n_146) );
AND2x4_ASAP7_75t_L g142 ( .A(n_51), .B(n_143), .Y(n_142) );
AND2x4_ASAP7_75t_L g587 ( .A(n_51), .B(n_143), .Y(n_587) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_52), .Y(n_128) );
INVx2_ASAP7_75t_L g295 ( .A(n_53), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g609 ( .A(n_54), .Y(n_609) );
O2A1O1Ixp33_ASAP7_75t_L g626 ( .A1(n_55), .A2(n_140), .B(n_627), .C(n_628), .Y(n_626) );
CKINVDCx5p33_ASAP7_75t_R g648 ( .A(n_56), .Y(n_648) );
INVx2_ASAP7_75t_L g704 ( .A(n_57), .Y(n_704) );
CKINVDCx5p33_ASAP7_75t_R g608 ( .A(n_58), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_59), .A2(n_76), .B1(n_120), .B2(n_189), .Y(n_229) );
CKINVDCx14_ASAP7_75t_R g251 ( .A(n_60), .Y(n_251) );
AND2x2_ASAP7_75t_L g163 ( .A(n_61), .B(n_138), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_62), .B(n_206), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_63), .A2(n_82), .B1(n_183), .B2(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_65), .B(n_217), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g612 ( .A(n_67), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_68), .B(n_206), .Y(n_205) );
NAND2xp33_ASAP7_75t_R g662 ( .A(n_70), .B(n_195), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_70), .A2(n_100), .B1(n_257), .B2(n_593), .Y(n_710) );
NAND2x1p5_ASAP7_75t_L g167 ( .A(n_71), .B(n_150), .Y(n_167) );
INVx1_ASAP7_75t_L g927 ( .A(n_74), .Y(n_927) );
CKINVDCx14_ASAP7_75t_R g197 ( .A(n_75), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_77), .B(n_121), .Y(n_211) );
OR2x6_ASAP7_75t_L g542 ( .A(n_78), .B(n_543), .Y(n_542) );
AND3x1_ASAP7_75t_L g956 ( .A(n_78), .B(n_957), .C(n_959), .Y(n_956) );
CKINVDCx5p33_ASAP7_75t_R g703 ( .A(n_79), .Y(n_703) );
CKINVDCx5p33_ASAP7_75t_R g700 ( .A(n_81), .Y(n_700) );
INVx1_ASAP7_75t_L g544 ( .A(n_83), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_83), .B(n_545), .Y(n_955) );
INVx1_ASAP7_75t_L g958 ( .A(n_85), .Y(n_958) );
BUFx5_ASAP7_75t_L g122 ( .A(n_86), .Y(n_122) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_86), .Y(n_132) );
INVx1_ASAP7_75t_L g185 ( .A(n_86), .Y(n_185) );
INVx2_ASAP7_75t_L g680 ( .A(n_87), .Y(n_680) );
INVx2_ASAP7_75t_L g273 ( .A(n_88), .Y(n_273) );
INVx2_ASAP7_75t_L g631 ( .A(n_89), .Y(n_631) );
CKINVDCx5p33_ASAP7_75t_R g677 ( .A(n_90), .Y(n_677) );
NAND2xp33_ASAP7_75t_L g159 ( .A(n_91), .B(n_160), .Y(n_159) );
INVx2_ASAP7_75t_SL g143 ( .A(n_92), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_93), .B(n_130), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_94), .B(n_166), .Y(n_210) );
INVx1_ASAP7_75t_L g646 ( .A(n_95), .Y(n_646) );
CKINVDCx5p33_ASAP7_75t_R g426 ( .A(n_97), .Y(n_426) );
INVx2_ASAP7_75t_L g652 ( .A(n_98), .Y(n_652) );
OAI21xp33_ASAP7_75t_SL g622 ( .A1(n_99), .A2(n_122), .B(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_100), .B(n_593), .Y(n_694) );
INVxp67_ASAP7_75t_SL g724 ( .A(n_100), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_101), .A2(n_104), .B1(n_949), .B2(n_960), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_102), .B(n_148), .Y(n_147) );
OA21x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_560), .B(n_561), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_535), .Y(n_106) );
OAI22xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_424), .B1(n_427), .B2(n_533), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_424), .Y(n_108) );
NAND3xp33_ASAP7_75t_L g550 ( .A(n_109), .B(n_548), .C(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g534 ( .A(n_111), .B(n_428), .Y(n_534) );
NAND4xp25_ASAP7_75t_SL g111 ( .A(n_112), .B(n_315), .C(n_361), .D(n_393), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_253), .B(n_274), .Y(n_112) );
OAI21xp33_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_199), .B(n_220), .Y(n_113) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_114), .A2(n_373), .B1(n_377), .B2(n_379), .Y(n_372) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_176), .Y(n_115) );
INVx2_ASAP7_75t_L g305 ( .A(n_116), .Y(n_305) );
AND2x2_ASAP7_75t_L g422 ( .A(n_116), .B(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_152), .Y(n_116) );
AND2x2_ASAP7_75t_L g339 ( .A(n_117), .B(n_224), .Y(n_339) );
AND2x2_ASAP7_75t_L g389 ( .A(n_117), .B(n_359), .Y(n_389) );
NAND2x1_ASAP7_75t_L g416 ( .A(n_117), .B(n_178), .Y(n_416) );
OA21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_144), .B(n_147), .Y(n_117) );
OA21x2_ASAP7_75t_L g284 ( .A1(n_118), .A2(n_144), .B(n_147), .Y(n_284) );
OAI21x1_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_133), .B(n_141), .Y(n_118) );
OAI22xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_123), .B1(n_127), .B2(n_129), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g138 ( .A(n_122), .Y(n_138) );
INVx2_ASAP7_75t_L g191 ( .A(n_122), .Y(n_191) );
INVx2_ASAP7_75t_L g217 ( .A(n_122), .Y(n_217) );
AOI22xp33_ASAP7_75t_SL g607 ( .A1(n_122), .A2(n_157), .B1(n_608), .B2(n_609), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_122), .A2(n_136), .B1(n_611), .B2(n_612), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_122), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_122), .B(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_122), .B(n_648), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_122), .A2(n_157), .B1(n_699), .B2(n_700), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_126), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI22x1_ASAP7_75t_L g180 ( .A1(n_126), .A2(n_181), .B1(n_186), .B2(n_188), .Y(n_180) );
INVx4_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_127), .A2(n_210), .B(n_211), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_127), .B(n_227), .Y(n_226) );
OA22x2_ASAP7_75t_L g588 ( .A1(n_127), .A2(n_187), .B1(n_589), .B2(n_590), .Y(n_588) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_128), .Y(n_140) );
INVxp67_ASAP7_75t_L g161 ( .A(n_128), .Y(n_161) );
INVx1_ASAP7_75t_L g187 ( .A(n_128), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_128), .B(n_262), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_128), .B(n_265), .Y(n_264) );
INVx4_ASAP7_75t_L g268 ( .A(n_128), .Y(n_268) );
INVx3_ASAP7_75t_L g299 ( .A(n_128), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_128), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_128), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g136 ( .A(n_132), .Y(n_136) );
INVx6_ASAP7_75t_L g157 ( .A(n_132), .Y(n_157) );
INVx3_ASAP7_75t_L g215 ( .A(n_132), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_137), .B(n_139), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_135), .B(n_264), .Y(n_263) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_135), .A2(n_138), .B1(n_267), .B2(n_270), .Y(n_266) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g675 ( .A(n_136), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g702 ( .A1(n_136), .A2(n_245), .B1(n_703), .B2(n_704), .Y(n_702) );
INVxp67_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_SL g169 ( .A(n_140), .Y(n_169) );
INVx1_ASAP7_75t_L g218 ( .A(n_140), .Y(n_218) );
INVx1_ASAP7_75t_L g241 ( .A(n_140), .Y(n_241) );
OAI221xp5_ASAP7_75t_L g606 ( .A1(n_140), .A2(n_142), .B1(n_299), .B2(n_607), .C(n_610), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_140), .A2(n_268), .B1(n_659), .B2(n_660), .Y(n_658) );
OAI22xp33_ASAP7_75t_L g722 ( .A1(n_140), .A2(n_268), .B1(n_698), .B2(n_702), .Y(n_722) );
AO31x2_ASAP7_75t_L g179 ( .A1(n_141), .A2(n_180), .A3(n_192), .B(n_196), .Y(n_179) );
AO31x2_ASAP7_75t_L g286 ( .A1(n_141), .A2(n_180), .A3(n_192), .B(n_196), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_141), .B(n_585), .Y(n_721) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx3_ASAP7_75t_L g174 ( .A(n_142), .Y(n_174) );
INVx3_ASAP7_75t_L g228 ( .A(n_142), .Y(n_228) );
INVx1_ASAP7_75t_L g239 ( .A(n_142), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_142), .B(n_151), .Y(n_603) );
INVx3_ASAP7_75t_L g198 ( .A(n_144), .Y(n_198) );
BUFx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx4_ASAP7_75t_L g151 ( .A(n_145), .Y(n_151) );
INVx2_ASAP7_75t_L g207 ( .A(n_145), .Y(n_207) );
OR2x2_ASAP7_75t_L g238 ( .A(n_148), .B(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
OR2x2_ASAP7_75t_L g294 ( .A(n_149), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g172 ( .A(n_151), .Y(n_172) );
INVx2_ASAP7_75t_L g593 ( .A(n_151), .Y(n_593) );
NOR2xp33_ASAP7_75t_SL g679 ( .A(n_151), .B(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g341 ( .A(n_152), .B(n_286), .Y(n_341) );
AND2x2_ASAP7_75t_L g364 ( .A(n_152), .B(n_286), .Y(n_364) );
AND2x4_ASAP7_75t_L g410 ( .A(n_152), .B(n_283), .Y(n_410) );
AO21x2_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_162), .B(n_170), .Y(n_152) );
AO21x2_ASAP7_75t_L g280 ( .A1(n_153), .A2(n_162), .B(n_170), .Y(n_280) );
OAI21x1_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_158), .B(n_161), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_155), .B(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g160 ( .A(n_157), .Y(n_160) );
INVx1_ASAP7_75t_L g166 ( .A(n_157), .Y(n_166) );
INVx2_ASAP7_75t_SL g591 ( .A(n_157), .Y(n_591) );
INVx2_ASAP7_75t_L g671 ( .A(n_157), .Y(n_671) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g189 ( .A(n_160), .Y(n_189) );
OAI21x1_ASAP7_75t_SL g162 ( .A1(n_163), .A2(n_164), .B(n_168), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_165), .B(n_167), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_167), .B(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g175 ( .A(n_167), .Y(n_175) );
AOI21x1_ASAP7_75t_L g246 ( .A1(n_169), .A2(n_247), .B(n_248), .Y(n_246) );
AOI21xp33_ASAP7_75t_SL g170 ( .A1(n_171), .A2(n_173), .B(n_175), .Y(n_170) );
INVx2_ASAP7_75t_L g605 ( .A(n_171), .Y(n_605) );
OR2x2_ASAP7_75t_L g723 ( .A(n_171), .B(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_SL g678 ( .A(n_172), .B(n_649), .Y(n_678) );
NAND3xp33_ASAP7_75t_SL g291 ( .A(n_173), .B(n_258), .C(n_268), .Y(n_291) );
NAND3xp33_ASAP7_75t_L g297 ( .A(n_173), .B(n_258), .C(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NOR2x1_ASAP7_75t_L g219 ( .A(n_174), .B(n_206), .Y(n_219) );
INVx1_ASAP7_75t_L g303 ( .A(n_176), .Y(n_303) );
AND2x2_ASAP7_75t_L g488 ( .A(n_176), .B(n_410), .Y(n_488) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g252 ( .A(n_177), .Y(n_252) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g411 ( .A(n_178), .B(n_400), .Y(n_411) );
INVx1_ASAP7_75t_L g483 ( .A(n_178), .Y(n_483) );
AND2x2_ASAP7_75t_L g530 ( .A(n_178), .B(n_280), .Y(n_530) );
INVx3_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g469 ( .A(n_179), .B(n_332), .Y(n_469) );
INVx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g669 ( .A(n_183), .Y(n_669) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g245 ( .A(n_185), .Y(n_245) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_187), .B(n_227), .Y(n_231) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_195), .B(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g258 ( .A(n_195), .Y(n_258) );
BUFx3_ASAP7_75t_L g586 ( .A(n_195), .Y(n_586) );
INVx1_ASAP7_75t_L g620 ( .A(n_195), .Y(n_620) );
INVx1_ASAP7_75t_L g653 ( .A(n_195), .Y(n_653) );
NOR2xp67_ASAP7_75t_SL g196 ( .A(n_197), .B(n_198), .Y(n_196) );
OR2x2_ASAP7_75t_L g250 ( .A(n_198), .B(n_251), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_198), .A2(n_731), .B(n_732), .Y(n_730) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
OR2x2_ASAP7_75t_L g439 ( .A(n_202), .B(n_323), .Y(n_439) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g353 ( .A(n_203), .B(n_237), .Y(n_353) );
AND2x2_ASAP7_75t_L g385 ( .A(n_203), .B(n_289), .Y(n_385) );
INVx3_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g236 ( .A(n_204), .B(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g313 ( .A(n_204), .B(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g368 ( .A(n_204), .Y(n_368) );
AND2x4_ASAP7_75t_L g204 ( .A(n_205), .B(n_208), .Y(n_204) );
NOR2xp67_ASAP7_75t_L g661 ( .A(n_206), .B(n_239), .Y(n_661) );
INVx3_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_207), .B(n_273), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_207), .B(n_631), .Y(n_630) );
BUFx3_ASAP7_75t_L g650 ( .A(n_207), .Y(n_650) );
OAI21x1_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_212), .B(n_219), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_216), .B(n_218), .Y(n_212) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g234 ( .A(n_215), .Y(n_234) );
INVx1_ASAP7_75t_L g249 ( .A(n_215), .Y(n_249) );
INVx1_ASAP7_75t_L g627 ( .A(n_215), .Y(n_627) );
INVx1_ASAP7_75t_L g641 ( .A(n_215), .Y(n_641) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_218), .A2(n_625), .B1(n_649), .B2(n_697), .C(n_701), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_221), .B(n_252), .Y(n_220) );
INVx1_ASAP7_75t_L g486 ( .A(n_221), .Y(n_486) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_236), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g363 ( .A(n_223), .Y(n_363) );
INVx1_ASAP7_75t_L g406 ( .A(n_223), .Y(n_406) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g307 ( .A(n_224), .Y(n_307) );
AND2x2_ASAP7_75t_L g331 ( .A(n_224), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_224), .B(n_279), .Y(n_378) );
INVx2_ASAP7_75t_L g400 ( .A(n_224), .Y(n_400) );
NAND2x1p5_ASAP7_75t_L g224 ( .A(n_225), .B(n_230), .Y(n_224) );
AND2x2_ASAP7_75t_L g359 ( .A(n_225), .B(n_230), .Y(n_359) );
OR2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_229), .Y(n_225) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_235), .Y(n_230) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g293 ( .A(n_234), .Y(n_293) );
AND2x2_ASAP7_75t_L g287 ( .A(n_236), .B(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g325 ( .A(n_236), .Y(n_325) );
AND2x2_ASAP7_75t_L g335 ( .A(n_236), .B(n_336), .Y(n_335) );
INVx2_ASAP7_75t_SL g314 ( .A(n_237), .Y(n_314) );
OAI21x1_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_240), .B(n_250), .Y(n_237) );
OAI21xp5_ASAP7_75t_L g346 ( .A1(n_238), .A2(n_240), .B(n_250), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_239), .B(n_257), .Y(n_256) );
AOI21x1_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B(n_246), .Y(n_240) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g628 ( .A(n_245), .B(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_245), .B(n_677), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_249), .A2(n_268), .B1(n_645), .B2(n_647), .Y(n_644) );
OR2x2_ASAP7_75t_L g329 ( .A(n_252), .B(n_330), .Y(n_329) );
NAND3xp33_ASAP7_75t_L g527 ( .A(n_253), .B(n_528), .C(n_531), .Y(n_527) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g473 ( .A(n_254), .B(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g477 ( .A(n_254), .B(n_374), .Y(n_477) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g288 ( .A(n_255), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g311 ( .A(n_255), .Y(n_311) );
OR2x2_ASAP7_75t_L g345 ( .A(n_255), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g352 ( .A(n_255), .Y(n_352) );
AND2x2_ASAP7_75t_L g384 ( .A(n_255), .B(n_314), .Y(n_384) );
AO21x2_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_259), .B(n_272), .Y(n_255) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND3xp33_ASAP7_75t_SL g259 ( .A(n_260), .B(n_263), .C(n_266), .Y(n_259) );
NOR2xp33_ASAP7_75t_SL g267 ( .A(n_268), .B(n_269), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_268), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g625 ( .A(n_268), .Y(n_625) );
AOI31xp33_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_301), .A3(n_306), .B(n_308), .Y(n_274) );
INVx1_ASAP7_75t_L g316 ( .A(n_275), .Y(n_316) );
OAI21xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_281), .B(n_287), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g514 ( .A(n_278), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVxp67_ASAP7_75t_L g360 ( .A(n_280), .Y(n_360) );
INVx2_ASAP7_75t_L g392 ( .A(n_280), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_281), .B(n_306), .Y(n_318) );
OAI21xp33_ASAP7_75t_L g502 ( .A1(n_281), .A2(n_503), .B(n_504), .Y(n_502) );
INVx2_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
INVxp67_ASAP7_75t_SL g398 ( .A(n_283), .Y(n_398) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g332 ( .A(n_284), .Y(n_332) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x4_ASAP7_75t_L g391 ( .A(n_286), .B(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g321 ( .A(n_288), .B(n_322), .Y(n_321) );
NAND2x1_ASAP7_75t_SL g386 ( .A(n_288), .B(n_313), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_288), .B(n_374), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_288), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g518 ( .A(n_288), .Y(n_518) );
INVx2_ASAP7_75t_L g312 ( .A(n_289), .Y(n_312) );
AND2x2_ASAP7_75t_L g327 ( .A(n_289), .B(n_311), .Y(n_327) );
INVx1_ASAP7_75t_L g337 ( .A(n_289), .Y(n_337) );
NOR2x1_ASAP7_75t_L g351 ( .A(n_289), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g355 ( .A(n_289), .Y(n_355) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_289), .Y(n_371) );
INVx1_ASAP7_75t_L g438 ( .A(n_289), .Y(n_438) );
OR2x6_ASAP7_75t_L g289 ( .A(n_290), .B(n_296), .Y(n_289) );
OAI21x1_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_292), .B(n_294), .Y(n_290) );
NOR2xp67_ASAP7_75t_L g296 ( .A(n_297), .B(n_300), .Y(n_296) );
INVx3_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_299), .A2(n_602), .B(n_603), .Y(n_601) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g520 ( .A(n_305), .B(n_423), .Y(n_520) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_308), .A2(n_397), .B1(n_399), .B2(n_401), .Y(n_396) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_313), .Y(n_309) );
AND2x2_ASAP7_75t_L g402 ( .A(n_310), .B(n_374), .Y(n_402) );
AND2x2_ASAP7_75t_L g504 ( .A(n_310), .B(n_353), .Y(n_504) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
AND2x2_ASAP7_75t_L g354 ( .A(n_313), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g323 ( .A(n_314), .Y(n_323) );
INVx1_ASAP7_75t_L g474 ( .A(n_314), .Y(n_474) );
AOI221x1_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_317), .B1(n_319), .B2(n_328), .C(n_333), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_324), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_321), .A2(n_335), .B1(n_413), .B2(n_414), .Y(n_412) );
INVxp67_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
OR2x2_ASAP7_75t_L g420 ( .A(n_325), .B(n_336), .Y(n_420) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g419 ( .A(n_327), .B(n_353), .Y(n_419) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g446 ( .A(n_331), .Y(n_446) );
INVx1_ASAP7_75t_L g348 ( .A(n_332), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_332), .B(n_400), .Y(n_515) );
OAI221xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_338), .B1(n_342), .B2(n_347), .C(n_349), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_SL g379 ( .A(n_336), .B(n_380), .Y(n_379) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_336), .Y(n_485) );
OR2x2_ASAP7_75t_L g523 ( .A(n_336), .B(n_439), .Y(n_523) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g343 ( .A(n_337), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_339), .B(n_390), .Y(n_460) );
AND2x2_ASAP7_75t_L g482 ( .A(n_339), .B(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_339), .B(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g405 ( .A(n_340), .B(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_340), .B(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g347 ( .A(n_341), .B(n_348), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g381 ( .A1(n_341), .A2(n_382), .B1(n_386), .B2(n_387), .Y(n_381) );
INVxp67_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OAI21xp33_ASAP7_75t_L g451 ( .A1(n_343), .A2(n_452), .B(n_457), .Y(n_451) );
AND2x2_ASAP7_75t_L g408 ( .A(n_344), .B(n_371), .Y(n_408) );
INVx1_ASAP7_75t_L g511 ( .A(n_344), .Y(n_511) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g367 ( .A(n_345), .B(n_368), .Y(n_367) );
BUFx2_ASAP7_75t_L g456 ( .A(n_346), .Y(n_456) );
AND3x2_ASAP7_75t_L g356 ( .A(n_348), .B(n_357), .C(n_360), .Y(n_356) );
OR2x2_ASAP7_75t_L g377 ( .A(n_348), .B(n_378), .Y(n_377) );
OAI21xp5_ASAP7_75t_SL g349 ( .A1(n_350), .A2(n_354), .B(n_356), .Y(n_349) );
AND2x4_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
INVx2_ASAP7_75t_L g376 ( .A(n_351), .Y(n_376) );
INVx2_ASAP7_75t_L g380 ( .A(n_353), .Y(n_380) );
INVx1_ASAP7_75t_L g442 ( .A(n_353), .Y(n_442) );
AND2x2_ASAP7_75t_L g490 ( .A(n_355), .B(n_368), .Y(n_490) );
AND2x2_ASAP7_75t_L g432 ( .A(n_357), .B(n_391), .Y(n_432) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g415 ( .A(n_358), .B(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g423 ( .A(n_358), .Y(n_423) );
INVx2_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_360), .Y(n_395) );
AOI211xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_365), .B(n_372), .C(n_381), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_369), .Y(n_366) );
OAI221xp5_ASAP7_75t_SL g403 ( .A1(n_367), .A2(n_404), .B1(n_407), .B2(n_409), .C(n_412), .Y(n_403) );
INVxp67_ASAP7_75t_L g433 ( .A(n_367), .Y(n_433) );
INVx2_ASAP7_75t_L g374 ( .A(n_368), .Y(n_374) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_368), .Y(n_472) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_369), .Y(n_498) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
OR2x2_ASAP7_75t_L g522 ( .A(n_374), .B(n_376), .Y(n_522) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g503 ( .A(n_378), .Y(n_503) );
OR2x2_ASAP7_75t_L g517 ( .A(n_380), .B(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_384), .B(n_438), .Y(n_462) );
BUFx3_ASAP7_75t_L g491 ( .A(n_384), .Y(n_491) );
INVx2_ASAP7_75t_L g510 ( .A(n_385), .Y(n_510) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NOR2xp67_ASAP7_75t_SL g388 ( .A(n_389), .B(n_390), .Y(n_388) );
AND2x4_ASAP7_75t_L g457 ( .A(n_389), .B(n_391), .Y(n_457) );
INVx3_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
BUFx3_ASAP7_75t_L g480 ( .A(n_391), .Y(n_480) );
INVx1_ASAP7_75t_L g468 ( .A(n_392), .Y(n_468) );
NOR3xp33_ASAP7_75t_L g393 ( .A(n_394), .B(n_403), .C(n_417), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g413 ( .A(n_400), .B(n_410), .Y(n_413) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_406), .B(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g496 ( .A(n_406), .Y(n_496) );
INVx2_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
BUFx3_ASAP7_75t_L g450 ( .A(n_410), .Y(n_450) );
AND2x4_ASAP7_75t_SL g497 ( .A(n_410), .B(n_483), .Y(n_497) );
INVx2_ASAP7_75t_L g435 ( .A(n_411), .Y(n_435) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_416), .Y(n_525) );
AOI21xp33_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_420), .B(n_421), .Y(n_417) );
OAI222xp33_ASAP7_75t_L g463 ( .A1(n_418), .A2(n_464), .B1(n_470), .B2(n_475), .C1(n_479), .C2(n_481), .Y(n_463) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_426), .Y(n_549) );
INVx1_ASAP7_75t_L g551 ( .A(n_427), .Y(n_551) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_492), .Y(n_428) );
NOR4xp25_ASAP7_75t_L g429 ( .A(n_430), .B(n_447), .C(n_463), .D(n_484), .Y(n_429) );
NAND2xp5_ASAP7_75t_SL g430 ( .A(n_431), .B(n_440), .Y(n_430) );
AOI21xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_433), .B(n_434), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
OR2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_439), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g478 ( .A(n_438), .B(n_456), .Y(n_478) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_439), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_443), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OAI211xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_449), .B(n_451), .C(n_458), .Y(n_447) );
INVx2_ASAP7_75t_L g507 ( .A(n_450), .Y(n_507) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVxp67_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_461), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_465), .B(n_496), .Y(n_526) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NAND2x1p5_ASAP7_75t_L g466 ( .A(n_467), .B(n_469), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
INVx1_ASAP7_75t_L g532 ( .A(n_474), .Y(n_532) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OAI32xp33_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .A3(n_487), .B1(n_489), .B2(n_963), .Y(n_484) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
OAI221xp5_ASAP7_75t_L g524 ( .A1(n_489), .A2(n_509), .B1(n_525), .B2(n_526), .C(n_527), .Y(n_524) );
NAND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
AOI211x1_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_499), .B(n_501), .C(n_524), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_498), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
NAND2xp67_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND3xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_505), .C(n_512), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_508), .Y(n_505) );
INVxp67_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_516), .B1(n_519), .B2(n_521), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_523), .Y(n_521) );
INVxp67_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
OAI21xp5_ASAP7_75t_L g547 ( .A1(n_533), .A2(n_548), .B(n_550), .Y(n_547) );
INVxp67_ASAP7_75t_L g564 ( .A(n_533), .Y(n_564) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AO22x2_ASAP7_75t_L g931 ( .A1(n_534), .A2(n_568), .B1(n_932), .B2(n_936), .Y(n_931) );
CKINVDCx11_ASAP7_75t_R g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_537), .B(n_559), .Y(n_558) );
BUFx10_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_538), .Y(n_557) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
OR2x6_ASAP7_75t_L g572 ( .A(n_541), .B(n_573), .Y(n_572) );
INVx8_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g568 ( .A(n_542), .B(n_569), .Y(n_568) );
OR2x6_ASAP7_75t_L g948 ( .A(n_542), .B(n_569), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
AOI21xp5_ASAP7_75t_SL g546 ( .A1(n_547), .A2(n_552), .B(n_558), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx5_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g939 ( .A(n_558), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_930), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_563), .B(n_924), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_565), .B1(n_570), .B2(n_574), .Y(n_563) );
INVx4_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
BUFx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
BUFx8_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g935 ( .A(n_572), .Y(n_935) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx2_ASAP7_75t_SL g936 ( .A(n_575), .Y(n_936) );
AND2x4_ASAP7_75t_L g575 ( .A(n_576), .B(n_794), .Y(n_575) );
AND4x1_ASAP7_75t_L g576 ( .A(n_577), .B(n_742), .C(n_762), .D(n_774), .Y(n_576) );
AOI311xp33_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_632), .A3(n_663), .B(n_681), .C(n_715), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_614), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_581), .B(n_594), .Y(n_580) );
INVx3_ASAP7_75t_L g714 ( .A(n_581), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_581), .B(n_735), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_581), .B(n_766), .Y(n_765) );
AND2x2_ASAP7_75t_L g864 ( .A(n_581), .B(n_848), .Y(n_864) );
INVx3_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g753 ( .A(n_582), .B(n_685), .Y(n_753) );
INVx1_ASAP7_75t_L g816 ( .A(n_582), .Y(n_816) );
AND2x2_ASAP7_75t_L g858 ( .A(n_582), .B(n_604), .Y(n_858) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g834 ( .A(n_583), .Y(n_834) );
OAI21x1_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_588), .B(n_592), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_587), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g619 ( .A(n_587), .B(n_620), .Y(n_619) );
INVx4_ASAP7_75t_L g649 ( .A(n_587), .Y(n_649) );
INVx1_ASAP7_75t_L g731 ( .A(n_588), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_592), .Y(n_732) );
AND2x2_ASAP7_75t_L g845 ( .A(n_594), .B(n_714), .Y(n_845) );
INVx1_ASAP7_75t_SL g869 ( .A(n_594), .Y(n_869) );
AND2x2_ASAP7_75t_L g882 ( .A(n_594), .B(n_833), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_594), .B(n_683), .Y(n_883) );
AND2x4_ASAP7_75t_L g594 ( .A(n_595), .B(n_604), .Y(n_594) );
AND2x2_ASAP7_75t_L g766 ( .A(n_595), .B(n_617), .Y(n_766) );
INVx3_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g685 ( .A(n_596), .Y(n_685) );
NAND2xp33_ASAP7_75t_R g727 ( .A(n_596), .B(n_617), .Y(n_727) );
AND2x2_ASAP7_75t_L g735 ( .A(n_596), .B(n_604), .Y(n_735) );
INVx1_ASAP7_75t_L g806 ( .A(n_596), .Y(n_806) );
AND2x2_ASAP7_75t_L g848 ( .A(n_596), .B(n_617), .Y(n_848) );
HB1xp67_ASAP7_75t_L g875 ( .A(n_596), .Y(n_875) );
AND2x4_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_601), .Y(n_598) );
OR2x2_ASAP7_75t_L g729 ( .A(n_604), .B(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_L g815 ( .A(n_604), .B(n_816), .Y(n_815) );
OA21x2_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_606), .B(n_613), .Y(n_604) );
OA21x2_ASAP7_75t_L g687 ( .A1(n_605), .A2(n_606), .B(n_613), .Y(n_687) );
AND2x2_ASAP7_75t_L g878 ( .A(n_614), .B(n_859), .Y(n_878) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g887 ( .A(n_615), .B(n_825), .Y(n_887) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g734 ( .A(n_616), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g828 ( .A(n_616), .Y(n_828) );
AND2x2_ASAP7_75t_L g833 ( .A(n_616), .B(n_834), .Y(n_833) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
BUFx2_ASAP7_75t_L g683 ( .A(n_617), .Y(n_683) );
INVx2_ASAP7_75t_L g748 ( .A(n_617), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_617), .B(n_687), .Y(n_751) );
INVx1_ASAP7_75t_L g778 ( .A(n_617), .Y(n_778) );
OR2x2_ASAP7_75t_L g785 ( .A(n_617), .B(n_685), .Y(n_785) );
AND2x2_ASAP7_75t_L g819 ( .A(n_617), .B(n_820), .Y(n_819) );
INVx3_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AOI21x1_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_621), .B(n_630), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_625), .B(n_626), .Y(n_621) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
BUFx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_634), .B(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g802 ( .A(n_635), .B(n_739), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_654), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g910 ( .A(n_636), .B(n_693), .Y(n_910) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g789 ( .A(n_637), .B(n_656), .Y(n_789) );
AND2x2_ASAP7_75t_L g810 ( .A(n_637), .B(n_708), .Y(n_810) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
BUFx2_ASAP7_75t_R g690 ( .A(n_638), .Y(n_690) );
INVx2_ASAP7_75t_L g741 ( .A(n_638), .Y(n_741) );
AND2x2_ASAP7_75t_L g791 ( .A(n_638), .B(n_792), .Y(n_791) );
HB1xp67_ASAP7_75t_L g800 ( .A(n_638), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_638), .B(n_666), .Y(n_839) );
AND2x2_ASAP7_75t_L g844 ( .A(n_638), .B(n_760), .Y(n_844) );
AO21x2_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_650), .B(n_651), .Y(n_638) );
NOR3xp33_ASAP7_75t_L g639 ( .A(n_640), .B(n_644), .C(n_649), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g695 ( .A(n_650), .B(n_696), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AND2x4_ASAP7_75t_L g740 ( .A(n_655), .B(n_741), .Y(n_740) );
AND2x2_ASAP7_75t_L g913 ( .A(n_655), .B(n_760), .Y(n_913) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g719 ( .A(n_656), .B(n_720), .Y(n_719) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_656), .Y(n_757) );
INVx1_ASAP7_75t_L g792 ( .A(n_656), .Y(n_792) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_662), .Y(n_656) );
AND2x2_ASAP7_75t_L g709 ( .A(n_657), .B(n_710), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_661), .Y(n_657) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx2_ASAP7_75t_SL g809 ( .A(n_665), .Y(n_809) );
INVx1_ASAP7_75t_L g831 ( .A(n_665), .Y(n_831) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OR2x2_ASAP7_75t_L g692 ( .A(n_666), .B(n_693), .Y(n_692) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_666), .Y(n_711) );
INVx1_ASAP7_75t_L g718 ( .A(n_666), .Y(n_718) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_666), .Y(n_739) );
AND2x4_ASAP7_75t_L g744 ( .A(n_666), .B(n_720), .Y(n_744) );
INVx2_ASAP7_75t_L g760 ( .A(n_666), .Y(n_760) );
AND2x2_ASAP7_75t_L g770 ( .A(n_666), .B(n_693), .Y(n_770) );
AO31x2_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_673), .A3(n_678), .B(n_679), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI22xp33_ASAP7_75t_SL g681 ( .A1(n_682), .A2(n_688), .B1(n_705), .B2(n_712), .Y(n_681) );
NAND2x1p5_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
AND2x2_ASAP7_75t_L g713 ( .A(n_684), .B(n_714), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_684), .A2(n_763), .B1(n_767), .B2(n_773), .Y(n_762) );
AND2x4_ASAP7_75t_L g859 ( .A(n_684), .B(n_860), .Y(n_859) );
NAND2x1p5_ASAP7_75t_L g904 ( .A(n_684), .B(n_827), .Y(n_904) );
AND2x4_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
AND2x4_ASAP7_75t_L g825 ( .A(n_686), .B(n_730), .Y(n_825) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g820 ( .A(n_687), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_691), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AND2x4_ASAP7_75t_L g894 ( .A(n_691), .B(n_791), .Y(n_894) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g798 ( .A(n_692), .B(n_799), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_693), .B(n_741), .Y(n_761) );
AND2x2_ASAP7_75t_L g793 ( .A(n_693), .B(n_718), .Y(n_793) );
AND2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
AND2x2_ASAP7_75t_L g708 ( .A(n_695), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AOI21xp33_ASAP7_75t_L g917 ( .A1(n_705), .A2(n_918), .B(n_921), .Y(n_917) );
HB1xp67_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
OR2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_711), .Y(n_706) );
OR2x2_ASAP7_75t_L g880 ( .A(n_707), .B(n_718), .Y(n_880) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g901 ( .A(n_708), .Y(n_901) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g775 ( .A(n_714), .B(n_776), .Y(n_775) );
AND2x2_ASAP7_75t_L g852 ( .A(n_714), .B(n_735), .Y(n_852) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_725), .B1(n_733), .B2(n_736), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
AND2x4_ASAP7_75t_L g837 ( .A(n_719), .B(n_838), .Y(n_837) );
AND2x2_ASAP7_75t_L g843 ( .A(n_719), .B(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g781 ( .A(n_720), .Y(n_781) );
OAI21x1_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_722), .B(n_723), .Y(n_720) );
INVxp67_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_728), .B(n_827), .Y(n_826) );
AND2x2_ASAP7_75t_L g922 ( .A(n_728), .B(n_923), .Y(n_922) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g786 ( .A(n_729), .Y(n_786) );
NAND2xp33_ASAP7_75t_L g862 ( .A(n_733), .B(n_863), .Y(n_862) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
BUFx3_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_740), .Y(n_737) );
INVxp67_ASAP7_75t_L g854 ( .A(n_738), .Y(n_854) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g743 ( .A(n_740), .B(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_L g769 ( .A(n_740), .B(n_770), .Y(n_769) );
AND2x2_ASAP7_75t_L g776 ( .A(n_740), .B(n_777), .Y(n_776) );
AND2x2_ASAP7_75t_L g850 ( .A(n_740), .B(n_809), .Y(n_850) );
OAI31xp33_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_745), .A3(n_747), .B(n_749), .Y(n_742) );
INVx2_ASAP7_75t_L g754 ( .A(n_743), .Y(n_754) );
INVx2_ASAP7_75t_SL g772 ( .A(n_744), .Y(n_772) );
AND2x2_ASAP7_75t_L g788 ( .A(n_744), .B(n_789), .Y(n_788) );
AND2x2_ASAP7_75t_L g885 ( .A(n_744), .B(n_799), .Y(n_885) );
AND2x4_ASAP7_75t_L g905 ( .A(n_744), .B(n_791), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_744), .B(n_756), .Y(n_920) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
BUFx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
A2O1A1Ixp33_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_752), .B(n_754), .C(n_755), .Y(n_749) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
NOR2xp67_ASAP7_75t_L g805 ( .A(n_751), .B(n_806), .Y(n_805) );
OAI22xp33_ASAP7_75t_L g782 ( .A1(n_752), .A2(n_783), .B1(n_787), .B2(n_790), .Y(n_782) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g773 ( .A(n_755), .Y(n_773) );
OR2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_758), .Y(n_755) );
OR2x2_ASAP7_75t_L g771 ( .A(n_756), .B(n_772), .Y(n_771) );
AOI322xp5_ASAP7_75t_L g855 ( .A1(n_756), .A2(n_779), .A3(n_856), .B1(n_859), .B2(n_861), .C1(n_862), .C2(n_865), .Y(n_855) );
INVx2_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g916 ( .A(n_758), .Y(n_916) );
OR2x2_ASAP7_75t_L g758 ( .A(n_759), .B(n_761), .Y(n_758) );
INVx1_ASAP7_75t_L g892 ( .A(n_759), .Y(n_892) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g914 ( .A(n_761), .Y(n_914) );
INVxp67_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
BUFx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx2_ASAP7_75t_L g823 ( .A(n_766), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_768), .B(n_771), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
AND2x2_ASAP7_75t_L g865 ( .A(n_770), .B(n_791), .Y(n_865) );
INVx2_ASAP7_75t_L g871 ( .A(n_771), .Y(n_871) );
AOI21xp5_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_779), .B(n_782), .Y(n_774) );
INVx1_ASAP7_75t_L g841 ( .A(n_776), .Y(n_841) );
INVx1_ASAP7_75t_L g813 ( .A(n_777), .Y(n_813) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_778), .B(n_820), .Y(n_898) );
HB1xp67_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
NOR2xp33_ASAP7_75t_L g861 ( .A(n_780), .B(n_822), .Y(n_861) );
INVx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_784), .B(n_786), .Y(n_783) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx2_ASAP7_75t_L g923 ( .A(n_785), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_786), .A2(n_912), .B1(n_915), .B2(n_916), .Y(n_911) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
AND2x2_ASAP7_75t_L g891 ( .A(n_789), .B(n_892), .Y(n_891) );
OAI22xp5_ASAP7_75t_L g807 ( .A1(n_790), .A2(n_808), .B1(n_811), .B2(n_817), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_791), .B(n_793), .Y(n_790) );
INVx2_ASAP7_75t_SL g822 ( .A(n_791), .Y(n_822) );
NOR2xp67_ASAP7_75t_L g794 ( .A(n_795), .B(n_876), .Y(n_794) );
NAND4xp25_ASAP7_75t_L g795 ( .A(n_796), .B(n_835), .C(n_855), .D(n_866), .Y(n_795) );
NOR3xp33_ASAP7_75t_L g796 ( .A(n_797), .B(n_807), .C(n_821), .Y(n_796) );
AOI21xp33_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_801), .B(n_803), .Y(n_797) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
HB1xp67_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
BUFx2_ASAP7_75t_SL g804 ( .A(n_805), .Y(n_804) );
NAND2x1p5_ASAP7_75t_SL g808 ( .A(n_809), .B(n_810), .Y(n_808) );
INVx1_ASAP7_75t_L g829 ( .A(n_810), .Y(n_829) );
HB1xp67_ASAP7_75t_L g888 ( .A(n_810), .Y(n_888) );
INVxp33_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
NOR2x1_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .Y(n_812) );
INVx3_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
HB1xp67_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
OAI322xp33_ASAP7_75t_L g821 ( .A1(n_822), .A2(n_823), .A3(n_824), .B1(n_826), .B2(n_829), .C1(n_830), .C2(n_832), .Y(n_821) );
OR2x2_ASAP7_75t_L g853 ( .A(n_822), .B(n_854), .Y(n_853) );
INVx2_ASAP7_75t_L g836 ( .A(n_824), .Y(n_836) );
INVx2_ASAP7_75t_SL g824 ( .A(n_825), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_825), .B(n_848), .Y(n_847) );
INVx2_ASAP7_75t_L g870 ( .A(n_827), .Y(n_870) );
INVx2_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
OAI21xp33_ASAP7_75t_L g840 ( .A1(n_831), .A2(n_841), .B(n_842), .Y(n_840) );
INVx2_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx2_ASAP7_75t_L g860 ( .A(n_834), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_834), .B(n_875), .Y(n_874) );
AOI221x1_ASAP7_75t_L g835 ( .A1(n_836), .A2(n_837), .B1(n_840), .B2(n_845), .C(n_846), .Y(n_835) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
OR2x2_ASAP7_75t_L g900 ( .A(n_839), .B(n_901), .Y(n_900) );
INVx2_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
AOI21xp5_ASAP7_75t_L g877 ( .A1(n_843), .A2(n_878), .B(n_879), .Y(n_877) );
OAI22xp5_ASAP7_75t_L g846 ( .A1(n_847), .A2(n_849), .B1(n_851), .B2(n_853), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_848), .B(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_850), .A2(n_867), .B1(n_871), .B2(n_872), .Y(n_866) );
OAI221xp5_ASAP7_75t_SL g906 ( .A1(n_851), .A2(n_900), .B1(n_907), .B2(n_908), .C(n_911), .Y(n_906) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx2_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
OR2x2_ASAP7_75t_L g868 ( .A(n_869), .B(n_870), .Y(n_868) );
NOR2xp33_ASAP7_75t_L g899 ( .A(n_869), .B(n_900), .Y(n_899) );
OR2x2_ASAP7_75t_L g873 ( .A(n_870), .B(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
HB1xp67_ASAP7_75t_L g907 ( .A(n_874), .Y(n_907) );
INVxp67_ASAP7_75t_L g897 ( .A(n_875), .Y(n_897) );
NAND3xp33_ASAP7_75t_L g876 ( .A(n_877), .B(n_886), .C(n_902), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g879 ( .A1(n_880), .A2(n_881), .B1(n_883), .B2(n_884), .Y(n_879) );
INVxp67_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
AOI221xp5_ASAP7_75t_L g886 ( .A1(n_887), .A2(n_888), .B1(n_889), .B2(n_895), .C(n_899), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_890), .B(n_893), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
OR2x2_ASAP7_75t_L g896 ( .A(n_897), .B(n_898), .Y(n_896) );
INVx1_ASAP7_75t_L g915 ( .A(n_898), .Y(n_915) );
AOI211xp5_ASAP7_75t_L g902 ( .A1(n_903), .A2(n_905), .B(n_906), .C(n_917), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
HB1xp67_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
AND2x2_ASAP7_75t_L g912 ( .A(n_913), .B(n_914), .Y(n_912) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx2_ASAP7_75t_SL g921 ( .A(n_922), .Y(n_921) );
INVxp67_ASAP7_75t_SL g937 ( .A(n_924), .Y(n_937) );
INVxp33_ASAP7_75t_SL g925 ( .A(n_926), .Y(n_925) );
AOI21xp5_ASAP7_75t_L g930 ( .A1(n_931), .A2(n_937), .B(n_938), .Y(n_930) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
BUFx12f_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
CKINVDCx11_ASAP7_75t_R g934 ( .A(n_935), .Y(n_934) );
NAND3xp33_ASAP7_75t_L g938 ( .A(n_939), .B(n_940), .C(n_943), .Y(n_938) );
CKINVDCx5p33_ASAP7_75t_R g940 ( .A(n_941), .Y(n_940) );
INVx1_ASAP7_75t_SL g941 ( .A(n_942), .Y(n_941) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
NOR2xp33_ASAP7_75t_L g944 ( .A(n_945), .B(n_946), .Y(n_944) );
BUFx3_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
HB1xp67_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
CKINVDCx5p33_ASAP7_75t_R g950 ( .A(n_951), .Y(n_950) );
BUFx2_ASAP7_75t_SL g951 ( .A(n_952), .Y(n_951) );
BUFx3_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
BUFx2_ASAP7_75t_L g961 ( .A(n_953), .Y(n_961) );
AND2x4_ASAP7_75t_L g953 ( .A(n_954), .B(n_956), .Y(n_953) );
CKINVDCx20_ASAP7_75t_R g954 ( .A(n_955), .Y(n_954) );
INVx1_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
endmodule