module real_aes_2950_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_503;
wire n_287;
wire n_357;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_417;
wire n_363;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_500;
wire n_307;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_0), .B(n_214), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_1), .A2(n_209), .B(n_256), .Y(n_255) );
AOI22xp33_ASAP7_75t_SL g85 ( .A1(n_2), .A2(n_54), .B1(n_86), .B2(n_104), .Y(n_85) );
AO22x2_ASAP7_75t_L g90 ( .A1(n_3), .A2(n_55), .B1(n_91), .B2(n_92), .Y(n_90) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_4), .B(n_225), .Y(n_300) );
INVx1_ASAP7_75t_L g189 ( .A(n_5), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_6), .B(n_225), .Y(n_264) );
AO22x2_ASAP7_75t_L g94 ( .A1(n_7), .A2(n_19), .B1(n_91), .B2(n_95), .Y(n_94) );
NAND2xp33_ASAP7_75t_L g276 ( .A(n_8), .B(n_223), .Y(n_276) );
INVx2_ASAP7_75t_L g206 ( .A(n_9), .Y(n_206) );
AOI221x1_ASAP7_75t_L g208 ( .A1(n_10), .A2(n_16), .B1(n_209), .B2(n_214), .C(n_221), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_11), .B(n_214), .Y(n_272) );
AO21x2_ASAP7_75t_L g269 ( .A1(n_12), .A2(n_270), .B(n_271), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_13), .B(n_204), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_14), .B(n_225), .Y(n_284) );
AO21x1_ASAP7_75t_L g295 ( .A1(n_15), .A2(n_214), .B(n_296), .Y(n_295) );
NAND2x1_ASAP7_75t_L g233 ( .A(n_17), .B(n_225), .Y(n_233) );
NAND2x1_ASAP7_75t_L g263 ( .A(n_18), .B(n_223), .Y(n_263) );
OAI221xp5_ASAP7_75t_L g181 ( .A1(n_19), .A2(n_55), .B1(n_59), .B2(n_182), .C(n_184), .Y(n_181) );
AOI22xp33_ASAP7_75t_SL g145 ( .A1(n_20), .A2(n_60), .B1(n_146), .B2(n_148), .Y(n_145) );
OR2x2_ASAP7_75t_L g207 ( .A(n_21), .B(n_67), .Y(n_207) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_21), .A2(n_67), .B(n_206), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_22), .B(n_223), .Y(n_258) );
INVx3_ASAP7_75t_L g91 ( .A(n_23), .Y(n_91) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_24), .B(n_225), .Y(n_275) );
AOI22xp33_ASAP7_75t_SL g137 ( .A1(n_25), .A2(n_47), .B1(n_138), .B2(n_142), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_26), .B(n_223), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_26), .A2(n_80), .B1(n_167), .B2(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_26), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g109 ( .A1(n_27), .A2(n_64), .B1(n_110), .B2(n_116), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_28), .A2(n_209), .B(n_244), .Y(n_243) );
INVx1_ASAP7_75t_SL g99 ( .A(n_29), .Y(n_99) );
INVx1_ASAP7_75t_L g191 ( .A(n_30), .Y(n_191) );
AND2x2_ASAP7_75t_L g210 ( .A(n_30), .B(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g220 ( .A(n_30), .B(n_189), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_31), .B(n_214), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_32), .A2(n_80), .B1(n_166), .B2(n_167), .Y(n_79) );
INVx1_ASAP7_75t_L g166 ( .A(n_32), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_33), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_34), .B(n_223), .Y(n_245) );
AOI22xp5_ASAP7_75t_L g168 ( .A1(n_35), .A2(n_169), .B1(n_176), .B2(n_177), .Y(n_168) );
CKINVDCx16_ASAP7_75t_R g176 ( .A(n_35), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_36), .A2(n_209), .B(n_262), .Y(n_261) );
AO22x2_ASAP7_75t_L g102 ( .A1(n_37), .A2(n_59), .B1(n_91), .B2(n_103), .Y(n_102) );
AOI22xp33_ASAP7_75t_L g128 ( .A1(n_38), .A2(n_73), .B1(n_129), .B2(n_131), .Y(n_128) );
AOI22xp5_ASAP7_75t_L g153 ( .A1(n_39), .A2(n_40), .B1(n_154), .B2(n_157), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_41), .B(n_223), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_42), .A2(n_80), .B1(n_167), .B2(n_511), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_42), .Y(n_511) );
INVx1_ASAP7_75t_L g213 ( .A(n_43), .Y(n_213) );
INVx1_ASAP7_75t_L g217 ( .A(n_43), .Y(n_217) );
INVx1_ASAP7_75t_L g100 ( .A(n_44), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_45), .B(n_225), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_46), .A2(n_209), .B(n_232), .Y(n_231) );
AO21x1_ASAP7_75t_L g297 ( .A1(n_48), .A2(n_209), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g523 ( .A(n_48), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_49), .B(n_214), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_50), .A2(n_172), .B1(n_173), .B2(n_174), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_50), .Y(n_172) );
AOI22xp33_ASAP7_75t_L g159 ( .A1(n_51), .A2(n_52), .B1(n_160), .B2(n_163), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_53), .B(n_214), .Y(n_265) );
INVxp33_ASAP7_75t_L g186 ( .A(n_55), .Y(n_186) );
AND2x2_ASAP7_75t_L g248 ( .A(n_56), .B(n_205), .Y(n_248) );
INVx1_ASAP7_75t_L g211 ( .A(n_57), .Y(n_211) );
INVx1_ASAP7_75t_L g219 ( .A(n_57), .Y(n_219) );
AND2x2_ASAP7_75t_L g267 ( .A(n_58), .B(n_237), .Y(n_267) );
INVxp67_ASAP7_75t_L g185 ( .A(n_59), .Y(n_185) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_61), .Y(n_174) );
AND2x2_ASAP7_75t_L g252 ( .A(n_62), .B(n_237), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_63), .B(n_214), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_65), .Y(n_127) );
AND2x2_ASAP7_75t_L g296 ( .A(n_66), .B(n_277), .Y(n_296) );
AND2x2_ASAP7_75t_L g240 ( .A(n_68), .B(n_237), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_69), .B(n_223), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_70), .B(n_225), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g169 ( .A1(n_71), .A2(n_170), .B1(n_171), .B2(n_175), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_71), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_71), .B(n_223), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_72), .A2(n_209), .B(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_74), .B(n_225), .Y(n_257) );
BUFx2_ASAP7_75t_SL g183 ( .A(n_75), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_76), .A2(n_209), .B(n_274), .Y(n_273) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_178), .B1(n_192), .B2(n_500), .C(n_501), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_168), .Y(n_78) );
INVx1_ASAP7_75t_L g167 ( .A(n_80), .Y(n_167) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NAND2xp5_ASAP7_75t_L g82 ( .A(n_83), .B(n_135), .Y(n_82) );
NOR2xp33_ASAP7_75t_L g83 ( .A(n_84), .B(n_120), .Y(n_83) );
NAND2xp5_ASAP7_75t_L g84 ( .A(n_85), .B(n_109), .Y(n_84) );
INVx2_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
INVx3_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_96), .Y(n_88) );
AND2x4_ASAP7_75t_L g144 ( .A(n_89), .B(n_141), .Y(n_144) );
AND2x2_ASAP7_75t_L g147 ( .A(n_89), .B(n_114), .Y(n_147) );
AND2x2_ASAP7_75t_L g89 ( .A(n_90), .B(n_93), .Y(n_89) );
INVx2_ASAP7_75t_L g113 ( .A(n_90), .Y(n_113) );
AND2x2_ASAP7_75t_L g133 ( .A(n_90), .B(n_94), .Y(n_133) );
INVx1_ASAP7_75t_L g92 ( .A(n_91), .Y(n_92) );
INVx2_ASAP7_75t_L g95 ( .A(n_91), .Y(n_95) );
OAI22x1_ASAP7_75t_L g97 ( .A1(n_91), .A2(n_98), .B1(n_99), .B2(n_100), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_91), .Y(n_98) );
INVx1_ASAP7_75t_L g103 ( .A(n_91), .Y(n_103) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_93), .Y(n_108) );
INVx1_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
AND2x4_ASAP7_75t_L g112 ( .A(n_94), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g126 ( .A(n_94), .Y(n_126) );
AND2x2_ASAP7_75t_L g130 ( .A(n_96), .B(n_112), .Y(n_130) );
AND2x4_ASAP7_75t_L g162 ( .A(n_96), .B(n_125), .Y(n_162) );
AND2x2_ASAP7_75t_L g96 ( .A(n_97), .B(n_101), .Y(n_96) );
AND2x2_ASAP7_75t_L g106 ( .A(n_97), .B(n_102), .Y(n_106) );
INVx2_ASAP7_75t_L g115 ( .A(n_97), .Y(n_115) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_97), .Y(n_134) );
AND2x4_ASAP7_75t_L g141 ( .A(n_101), .B(n_115), .Y(n_141) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_L g114 ( .A(n_102), .B(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g151 ( .A(n_102), .Y(n_151) );
BUFx6f_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
AND2x4_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
AND2x4_ASAP7_75t_L g118 ( .A(n_106), .B(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g124 ( .A(n_106), .B(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AND2x4_ASAP7_75t_L g111 ( .A(n_112), .B(n_114), .Y(n_111) );
AND2x4_ASAP7_75t_L g158 ( .A(n_112), .B(n_141), .Y(n_158) );
INVxp67_ASAP7_75t_L g119 ( .A(n_113), .Y(n_119) );
AND2x4_ASAP7_75t_L g125 ( .A(n_113), .B(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g156 ( .A(n_114), .B(n_125), .Y(n_156) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx6_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI21xp33_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_127), .B(n_128), .Y(n_120) );
INVx1_ASAP7_75t_SL g121 ( .A(n_122), .Y(n_121) );
INVx4_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
INVx6_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x4_ASAP7_75t_L g140 ( .A(n_125), .B(n_141), .Y(n_140) );
BUFx5_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
BUFx12f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
AND2x4_ASAP7_75t_L g150 ( .A(n_133), .B(n_151), .Y(n_150) );
AND2x4_ASAP7_75t_L g165 ( .A(n_133), .B(n_141), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_136), .B(n_152), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_145), .Y(n_136) );
INVx2_ASAP7_75t_SL g138 ( .A(n_139), .Y(n_138) );
INVx8_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_SL g142 ( .A(n_143), .Y(n_142) );
INVx8_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx5_ASAP7_75t_SL g149 ( .A(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_153), .B(n_159), .Y(n_152) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx6_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_SL g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_169), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_171), .Y(n_175) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_179), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_180), .Y(n_179) );
AND3x1_ASAP7_75t_SL g180 ( .A(n_181), .B(n_187), .C(n_190), .Y(n_180) );
INVxp67_ASAP7_75t_L g509 ( .A(n_181), .Y(n_509) );
CKINVDCx8_ASAP7_75t_R g182 ( .A(n_183), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_185), .B(n_186), .Y(n_184) );
CKINVDCx16_ASAP7_75t_R g507 ( .A(n_187), .Y(n_507) );
OAI21xp5_ASAP7_75t_L g516 ( .A1(n_187), .A2(n_517), .B(n_520), .Y(n_516) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
OR2x2_ASAP7_75t_SL g514 ( .A(n_188), .B(n_190), .Y(n_514) );
AND2x2_ASAP7_75t_L g521 ( .A(n_188), .B(n_522), .Y(n_521) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g212 ( .A(n_189), .B(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_190), .B(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx3_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_196), .B(n_412), .Y(n_195) );
AND4x1_ASAP7_75t_L g196 ( .A(n_197), .B(n_324), .C(n_351), .D(n_386), .Y(n_196) );
AOI221xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_249), .B1(n_289), .B2(n_304), .C(n_308), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_200), .B(n_228), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_200), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
OR2x2_ASAP7_75t_L g365 ( .A(n_201), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g420 ( .A(n_201), .B(n_375), .Y(n_420) );
BUFx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g323 ( .A(n_202), .B(n_241), .Y(n_323) );
AND2x4_ASAP7_75t_L g359 ( .A(n_202), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g373 ( .A(n_202), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g290 ( .A(n_203), .Y(n_290) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_203), .Y(n_462) );
OA21x2_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_208), .B(n_227), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_204), .A2(n_254), .B(n_255), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_204), .Y(n_266) );
OA21x2_ASAP7_75t_L g336 ( .A1(n_204), .A2(n_208), .B(n_227), .Y(n_336) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_SL g205 ( .A(n_206), .B(n_207), .Y(n_205) );
AND2x4_ASAP7_75t_L g277 ( .A(n_206), .B(n_207), .Y(n_277) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_209), .Y(n_500) );
AND2x6_ASAP7_75t_L g209 ( .A(n_210), .B(n_212), .Y(n_209) );
BUFx3_ASAP7_75t_L g519 ( .A(n_210), .Y(n_519) );
AND2x6_ASAP7_75t_L g223 ( .A(n_211), .B(n_216), .Y(n_223) );
AND2x4_ASAP7_75t_L g225 ( .A(n_213), .B(n_218), .Y(n_225) );
INVx2_ASAP7_75t_L g522 ( .A(n_213), .Y(n_522) );
AND2x4_ASAP7_75t_L g214 ( .A(n_215), .B(n_220), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_216), .B(n_218), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx5_ASAP7_75t_L g226 ( .A(n_220), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_224), .B(n_226), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_226), .A2(n_233), .B(n_234), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_226), .A2(n_245), .B(n_246), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_226), .A2(n_257), .B(n_258), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_226), .A2(n_263), .B(n_264), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_226), .A2(n_275), .B(n_276), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_226), .A2(n_284), .B(n_285), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_226), .A2(n_299), .B(n_300), .Y(n_298) );
A2O1A1Ixp33_ASAP7_75t_SL g317 ( .A1(n_228), .A2(n_290), .B(n_318), .C(n_322), .Y(n_317) );
AND2x2_ASAP7_75t_L g338 ( .A(n_228), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_228), .B(n_290), .Y(n_478) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_241), .Y(n_228) );
INVx2_ASAP7_75t_L g358 ( .A(n_229), .Y(n_358) );
BUFx3_ASAP7_75t_L g374 ( .A(n_229), .Y(n_374) );
INVxp67_ASAP7_75t_L g378 ( .A(n_229), .Y(n_378) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_236), .B(n_240), .Y(n_229) );
AO21x2_ASAP7_75t_L g328 ( .A1(n_230), .A2(n_236), .B(n_240), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_235), .Y(n_230) );
AO21x2_ASAP7_75t_L g241 ( .A1(n_236), .A2(n_242), .B(n_248), .Y(n_241) );
AO21x2_ASAP7_75t_L g303 ( .A1(n_236), .A2(n_242), .B(n_248), .Y(n_303) );
INVx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx4_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx3_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
BUFx4f_ASAP7_75t_L g270 ( .A(n_239), .Y(n_270) );
INVx2_ASAP7_75t_L g357 ( .A(n_241), .Y(n_357) );
AND2x2_ASAP7_75t_L g363 ( .A(n_241), .B(n_336), .Y(n_363) );
AND2x2_ASAP7_75t_L g389 ( .A(n_241), .B(n_358), .Y(n_389) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_243), .B(n_247), .Y(n_242) );
AOI211xp5_ASAP7_75t_L g386 ( .A1(n_249), .A2(n_387), .B(n_390), .C(n_400), .Y(n_386) );
AND2x2_ASAP7_75t_SL g249 ( .A(n_250), .B(n_268), .Y(n_249) );
OAI321xp33_ASAP7_75t_L g361 ( .A1(n_250), .A2(n_309), .A3(n_362), .B1(n_364), .B2(n_365), .C(n_367), .Y(n_361) );
AND2x2_ASAP7_75t_L g482 ( .A(n_250), .B(n_457), .Y(n_482) );
INVx1_ASAP7_75t_L g485 ( .A(n_250), .Y(n_485) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_259), .Y(n_250) );
INVx5_ASAP7_75t_L g307 ( .A(n_251), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_251), .B(n_321), .Y(n_320) );
NOR2x1_ASAP7_75t_SL g352 ( .A(n_251), .B(n_353), .Y(n_352) );
BUFx2_ASAP7_75t_L g397 ( .A(n_251), .Y(n_397) );
AND2x2_ASAP7_75t_L g499 ( .A(n_251), .B(n_269), .Y(n_499) );
OR2x6_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
AND2x2_ASAP7_75t_L g306 ( .A(n_259), .B(n_307), .Y(n_306) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_259), .Y(n_316) );
INVx4_ASAP7_75t_L g321 ( .A(n_259), .Y(n_321) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_266), .B(n_267), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_265), .Y(n_260) );
INVx1_ASAP7_75t_L g364 ( .A(n_268), .Y(n_364) );
A2O1A1Ixp33_ASAP7_75t_R g467 ( .A1(n_268), .A2(n_306), .B(n_338), .C(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g487 ( .A(n_268), .B(n_312), .Y(n_487) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_278), .Y(n_268) );
INVx1_ASAP7_75t_L g305 ( .A(n_269), .Y(n_305) );
INVx2_ASAP7_75t_L g311 ( .A(n_269), .Y(n_311) );
OR2x2_ASAP7_75t_L g330 ( .A(n_269), .B(n_321), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_269), .B(n_353), .Y(n_399) );
BUFx3_ASAP7_75t_L g406 ( .A(n_269), .Y(n_406) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_273), .B(n_277), .Y(n_271) );
INVx1_ASAP7_75t_SL g280 ( .A(n_277), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_277), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g369 ( .A(n_278), .Y(n_369) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_278), .Y(n_382) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g315 ( .A(n_279), .Y(n_315) );
INVx1_ASAP7_75t_L g424 ( .A(n_279), .Y(n_424) );
AO21x2_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_281), .B(n_287), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_280), .B(n_288), .Y(n_287) );
AO21x2_ASAP7_75t_L g353 ( .A1(n_280), .A2(n_281), .B(n_287), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_286), .Y(n_281) );
AND2x2_ASAP7_75t_L g325 ( .A(n_289), .B(n_326), .Y(n_325) );
OAI31xp33_ASAP7_75t_L g476 ( .A1(n_289), .A2(n_477), .A3(n_479), .B(n_482), .Y(n_476) );
INVx1_ASAP7_75t_SL g494 ( .A(n_289), .Y(n_494) );
AND2x4_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
AOI21xp33_ASAP7_75t_L g308 ( .A1(n_290), .A2(n_309), .B(n_317), .Y(n_308) );
NAND2x1_ASAP7_75t_L g388 ( .A(n_290), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_SL g417 ( .A(n_290), .Y(n_417) );
INVx2_ASAP7_75t_L g366 ( .A(n_291), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_291), .B(n_349), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_291), .B(n_348), .Y(n_458) );
NOR2xp33_ASAP7_75t_SL g466 ( .A(n_291), .B(n_417), .Y(n_466) );
AND2x4_ASAP7_75t_L g291 ( .A(n_292), .B(n_303), .Y(n_291) );
AND2x2_ASAP7_75t_SL g335 ( .A(n_292), .B(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g346 ( .A(n_292), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g375 ( .A(n_292), .B(n_357), .Y(n_375) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
BUFx2_ASAP7_75t_L g339 ( .A(n_293), .Y(n_339) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g360 ( .A(n_294), .Y(n_360) );
OAI21x1_ASAP7_75t_SL g294 ( .A1(n_295), .A2(n_297), .B(n_301), .Y(n_294) );
INVx1_ASAP7_75t_L g302 ( .A(n_296), .Y(n_302) );
INVx2_ASAP7_75t_L g347 ( .A(n_303), .Y(n_347) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_303), .Y(n_407) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx1_ASAP7_75t_L g343 ( .A(n_305), .Y(n_343) );
AND2x2_ASAP7_75t_L g422 ( .A(n_305), .B(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g333 ( .A(n_306), .B(n_327), .Y(n_333) );
INVx2_ASAP7_75t_SL g381 ( .A(n_306), .Y(n_381) );
INVx4_ASAP7_75t_L g312 ( .A(n_307), .Y(n_312) );
AND2x2_ASAP7_75t_L g410 ( .A(n_307), .B(n_353), .Y(n_410) );
AND2x2_ASAP7_75t_SL g428 ( .A(n_307), .B(n_423), .Y(n_428) );
NAND2x1p5_ASAP7_75t_L g445 ( .A(n_307), .B(n_321), .Y(n_445) );
INVx1_ASAP7_75t_L g451 ( .A(n_309), .Y(n_451) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_313), .Y(n_309) );
INVx1_ASAP7_75t_L g370 ( .A(n_310), .Y(n_370) );
OR2x2_ASAP7_75t_L g383 ( .A(n_310), .B(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
OR2x2_ASAP7_75t_L g435 ( .A(n_311), .B(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g465 ( .A(n_311), .B(n_353), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_312), .B(n_315), .Y(n_341) );
AND2x2_ASAP7_75t_L g433 ( .A(n_312), .B(n_423), .Y(n_433) );
AND2x4_ASAP7_75t_L g495 ( .A(n_312), .B(n_374), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
INVx2_ASAP7_75t_L g319 ( .A(n_314), .Y(n_319) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NOR2xp67_ASAP7_75t_SL g318 ( .A(n_319), .B(n_320), .Y(n_318) );
OAI322xp33_ASAP7_75t_SL g331 ( .A1(n_319), .A2(n_332), .A3(n_334), .B1(n_337), .B2(n_340), .C1(n_342), .C2(n_344), .Y(n_331) );
INVx1_ASAP7_75t_L g489 ( .A(n_319), .Y(n_489) );
OR2x2_ASAP7_75t_L g342 ( .A(n_320), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g368 ( .A(n_321), .B(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_321), .B(n_369), .Y(n_384) );
INVx2_ASAP7_75t_L g411 ( .A(n_321), .Y(n_411) );
AND2x4_ASAP7_75t_L g423 ( .A(n_321), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_SL g426 ( .A(n_323), .B(n_339), .Y(n_426) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_329), .B(n_331), .Y(n_324) );
AND2x2_ASAP7_75t_L g392 ( .A(n_326), .B(n_359), .Y(n_392) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_327), .B(n_481), .Y(n_480) );
BUFx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g350 ( .A(n_328), .Y(n_350) );
AND2x4_ASAP7_75t_SL g432 ( .A(n_328), .B(n_347), .Y(n_432) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g340 ( .A(n_330), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_333), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g468 ( .A(n_335), .B(n_432), .Y(n_468) );
NOR4xp25_ASAP7_75t_L g472 ( .A(n_335), .B(n_349), .C(n_389), .D(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g349 ( .A(n_336), .B(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g385 ( .A(n_336), .B(n_360), .Y(n_385) );
AND2x4_ASAP7_75t_L g449 ( .A(n_336), .B(n_360), .Y(n_449) );
INVx1_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_339), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
OR2x2_ASAP7_75t_L g438 ( .A(n_346), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g492 ( .A(n_346), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_347), .B(n_359), .Y(n_393) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
AOI211xp5_ASAP7_75t_SL g351 ( .A1(n_352), .A2(n_354), .B(n_361), .C(n_376), .Y(n_351) );
INVx1_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_359), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_357), .B(n_360), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_358), .B(n_363), .Y(n_362) );
BUFx2_ASAP7_75t_L g440 ( .A(n_358), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_359), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g455 ( .A(n_359), .Y(n_455) );
OAI21xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_370), .B(n_371), .Y(n_367) );
AND2x4_ASAP7_75t_L g404 ( .A(n_368), .B(n_405), .Y(n_404) );
AND2x4_ASAP7_75t_L g498 ( .A(n_368), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_375), .Y(n_372) );
INVx1_ASAP7_75t_SL g402 ( .A(n_374), .Y(n_402) );
AND2x2_ASAP7_75t_L g461 ( .A(n_375), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g475 ( .A(n_375), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_SL g376 ( .A1(n_377), .A2(n_379), .B(n_383), .C(n_385), .Y(n_376) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_377), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g453 ( .A(n_378), .B(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g474 ( .A(n_378), .B(n_475), .Y(n_474) );
INVxp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
OR2x2_ASAP7_75t_L g463 ( .A(n_381), .B(n_405), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_384), .A2(n_391), .B1(n_393), .B2(n_394), .Y(n_390) );
INVx1_ASAP7_75t_SL g481 ( .A(n_385), .Y(n_481) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVxp67_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_398), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_396), .B(n_405), .Y(n_447) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVxp67_ASAP7_75t_SL g457 ( .A(n_399), .Y(n_457) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_403), .B1(n_407), .B2(n_408), .Y(n_400) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AOI21xp5_ASAP7_75t_SL g414 ( .A1(n_405), .A2(n_415), .B(n_418), .Y(n_414) );
AND2x2_ASAP7_75t_L g443 ( .A(n_405), .B(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND3x2_ASAP7_75t_L g409 ( .A(n_406), .B(n_410), .C(n_411), .Y(n_409) );
AND2x2_ASAP7_75t_L g471 ( .A(n_406), .B(n_428), .Y(n_471) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g456 ( .A(n_411), .B(n_457), .Y(n_456) );
NOR2xp67_ASAP7_75t_L g412 ( .A(n_413), .B(n_469), .Y(n_412) );
NAND4xp25_ASAP7_75t_L g413 ( .A(n_414), .B(n_429), .C(n_450), .D(n_467), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_421), .B1(n_425), .B2(n_427), .Y(n_418) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_421), .A2(n_435), .B1(n_455), .B2(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g436 ( .A(n_423), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_425), .A2(n_448), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx3_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
AOI221xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_433), .B1(n_434), .B2(n_437), .C(n_441), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_446), .B1(n_447), .B2(n_448), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_444), .B(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_444), .B(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AOI221xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_452), .B1(n_456), .B2(n_458), .C(n_459), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_453), .B(n_455), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_463), .B1(n_464), .B2(n_466), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OAI211xp5_ASAP7_75t_SL g484 ( .A1(n_465), .A2(n_485), .B(n_486), .C(n_488), .Y(n_484) );
OAI211xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_472), .B(n_476), .C(n_483), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_SL g479 ( .A(n_480), .Y(n_479) );
AOI221xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_490), .B1(n_493), .B2(n_495), .C(n_496), .Y(n_483) );
INVx1_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
OAI222xp33_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_504), .B1(n_510), .B2(n_512), .C1(n_515), .C2(n_523), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_505), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_506), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
CKINVDCx16_ASAP7_75t_R g515 ( .A(n_516), .Y(n_515) );
INVxp67_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
endmodule