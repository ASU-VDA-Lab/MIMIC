module fake_jpeg_25721_n_146 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_146);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_9),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_7),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_23),
.Y(n_35)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

AOI21xp33_ASAP7_75t_L g23 ( 
.A1(n_13),
.A2(n_7),
.B(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_13),
.B(n_19),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_21),
.A2(n_18),
.B1(n_16),
.B2(n_15),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_29),
.A2(n_32),
.B1(n_26),
.B2(n_12),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_21),
.A2(n_18),
.B1(n_16),
.B2(n_15),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_33),
.A2(n_34),
.B1(n_17),
.B2(n_10),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_20),
.A2(n_19),
.B1(n_17),
.B2(n_10),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_36),
.A2(n_37),
.B1(n_31),
.B2(n_28),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_17),
.B1(n_10),
.B2(n_24),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_44),
.Y(n_48)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_45),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_31),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_11),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_35),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_11),
.B1(n_12),
.B2(n_24),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_47),
.A2(n_31),
.B1(n_28),
.B2(n_27),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_54),
.Y(n_62)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_41),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_33),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_59),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_11),
.B(n_12),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_58),
.B1(n_47),
.B2(n_40),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_46),
.B(n_25),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_53),
.B1(n_39),
.B2(n_42),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_64),
.B1(n_65),
.B2(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_51),
.B(n_44),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_66),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_44),
.B1(n_36),
.B2(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_55),
.B(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_11),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_69),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_70),
.A2(n_50),
.B(n_45),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_68),
.Y(n_85)
);

AOI322xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_54),
.A3(n_58),
.B1(n_59),
.B2(n_50),
.C1(n_52),
.C2(n_25),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_30),
.Y(n_93)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_59),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_80),
.Y(n_83)
);

OA21x2_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_59),
.B(n_31),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_68),
.B(n_30),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_22),
.C(n_25),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_43),
.B1(n_28),
.B2(n_31),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_81),
.A2(n_67),
.B1(n_43),
.B2(n_65),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_73),
.A2(n_60),
.B1(n_70),
.B2(n_66),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_82),
.A2(n_89),
.B1(n_90),
.B2(n_28),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_84),
.A2(n_71),
.B1(n_81),
.B2(n_75),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_79),
.A2(n_0),
.B(n_1),
.Y(n_89)
);

NAND2xp33_ASAP7_75t_R g90 ( 
.A(n_79),
.B(n_73),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_24),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_77),
.Y(n_95)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_72),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_78),
.Y(n_94)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_102),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_97),
.A2(n_104),
.B1(n_30),
.B2(n_22),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_80),
.C(n_79),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_101),
.C(n_85),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_75),
.C(n_76),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_76),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_89),
.Y(n_109)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_82),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_108),
.C(n_109),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_84),
.C(n_86),
.Y(n_108)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_104),
.A2(n_9),
.B(n_1),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_114),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_99),
.A2(n_9),
.B1(n_30),
.B2(n_2),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_98),
.A2(n_0),
.B(n_1),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_115),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_101),
.B(n_0),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_108),
.A2(n_96),
.B1(n_106),
.B2(n_95),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_22),
.Y(n_127)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_111),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_118),
.A2(n_107),
.B(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_126),
.A2(n_127),
.B(n_129),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_0),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_130),
.C(n_121),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_123),
.A2(n_2),
.B(n_3),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_2),
.C(n_3),
.Y(n_130)
);

OAI321xp33_ASAP7_75t_L g131 ( 
.A1(n_126),
.A2(n_117),
.A3(n_120),
.B1(n_123),
.B2(n_118),
.C(n_121),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_132),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_133),
.B(n_124),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_117),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_139),
.C(n_5),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_122),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_138),
.Y(n_140)
);

AOI21x1_ASAP7_75t_L g141 ( 
.A1(n_137),
.A2(n_124),
.B(n_3),
.Y(n_141)
);

AOI31xp33_ASAP7_75t_L g144 ( 
.A1(n_141),
.A2(n_4),
.A3(n_5),
.B(n_140),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_2),
.C(n_4),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_143),
.A2(n_144),
.B(n_4),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_5),
.Y(n_146)
);


endmodule