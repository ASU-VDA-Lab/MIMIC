module fake_jpeg_20398_n_292 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_292);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_292;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_247;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_273;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_9),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_40),
.Y(n_47)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_0),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_21),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_25),
.B1(n_19),
.B2(n_23),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_44),
.A2(n_54),
.B1(n_38),
.B2(n_39),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_25),
.B1(n_41),
.B2(n_35),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_45),
.A2(n_58),
.B1(n_39),
.B2(n_38),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_27),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_49),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_21),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_59),
.Y(n_76)
);

AO22x1_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_42),
.B1(n_41),
.B2(n_35),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_25),
.B1(n_30),
.B2(n_22),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_41),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_30),
.B1(n_26),
.B2(n_32),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_34),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_29),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_60),
.B(n_26),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_63),
.B(n_68),
.Y(n_102)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_64),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_SL g110 ( 
.A(n_65),
.B(n_79),
.C(n_81),
.Y(n_110)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVxp67_ASAP7_75t_SL g99 ( 
.A(n_66),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_43),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_57),
.A2(n_41),
.B1(n_35),
.B2(n_40),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_69),
.A2(n_72),
.B1(n_79),
.B2(n_82),
.Y(n_121)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g115 ( 
.A(n_70),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_74),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_54),
.A2(n_40),
.B(n_33),
.C(n_31),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_59),
.B(n_23),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_73),
.B(n_88),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_22),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

OAI32xp33_ASAP7_75t_L g77 ( 
.A1(n_49),
.A2(n_46),
.A3(n_44),
.B1(n_47),
.B2(n_60),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_95),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_28),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_83),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_39),
.B1(n_38),
.B2(n_40),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_80),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_39),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_45),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_52),
.A2(n_39),
.B1(n_38),
.B2(n_28),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_85),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_48),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_54),
.A2(n_39),
.B1(n_38),
.B2(n_33),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_55),
.A2(n_38),
.B1(n_33),
.B2(n_31),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_55),
.A2(n_17),
.B1(n_36),
.B2(n_21),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_58),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_92),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_55),
.B(n_26),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_48),
.B(n_21),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_96),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_22),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_77),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_62),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_106),
.B(n_122),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_61),
.B1(n_51),
.B2(n_31),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_98),
.B1(n_111),
.B2(n_121),
.Y(n_130)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_110),
.A2(n_74),
.B(n_72),
.Y(n_127)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_91),
.A2(n_24),
.B1(n_32),
.B2(n_51),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_112),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_81),
.A2(n_24),
.B(n_21),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_113),
.A2(n_65),
.B(n_67),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

INVxp67_ASAP7_75t_SL g132 ( 
.A(n_116),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_21),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_120),
.Y(n_138)
);

OAI32xp33_ASAP7_75t_L g120 ( 
.A1(n_67),
.A2(n_24),
.A3(n_18),
.B1(n_12),
.B2(n_16),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_69),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_76),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_125),
.B(n_129),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_127),
.A2(n_133),
.B(n_136),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_128),
.B(n_120),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_76),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_130),
.A2(n_122),
.B1(n_110),
.B2(n_113),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_71),
.B(n_114),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_97),
.B(n_68),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_146),
.Y(n_180)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_65),
.B1(n_90),
.B2(n_66),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_141),
.A2(n_143),
.B1(n_98),
.B2(n_121),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_64),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_112),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_75),
.B1(n_70),
.B2(n_96),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_97),
.B(n_93),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_99),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_148),
.B(n_149),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_102),
.B(n_114),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_150),
.Y(n_168)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_151),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_100),
.B(n_93),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_152),
.B(n_154),
.Y(n_179)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_153),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_109),
.B(n_61),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_101),
.B(n_109),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_155),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_156),
.A2(n_51),
.B1(n_84),
.B2(n_83),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_158),
.A2(n_153),
.B1(n_151),
.B2(n_150),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_102),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_161),
.B(n_167),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_118),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_163),
.B(n_176),
.Y(n_198)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_173),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_141),
.B1(n_130),
.B2(n_145),
.Y(n_170)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_181),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_178),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_135),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_117),
.C(n_107),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_131),
.C(n_138),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_126),
.B(n_117),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_115),
.Y(n_191)
);

AO22x1_ASAP7_75t_L g178 ( 
.A1(n_138),
.A2(n_106),
.B1(n_115),
.B2(n_123),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_115),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_131),
.A2(n_134),
.B(n_127),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_148),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_175),
.C(n_176),
.Y(n_215)
);

AOI322xp5_ASAP7_75t_L g187 ( 
.A1(n_159),
.A2(n_139),
.A3(n_126),
.B1(n_137),
.B2(n_146),
.C1(n_140),
.C2(n_135),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_202),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_188),
.A2(n_183),
.B(n_155),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_194),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_193),
.A2(n_201),
.B1(n_204),
.B2(n_0),
.Y(n_228)
);

INVxp67_ASAP7_75t_SL g194 ( 
.A(n_169),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_172),
.Y(n_195)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

AOI221xp5_ASAP7_75t_L g197 ( 
.A1(n_159),
.A2(n_147),
.B1(n_18),
.B2(n_123),
.C(n_13),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_179),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_199),
.A2(n_200),
.B1(n_206),
.B2(n_157),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_156),
.A2(n_93),
.B1(n_17),
.B2(n_36),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_158),
.A2(n_10),
.B1(n_16),
.B2(n_15),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_157),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_205),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_167),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_162),
.B(n_8),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_170),
.A2(n_17),
.B1(n_36),
.B2(n_18),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_163),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_212),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_211),
.A2(n_209),
.B1(n_195),
.B2(n_207),
.Y(n_234)
);

XNOR2x1_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_171),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_214),
.A2(n_205),
.B(n_13),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_229),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_181),
.C(n_178),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_218),
.C(n_222),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_207),
.A2(n_174),
.B1(n_165),
.B2(n_164),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_217),
.A2(n_221),
.B1(n_203),
.B2(n_193),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_178),
.C(n_180),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_219),
.B(n_228),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_188),
.A2(n_170),
.B(n_180),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_220),
.A2(n_185),
.B(n_221),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_189),
.A2(n_170),
.B1(n_166),
.B2(n_168),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_182),
.C(n_168),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_201),
.A2(n_17),
.B1(n_7),
.B2(n_9),
.Y(n_224)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_224),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_185),
.B(n_13),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_230),
.A2(n_244),
.B(n_0),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_222),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_237),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_225),
.A2(n_189),
.B1(n_200),
.B2(n_206),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_232),
.A2(n_241),
.B1(n_246),
.B2(n_1),
.Y(n_256)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_234),
.B(n_2),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_213),
.A2(n_192),
.B(n_202),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_236),
.A2(n_0),
.B(n_1),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_192),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_220),
.A2(n_204),
.B1(n_199),
.B2(n_196),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_190),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_212),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_12),
.C(n_11),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_219),
.C(n_229),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_211),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_214),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_249),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_251),
.B(n_242),
.Y(n_268)
);

NAND4xp25_ASAP7_75t_SL g252 ( 
.A(n_236),
.B(n_217),
.C(n_223),
.D(n_227),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_256),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_226),
.C(n_1),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_258),
.C(n_259),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_254),
.A2(n_244),
.B(n_255),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_255),
.A2(n_257),
.B1(n_3),
.B2(n_5),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_2),
.C(n_3),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_2),
.C(n_3),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

A2O1A1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_250),
.A2(n_230),
.B(n_233),
.C(n_241),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_261),
.A2(n_263),
.B(n_242),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_232),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_265),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_235),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_245),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_248),
.A2(n_238),
.B(n_243),
.Y(n_266)
);

OAI21x1_ASAP7_75t_SL g276 ( 
.A1(n_266),
.A2(n_269),
.B(n_267),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_239),
.C(n_249),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_270),
.B(n_251),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_273),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_259),
.B(n_247),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_275),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_247),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_276),
.A2(n_278),
.B1(n_267),
.B2(n_260),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_280),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_277),
.A2(n_269),
.B(n_261),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_239),
.C(n_5),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_284),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_5),
.Y(n_284)
);

INVxp33_ASAP7_75t_L g287 ( 
.A(n_284),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_281),
.A2(n_5),
.B(n_6),
.Y(n_285)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_285),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_288),
.A2(n_6),
.B1(n_282),
.B2(n_287),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_289),
.A2(n_6),
.B(n_286),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_290),
.Y(n_292)
);


endmodule