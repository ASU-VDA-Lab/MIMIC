module fake_jpeg_2731_n_584 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_584);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_584;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_548;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_17),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_18),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_4),
.B(n_0),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_54),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_22),
.B(n_29),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_55),
.B(n_71),
.Y(n_114)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_34),
.Y(n_56)
);

CKINVDCx12_ASAP7_75t_R g150 ( 
.A(n_56),
.Y(n_150)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_58),
.Y(n_141)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_60),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_61),
.Y(n_149)
);

NAND2xp67_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_0),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_62),
.B(n_48),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_64),
.Y(n_156)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_66),
.Y(n_148)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_67),
.Y(n_146)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_17),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_74),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_75),
.Y(n_154)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_76),
.Y(n_171)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_77),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_79),
.Y(n_145)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_80),
.Y(n_170)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_81),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_83),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_47),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_88),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_22),
.B(n_16),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_94),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_90),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_91),
.Y(n_159)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

BUFx24_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_93),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_29),
.B(n_16),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_49),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_104),
.Y(n_112)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_97),
.Y(n_162)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_32),
.B(n_15),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_103),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_35),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_100),
.Y(n_139)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_40),
.Y(n_102)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_32),
.B(n_0),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_25),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_35),
.Y(n_105)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_21),
.B(n_0),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_107),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_36),
.B(n_1),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_44),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_27),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_27),
.C(n_46),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_110),
.B(n_113),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_27),
.C(n_46),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_115),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_63),
.A2(n_72),
.B1(n_74),
.B2(n_73),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_120),
.A2(n_142),
.B1(n_155),
.B2(n_83),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_85),
.A2(n_36),
.B(n_24),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_125),
.A2(n_112),
.B(n_48),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_57),
.B(n_24),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_126),
.B(n_168),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_88),
.A2(n_36),
.B1(n_50),
.B2(n_44),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_140),
.A2(n_93),
.B1(n_92),
.B2(n_54),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_97),
.A2(n_53),
.B1(n_50),
.B2(n_44),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_144),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_56),
.B(n_21),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_152),
.B(n_166),
.Y(n_203)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_67),
.A2(n_53),
.B1(n_50),
.B2(n_48),
.Y(n_153)
);

O2A1O1Ixp33_ASAP7_75t_SL g195 ( 
.A1(n_153),
.A2(n_167),
.B(n_142),
.C(n_140),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_100),
.A2(n_53),
.B1(n_38),
.B2(n_23),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_76),
.Y(n_166)
);

OA22x2_ASAP7_75t_L g167 ( 
.A1(n_102),
.A2(n_62),
.B1(n_79),
.B2(n_105),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_78),
.B(n_42),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_58),
.B(n_42),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_169),
.B(n_60),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_82),
.B(n_39),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_L g186 ( 
.A1(n_173),
.A2(n_48),
.B(n_37),
.Y(n_186)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_174),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_175),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_115),
.B(n_39),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_176),
.B(n_185),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_177),
.A2(n_189),
.B1(n_193),
.B2(n_201),
.Y(n_290)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_178),
.Y(n_237)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_179),
.Y(n_255)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_181),
.Y(n_254)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_182),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_133),
.A2(n_38),
.B(n_31),
.C(n_23),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_183),
.A2(n_185),
.B(n_176),
.C(n_187),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_141),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_184),
.B(n_190),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_132),
.B(n_26),
.Y(n_185)
);

AOI21xp33_ASAP7_75t_L g289 ( 
.A1(n_186),
.A2(n_9),
.B(n_10),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_117),
.B(n_26),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_187),
.B(n_196),
.Y(n_249)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_188),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_162),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_191),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_148),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_192),
.B(n_213),
.Y(n_282)
);

INVx11_ASAP7_75t_L g193 ( 
.A(n_122),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_194),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_195),
.A2(n_222),
.B1(n_165),
.B2(n_157),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_119),
.B(n_30),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_124),
.B(n_30),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_197),
.B(n_224),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_198),
.A2(n_116),
.B(n_122),
.Y(n_269)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_199),
.Y(n_286)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_159),
.Y(n_200)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_200),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_137),
.A2(n_31),
.B1(n_104),
.B2(n_61),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_162),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_202),
.B(n_208),
.Y(n_245)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_204),
.Y(n_240)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_127),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_205),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_167),
.A2(n_104),
.B1(n_61),
.B2(n_75),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_206),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_154),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_207),
.Y(n_263)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_127),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_209),
.Y(n_284)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_172),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_210),
.B(n_215),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_167),
.A2(n_108),
.B1(n_91),
.B2(n_90),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_211),
.A2(n_229),
.B1(n_233),
.B2(n_165),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_131),
.B(n_114),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_212),
.B(n_221),
.Y(n_258)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_161),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_153),
.A2(n_87),
.B1(n_84),
.B2(n_37),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_216),
.A2(n_136),
.B1(n_111),
.B2(n_157),
.Y(n_244)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_135),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_217),
.B(n_218),
.Y(n_260)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_135),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_156),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_219),
.B(n_220),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_150),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_123),
.B(n_64),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_153),
.A2(n_75),
.B1(n_86),
.B2(n_37),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_149),
.A2(n_148),
.B1(n_143),
.B2(n_130),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_223),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_109),
.B(n_2),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_164),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_225),
.B(n_228),
.Y(n_267)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_111),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_226),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_129),
.B(n_2),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_227),
.B(n_234),
.Y(n_283)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_156),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_118),
.A2(n_43),
.B1(n_66),
.B2(n_5),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_130),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_230),
.B(n_232),
.Y(n_279)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_128),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_139),
.A2(n_43),
.B1(n_3),
.B2(n_5),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_138),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_134),
.B(n_2),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_236),
.B(n_7),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_180),
.B(n_170),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_238),
.B(n_239),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_180),
.B(n_149),
.C(n_143),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g328 ( 
.A1(n_244),
.A2(n_287),
.B1(n_193),
.B2(n_179),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_247),
.A2(n_253),
.B1(n_222),
.B2(n_229),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_248),
.B(n_281),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_203),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_251),
.Y(n_329)
);

A2O1A1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_214),
.A2(n_116),
.B(n_5),
.C(n_6),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_259),
.A2(n_269),
.B(n_289),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_180),
.B(n_171),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_261),
.B(n_268),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_211),
.A2(n_171),
.B1(n_147),
.B2(n_121),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_264),
.A2(n_270),
.B1(n_280),
.B2(n_184),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_231),
.B(n_138),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_177),
.A2(n_147),
.B1(n_121),
.B2(n_122),
.Y(n_270)
);

NOR2x1_ASAP7_75t_L g273 ( 
.A(n_196),
.B(n_116),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_273),
.B(n_291),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_235),
.B(n_2),
.C(n_6),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_274),
.B(n_218),
.Y(n_310)
);

AND2x2_ASAP7_75t_SL g276 ( 
.A(n_178),
.B(n_6),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_276),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_235),
.B(n_15),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_188),
.Y(n_303)
);

AOI32xp33_ASAP7_75t_L g278 ( 
.A1(n_198),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_233),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_195),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_280)
);

INVx13_ASAP7_75t_L g285 ( 
.A(n_220),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_285),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_197),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_207),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_288),
.B(n_228),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_293),
.A2(n_302),
.B1(n_305),
.B2(n_308),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_294),
.B(n_317),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_269),
.A2(n_195),
.B(n_192),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_295),
.A2(n_306),
.B(n_325),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_251),
.B(n_258),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_296),
.B(n_300),
.Y(n_345)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_241),
.Y(n_298)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_298),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_258),
.B(n_204),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_247),
.A2(n_224),
.B1(n_236),
.B2(n_234),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_303),
.B(n_313),
.Y(n_349)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_241),
.Y(n_304)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_304),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_259),
.A2(n_230),
.B(n_183),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_255),
.Y(n_307)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_307),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_261),
.A2(n_202),
.B1(n_190),
.B2(n_225),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_310),
.B(n_332),
.Y(n_360)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_256),
.Y(n_311)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_311),
.Y(n_380)
);

INVx2_ASAP7_75t_R g312 ( 
.A(n_259),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_312),
.B(n_342),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_275),
.B(n_200),
.Y(n_313)
);

AO22x1_ASAP7_75t_SL g315 ( 
.A1(n_253),
.A2(n_194),
.B1(n_215),
.B2(n_213),
.Y(n_315)
);

OA21x2_ASAP7_75t_L g358 ( 
.A1(n_315),
.A2(n_237),
.B(n_262),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_238),
.A2(n_209),
.B1(n_205),
.B2(n_232),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_316),
.A2(n_237),
.B1(n_262),
.B2(n_279),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_245),
.B(n_182),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_270),
.A2(n_264),
.B1(n_275),
.B2(n_249),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_318),
.A2(n_337),
.B1(n_339),
.B2(n_274),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_245),
.B(n_191),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_319),
.B(n_322),
.Y(n_362)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_272),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_320),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_281),
.B(n_174),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_321),
.B(n_326),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_268),
.B(n_283),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_255),
.Y(n_323)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_323),
.Y(n_381)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_324),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_273),
.A2(n_217),
.B(n_207),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_283),
.B(n_210),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_249),
.B(n_199),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_327),
.B(n_331),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_328),
.B(n_333),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_276),
.B(n_219),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_248),
.B(n_181),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_265),
.B(n_226),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_276),
.B(n_12),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_335),
.B(n_336),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_276),
.B(n_12),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_290),
.A2(n_13),
.B1(n_14),
.B2(n_257),
.Y(n_337)
);

BUFx12_ASAP7_75t_L g338 ( 
.A(n_285),
.Y(n_338)
);

INVx13_ASAP7_75t_L g368 ( 
.A(n_338),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_246),
.A2(n_13),
.B1(n_248),
.B2(n_273),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_277),
.B(n_246),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_340),
.B(n_282),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_256),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_341),
.B(n_343),
.Y(n_369)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_272),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_265),
.B(n_240),
.Y(n_343)
);

NAND2xp33_ASAP7_75t_SL g344 ( 
.A(n_325),
.B(n_239),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_344),
.A2(n_374),
.B(n_338),
.Y(n_425)
);

XOR2x2_ASAP7_75t_L g350 ( 
.A(n_330),
.B(n_278),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_350),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_329),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_351),
.B(n_355),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_354),
.A2(n_373),
.B1(n_327),
.B2(n_341),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_329),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_330),
.B(n_279),
.C(n_267),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_356),
.B(n_370),
.C(n_379),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_358),
.B(n_372),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_308),
.Y(n_364)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_364),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_315),
.B(n_267),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_365),
.Y(n_411)
);

CKINVDCx12_ASAP7_75t_R g367 ( 
.A(n_338),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_367),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_310),
.B(n_292),
.C(n_260),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_371),
.A2(n_375),
.B1(n_384),
.B2(n_305),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_324),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_293),
.A2(n_291),
.B1(n_250),
.B2(n_260),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_332),
.A2(n_285),
.B(n_288),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_302),
.A2(n_250),
.B1(n_254),
.B2(n_292),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_298),
.B(n_243),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_376),
.B(n_382),
.Y(n_424)
);

A2O1A1Ixp33_ASAP7_75t_L g378 ( 
.A1(n_309),
.A2(n_282),
.B(n_252),
.C(n_284),
.Y(n_378)
);

OAI21xp33_ASAP7_75t_L g413 ( 
.A1(n_378),
.A2(n_344),
.B(n_353),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_313),
.B(n_243),
.C(n_282),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_304),
.B(n_242),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_383),
.B(n_299),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_318),
.A2(n_254),
.B1(n_255),
.B2(n_242),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_339),
.B(n_271),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_385),
.B(n_271),
.Y(n_426)
);

AND2x6_ASAP7_75t_L g387 ( 
.A(n_309),
.B(n_263),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_387),
.B(n_301),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_389),
.B(n_375),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_390),
.B(n_359),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_363),
.A2(n_295),
.B(n_297),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_391),
.A2(n_409),
.B(n_414),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_357),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_392),
.B(n_415),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_361),
.A2(n_364),
.B1(n_371),
.B2(n_347),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_394),
.A2(n_406),
.B1(n_420),
.B2(n_427),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_395),
.A2(n_401),
.B1(n_423),
.B2(n_365),
.Y(n_446)
);

NAND3xp33_ASAP7_75t_L g397 ( 
.A(n_345),
.B(n_340),
.C(n_326),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_397),
.B(n_359),
.Y(n_454)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_386),
.Y(n_399)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_399),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_360),
.B(n_299),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_400),
.B(n_379),
.C(n_378),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_361),
.A2(n_312),
.B1(n_297),
.B2(n_306),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_383),
.B(n_311),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_402),
.B(n_403),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_356),
.B(n_316),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_405),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_363),
.A2(n_301),
.B1(n_334),
.B2(n_331),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_386),
.Y(n_407)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_407),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_370),
.B(n_303),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_408),
.B(n_360),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_374),
.A2(n_301),
.B(n_334),
.Y(n_409)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_357),
.Y(n_412)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_412),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_413),
.B(n_426),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_373),
.A2(n_337),
.B1(n_312),
.B2(n_314),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_380),
.Y(n_415)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_380),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_417),
.B(n_418),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_345),
.B(n_321),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_352),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_419),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_346),
.A2(n_315),
.B1(n_336),
.B2(n_335),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_349),
.B(n_342),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_421),
.B(n_384),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_351),
.A2(n_314),
.B(n_338),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_422),
.A2(n_425),
.B(n_355),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_365),
.A2(n_315),
.B1(n_320),
.B2(n_307),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_346),
.A2(n_307),
.B1(n_323),
.B2(n_286),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_430),
.B(n_433),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_396),
.B(n_350),
.C(n_369),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_435),
.B(n_436),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_396),
.B(n_350),
.C(n_349),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_404),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_437),
.B(n_443),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_403),
.B(n_353),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_439),
.B(n_440),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_408),
.B(n_402),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_398),
.B(n_348),
.C(n_377),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_442),
.B(n_444),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_404),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_446),
.A2(n_416),
.B1(n_411),
.B2(n_420),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_400),
.B(n_362),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_447),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_448),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_390),
.B(n_377),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_449),
.B(n_450),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_398),
.B(n_394),
.C(n_406),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_395),
.B(n_348),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_451),
.B(n_457),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_452),
.A2(n_423),
.B1(n_416),
.B2(n_414),
.Y(n_480)
);

NAND3xp33_ASAP7_75t_L g484 ( 
.A(n_454),
.B(n_456),
.C(n_460),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_424),
.B(n_372),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_409),
.B(n_346),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_393),
.B(n_388),
.C(n_354),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_458),
.B(n_416),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_404),
.B(n_388),
.Y(n_460)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_461),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_434),
.A2(n_428),
.B1(n_401),
.B2(n_452),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_462),
.A2(n_480),
.B1(n_457),
.B2(n_458),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_431),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_463),
.B(n_467),
.Y(n_491)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_432),
.Y(n_465)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_465),
.Y(n_493)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_455),
.Y(n_468)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_468),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_453),
.B(n_405),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_471),
.B(n_482),
.Y(n_505)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_445),
.Y(n_474)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_474),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_451),
.B(n_421),
.Y(n_475)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_475),
.Y(n_512)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_459),
.Y(n_476)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_476),
.Y(n_503)
);

FAx1_ASAP7_75t_SL g478 ( 
.A(n_433),
.B(n_411),
.CI(n_391),
.CON(n_478),
.SN(n_478)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_478),
.B(n_486),
.Y(n_499)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_442),
.Y(n_479)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_479),
.Y(n_504)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_445),
.Y(n_481)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_481),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_447),
.B(n_366),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_483),
.A2(n_434),
.B1(n_452),
.B2(n_441),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_428),
.A2(n_358),
.B1(n_387),
.B2(n_422),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_448),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_488),
.B(n_490),
.Y(n_509)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_446),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_492),
.A2(n_500),
.B1(n_510),
.B2(n_515),
.Y(n_532)
);

O2A1O1Ixp33_ASAP7_75t_L g494 ( 
.A1(n_487),
.A2(n_450),
.B(n_438),
.C(n_358),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_494),
.A2(n_502),
.B(n_472),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_469),
.B(n_429),
.C(n_430),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_496),
.B(n_501),
.C(n_506),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_477),
.B(n_429),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_497),
.B(n_507),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_469),
.B(n_436),
.C(n_440),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_487),
.A2(n_438),
.B(n_425),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_464),
.B(n_435),
.C(n_439),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_SL g507 ( 
.A(n_477),
.B(n_444),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_473),
.B(n_449),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_508),
.B(n_473),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_490),
.A2(n_483),
.B1(n_466),
.B2(n_485),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_481),
.B(n_427),
.Y(n_511)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_511),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_464),
.B(n_410),
.C(n_367),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_513),
.B(n_470),
.C(n_489),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_462),
.A2(n_410),
.B1(n_419),
.B2(n_381),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_504),
.B(n_484),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_516),
.B(n_522),
.Y(n_545)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_495),
.Y(n_517)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_517),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_SL g539 ( 
.A(n_518),
.B(n_508),
.Y(n_539)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_495),
.Y(n_519)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_519),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_521),
.B(n_531),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_491),
.B(n_474),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_SL g550 ( 
.A1(n_523),
.A2(n_502),
.B(n_529),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_509),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_524),
.B(n_525),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_504),
.B(n_476),
.Y(n_525)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_514),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_527),
.A2(n_533),
.B1(n_498),
.B2(n_465),
.Y(n_546)
);

CKINVDCx16_ASAP7_75t_R g528 ( 
.A(n_505),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_528),
.B(n_534),
.Y(n_540)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_503),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_530),
.B(n_468),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_514),
.B(n_475),
.Y(n_531)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_503),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_501),
.B(n_472),
.C(n_478),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_SL g535 ( 
.A1(n_527),
.A2(n_510),
.B1(n_492),
.B2(n_509),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_535),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_537),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_520),
.B(n_506),
.C(n_496),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_538),
.B(n_541),
.C(n_542),
.Y(n_556)
);

MAJx2_ASAP7_75t_L g563 ( 
.A(n_539),
.B(n_526),
.C(n_478),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_520),
.B(n_497),
.C(n_500),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_521),
.B(n_513),
.C(n_499),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_522),
.B(n_499),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_543),
.A2(n_544),
.B(n_523),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_534),
.B(n_493),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_546),
.B(n_551),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_550),
.B(n_531),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_532),
.A2(n_515),
.B1(n_511),
.B2(n_512),
.Y(n_551)
);

AOI31xp67_ASAP7_75t_L g571 ( 
.A1(n_552),
.A2(n_560),
.A3(n_562),
.B(n_535),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_545),
.B(n_532),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_557),
.B(n_558),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_548),
.B(n_518),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_559),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_540),
.A2(n_494),
.B(n_519),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_538),
.B(n_507),
.C(n_517),
.Y(n_561)
);

AOI31xp33_ASAP7_75t_L g568 ( 
.A1(n_561),
.A2(n_564),
.A3(n_549),
.B(n_536),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_542),
.A2(n_526),
.B(n_533),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_563),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_548),
.B(n_541),
.C(n_539),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_556),
.A2(n_550),
.B(n_547),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_L g573 ( 
.A1(n_566),
.A2(n_568),
.B(n_571),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_561),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_569),
.B(n_572),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_555),
.B(n_381),
.Y(n_572)
);

INVxp67_ASAP7_75t_L g575 ( 
.A(n_567),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_575),
.B(n_577),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_SL g576 ( 
.A1(n_565),
.A2(n_554),
.B(n_553),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_SL g578 ( 
.A1(n_576),
.A2(n_563),
.B(n_352),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_SL g577 ( 
.A1(n_570),
.A2(n_554),
.B1(n_559),
.B2(n_564),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_578),
.A2(n_579),
.B(n_573),
.Y(n_581)
);

OAI21xp33_ASAP7_75t_L g579 ( 
.A1(n_574),
.A2(n_368),
.B(n_323),
.Y(n_579)
);

OAI21xp5_ASAP7_75t_L g583 ( 
.A1(n_581),
.A2(n_582),
.B(n_266),
.Y(n_583)
);

AOI21xp5_ASAP7_75t_L g582 ( 
.A1(n_580),
.A2(n_368),
.B(n_286),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_583),
.B(n_266),
.Y(n_584)
);


endmodule