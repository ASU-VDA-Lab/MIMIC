module real_jpeg_25456_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_0),
.A2(n_37),
.B1(n_38),
.B2(n_44),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_0),
.A2(n_23),
.B1(n_24),
.B2(n_44),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_0),
.A2(n_44),
.B1(n_51),
.B2(n_55),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_22)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_5),
.A2(n_26),
.B1(n_37),
.B2(n_38),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_6),
.A2(n_37),
.B1(n_38),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_6),
.A2(n_42),
.B1(n_58),
.B2(n_59),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_6),
.A2(n_42),
.B1(n_51),
.B2(n_55),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_42),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_6),
.B(n_51),
.C(n_54),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_6),
.B(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_6),
.B(n_38),
.C(n_67),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_6),
.B(n_24),
.C(n_34),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_6),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_6),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_6),
.B(n_75),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_10),
.Y(n_84)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

OAI22xp5_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_107),
.B1(n_230),
.B2(n_231),
.Y(n_12)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_13),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_106),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_90),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_15),
.B(n_90),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_61),
.C(n_79),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_16),
.A2(n_61),
.B1(n_62),
.B2(n_111),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_16),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_45),
.B2(n_46),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_17),
.A2(n_20),
.B(n_48),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_31),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_19),
.A2(n_20),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_19),
.A2(n_20),
.B1(n_31),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_27),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_22),
.A2(n_28),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_24),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_24),
.B(n_193),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_27),
.B(n_126),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_28),
.A2(n_83),
.B1(n_125),
.B2(n_127),
.Y(n_124)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_29),
.Y(n_128)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_30),
.Y(n_194)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_31),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_40),
.B2(n_43),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_32),
.B(n_33),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_37),
.A2(n_38),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

INVx5_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_38),
.B(n_182),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_41),
.B(n_86),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_63),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_47),
.A2(n_48),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_47),
.A2(n_48),
.B1(n_63),
.B2(n_64),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_47),
.A2(n_48),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_64),
.Y(n_87)
);

AOI211xp5_ASAP7_75t_L g139 ( 
.A1(n_48),
.A2(n_85),
.B(n_89),
.C(n_140),
.Y(n_139)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_60),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_56),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_50),
.B(n_57),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_50),
.Y(n_160)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_51),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_55),
.B1(n_67),
.B2(n_68),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_51),
.B(n_171),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_54),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_58),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_72),
.B(n_78),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_72),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_63),
.B(n_138),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_63),
.A2(n_64),
.B1(n_85),
.B2(n_138),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_63),
.A2(n_64),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_64),
.B(n_143),
.C(n_158),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_64),
.A2(n_85),
.B(n_140),
.C(n_204),
.Y(n_207)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_71),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_66),
.B(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_66),
.A2(n_69),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_66),
.Y(n_188)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_77),
.B(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_78),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_79),
.A2(n_80),
.B1(n_110),
.B2(n_112),
.Y(n_109)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_87),
.B(n_88),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_81),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_81),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_82),
.A2(n_85),
.B1(n_138),
.B2(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_82),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_85),
.A2(n_124),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_85),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_85),
.B(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_85),
.A2(n_138),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_85),
.A2(n_138),
.B1(n_180),
.B2(n_181),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_85),
.A2(n_138),
.B1(n_168),
.B2(n_210),
.Y(n_209)
);

INVxp33_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_87),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_87),
.A2(n_88),
.B(n_142),
.Y(n_221)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_89),
.A2(n_122),
.B(n_129),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_98),
.Y(n_105)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_107),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_130),
.B(n_229),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_113),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_109),
.B(n_113),
.Y(n_229)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.C(n_121),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_114),
.A2(n_115),
.B1(n_119),
.B2(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_116),
.A2(n_117),
.B1(n_142),
.B2(n_149),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_116),
.A2(n_117),
.B1(n_122),
.B2(n_123),
.Y(n_218)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_119),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_121),
.B(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_223),
.B(n_228),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_161),
.B(n_214),
.C(n_222),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_151),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_133),
.B(n_151),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_141),
.B2(n_150),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_136),
.B(n_139),
.C(n_150),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_165),
.C(n_168),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_138),
.B(n_144),
.C(n_187),
.Y(n_201)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_142),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_145),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_143),
.A2(n_144),
.B1(n_158),
.B2(n_159),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_143),
.A2(n_144),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_143),
.B(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_143),
.A2(n_144),
.B1(n_169),
.B2(n_170),
.Y(n_204)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_144),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_144),
.B(n_196),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.C(n_156),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_153),
.A2(n_154),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_174),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_155),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_213),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_175),
.B(n_212),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_172),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_164),
.B(n_172),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_165),
.B(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_168),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_206),
.B(n_211),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_200),
.B(n_205),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_189),
.B(n_199),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_179),
.B(n_183),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_197),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_195),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_201),
.B(n_202),
.Y(n_205)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_207),
.B(n_208),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_216),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_221),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_219),
.C(n_221),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_227),
.Y(n_228)
);


endmodule