module fake_netlist_6_3011_n_1132 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1132);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1132;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_680;
wire n_741;
wire n_1008;
wire n_1027;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_988;
wire n_969;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_1074;
wire n_898;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_1099;
wire n_1026;
wire n_443;
wire n_1101;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_1127;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_222;
wire n_718;
wire n_248;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_1015;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_1116;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_886;
wire n_448;
wire n_953;
wire n_1017;
wire n_1004;
wire n_844;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_1084;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_1121;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_1090;
wire n_592;
wire n_813;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_984;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_1078;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_982;
wire n_964;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_1125;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_518;
wire n_299;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_401;
wire n_324;
wire n_743;
wire n_816;
wire n_766;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_1001;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_1129;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_32),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_176),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_151),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_2),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_139),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_19),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_211),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_0),
.Y(n_226)
);

BUFx8_ASAP7_75t_SL g227 ( 
.A(n_43),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_118),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_158),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_195),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_52),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_101),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_17),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_205),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_13),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_100),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_215),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_97),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_3),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_27),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_209),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_16),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_153),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_22),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_85),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_79),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_50),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_187),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_193),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_61),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_194),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_134),
.Y(n_252)
);

BUFx5_ASAP7_75t_L g253 ( 
.A(n_112),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_28),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_212),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_191),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_110),
.Y(n_257)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_33),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_60),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_44),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_14),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_70),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_125),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_0),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_177),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_159),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_87),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_135),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_5),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_35),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_169),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_173),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_25),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_167),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_53),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_5),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_30),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_69),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_121),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_119),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_150),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_59),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_2),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_47),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_217),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_105),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_109),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_22),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_37),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_92),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_244),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g292 ( 
.A(n_250),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_273),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_253),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_219),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_221),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_273),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_226),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_237),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_250),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_224),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_264),
.Y(n_302)
);

INVxp67_ASAP7_75t_SL g303 ( 
.A(n_277),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_235),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_286),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_242),
.Y(n_306)
);

INVxp33_ASAP7_75t_SL g307 ( 
.A(n_239),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_261),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_269),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_283),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_277),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_220),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_246),
.Y(n_313)
);

INVxp33_ASAP7_75t_SL g314 ( 
.A(n_240),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_222),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_289),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_231),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_227),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_236),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_254),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_276),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_238),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_218),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g324 ( 
.A(n_286),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_233),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_288),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_245),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_225),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_251),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_266),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_271),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_274),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_282),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_285),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_228),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_287),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_290),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_253),
.Y(n_338)
);

INVxp33_ASAP7_75t_SL g339 ( 
.A(n_229),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_304),
.Y(n_340)
);

AOI22x1_ASAP7_75t_SL g341 ( 
.A1(n_295),
.A2(n_234),
.B1(n_241),
.B2(n_230),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_292),
.B(n_223),
.Y(n_342)
);

CKINVDCx11_ASAP7_75t_R g343 ( 
.A(n_318),
.Y(n_343)
);

OAI21x1_ASAP7_75t_L g344 ( 
.A1(n_294),
.A2(n_281),
.B(n_258),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_312),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_317),
.Y(n_346)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_328),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_294),
.Y(n_348)
);

AND2x4_ASAP7_75t_L g349 ( 
.A(n_315),
.B(n_232),
.Y(n_349)
);

BUFx8_ASAP7_75t_SL g350 ( 
.A(n_313),
.Y(n_350)
);

BUFx12f_ASAP7_75t_L g351 ( 
.A(n_328),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_319),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_339),
.B(n_260),
.Y(n_353)
);

INVx5_ASAP7_75t_L g354 ( 
.A(n_320),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_338),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_307),
.A2(n_284),
.B1(n_280),
.B2(n_279),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_338),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_334),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_334),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_336),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_336),
.Y(n_361)
);

INVx6_ASAP7_75t_L g362 ( 
.A(n_322),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_337),
.Y(n_363)
);

INVx6_ASAP7_75t_L g364 ( 
.A(n_327),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_293),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_325),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_337),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_330),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_331),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_332),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_333),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_297),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_304),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_300),
.B(n_278),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_298),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_306),
.Y(n_376)
);

AOI22x1_ASAP7_75t_SL g377 ( 
.A1(n_316),
.A2(n_275),
.B1(n_272),
.B2(n_270),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_291),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_303),
.B(n_268),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_308),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_306),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_309),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_291),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_302),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_339),
.B(n_243),
.Y(n_385)
);

AND2x6_ASAP7_75t_L g386 ( 
.A(n_310),
.B(n_255),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_311),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_329),
.B(n_255),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_302),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_296),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_301),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_335),
.B(n_267),
.Y(n_392)
);

OA21x2_ASAP7_75t_L g393 ( 
.A1(n_320),
.A2(n_248),
.B(n_247),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_326),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_366),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_375),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_348),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_350),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_380),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_350),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_382),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_343),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_348),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_345),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_343),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_351),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_348),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_346),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_352),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_366),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_351),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_370),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_R g413 ( 
.A(n_394),
.B(n_323),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_385),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_394),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_362),
.B(n_335),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_371),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_347),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_347),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_347),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_362),
.B(n_307),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_355),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_341),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_365),
.Y(n_424)
);

INVx2_ASAP7_75t_SL g425 ( 
.A(n_390),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_365),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_341),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_377),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_377),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_392),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_372),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_356),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_362),
.B(n_314),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_354),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_354),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_R g436 ( 
.A(n_391),
.B(n_305),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_372),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_354),
.Y(n_438)
);

INVx6_ASAP7_75t_L g439 ( 
.A(n_362),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_369),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_355),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_354),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_369),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_369),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_354),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_393),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_353),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_390),
.B(n_342),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_387),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_374),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_379),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_364),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_393),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_357),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_342),
.B(n_321),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_364),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_357),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_373),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_393),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_364),
.Y(n_460)
);

INVxp67_ASAP7_75t_SL g461 ( 
.A(n_358),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_364),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_349),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_349),
.Y(n_464)
);

NAND2xp33_ASAP7_75t_R g465 ( 
.A(n_349),
.B(n_326),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_373),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_388),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_388),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_388),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_R g470 ( 
.A(n_340),
.B(n_324),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_414),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_439),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_448),
.B(n_321),
.Y(n_473)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_395),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_450),
.B(n_358),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_424),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_422),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_410),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_452),
.B(n_299),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_426),
.B(n_340),
.Y(n_480)
);

NAND3xp33_ASAP7_75t_L g481 ( 
.A(n_449),
.B(n_368),
.C(n_389),
.Y(n_481)
);

OR2x2_ASAP7_75t_L g482 ( 
.A(n_425),
.B(n_368),
.Y(n_482)
);

OR2x6_ASAP7_75t_L g483 ( 
.A(n_455),
.B(n_381),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_451),
.B(n_358),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_465),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_439),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_439),
.Y(n_487)
);

INVx4_ASAP7_75t_L g488 ( 
.A(n_456),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_441),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_431),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_437),
.B(n_381),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_460),
.B(n_358),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_447),
.B(n_314),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_463),
.Y(n_494)
);

BUFx6f_ASAP7_75t_SL g495 ( 
.A(n_396),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_430),
.A2(n_249),
.B1(n_252),
.B2(n_256),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_399),
.B(n_359),
.Y(n_497)
);

INVx4_ASAP7_75t_L g498 ( 
.A(n_462),
.Y(n_498)
);

OR2x6_ASAP7_75t_L g499 ( 
.A(n_416),
.B(n_359),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_464),
.B(n_358),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_401),
.Y(n_501)
);

INVx4_ASAP7_75t_SL g502 ( 
.A(n_404),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_408),
.Y(n_503)
);

INVx1_ASAP7_75t_SL g504 ( 
.A(n_413),
.Y(n_504)
);

INVx1_ASAP7_75t_SL g505 ( 
.A(n_415),
.Y(n_505)
);

INVxp33_ASAP7_75t_L g506 ( 
.A(n_436),
.Y(n_506)
);

OR2x6_ASAP7_75t_L g507 ( 
.A(n_409),
.B(n_363),
.Y(n_507)
);

BUFx4f_ASAP7_75t_L g508 ( 
.A(n_412),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_467),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_417),
.Y(n_510)
);

INVx8_ASAP7_75t_L g511 ( 
.A(n_406),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_421),
.B(n_360),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_433),
.B(n_378),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_458),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_397),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_441),
.Y(n_516)
);

INVx6_ASAP7_75t_L g517 ( 
.A(n_411),
.Y(n_517)
);

NAND2xp33_ASAP7_75t_L g518 ( 
.A(n_418),
.B(n_253),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_468),
.B(n_363),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_458),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_454),
.Y(n_521)
);

INVxp67_ASAP7_75t_SL g522 ( 
.A(n_422),
.Y(n_522)
);

NAND2xp33_ASAP7_75t_L g523 ( 
.A(n_419),
.B(n_253),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_403),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_454),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_403),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_407),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_407),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_469),
.B(n_367),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_457),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_457),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_461),
.B(n_360),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_422),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_466),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_420),
.B(n_360),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_466),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_440),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_443),
.B(n_444),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_446),
.A2(n_265),
.B1(n_257),
.B2(n_259),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_434),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_SL g541 ( 
.A(n_435),
.B(n_262),
.Y(n_541)
);

AND2x2_ASAP7_75t_SL g542 ( 
.A(n_432),
.B(n_255),
.Y(n_542)
);

AND2x6_ASAP7_75t_L g543 ( 
.A(n_435),
.B(n_255),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_446),
.Y(n_544)
);

NAND3x1_ASAP7_75t_L g545 ( 
.A(n_423),
.B(n_378),
.C(n_1),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_400),
.Y(n_546)
);

INVx1_ASAP7_75t_SL g547 ( 
.A(n_470),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_438),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_442),
.B(n_360),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_445),
.B(n_453),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_459),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_453),
.B(n_360),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_400),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_459),
.B(n_361),
.Y(n_554)
);

AO22x2_ASAP7_75t_L g555 ( 
.A1(n_551),
.A2(n_429),
.B1(n_428),
.B2(n_427),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_489),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_513),
.B(n_361),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_472),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_489),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_516),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_516),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_475),
.B(n_361),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_521),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_521),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_525),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_502),
.B(n_384),
.Y(n_566)
);

AO22x2_ASAP7_75t_L g567 ( 
.A1(n_551),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_525),
.Y(n_568)
);

OAI221xp5_ASAP7_75t_L g569 ( 
.A1(n_485),
.A2(n_367),
.B1(n_384),
.B2(n_378),
.C(n_263),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_530),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_542),
.A2(n_253),
.B1(n_258),
.B2(n_369),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_478),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_493),
.B(n_488),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_473),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_530),
.Y(n_575)
);

INVxp67_ASAP7_75t_L g576 ( 
.A(n_474),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_484),
.B(n_361),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_531),
.Y(n_578)
);

BUFx8_ASAP7_75t_L g579 ( 
.A(n_495),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_519),
.B(n_361),
.Y(n_580)
);

AO22x2_ASAP7_75t_L g581 ( 
.A1(n_544),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_471),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_531),
.Y(n_583)
);

NAND2x1p5_ASAP7_75t_L g584 ( 
.A(n_488),
.B(n_373),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_552),
.A2(n_554),
.B1(n_499),
.B2(n_512),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_502),
.B(n_373),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_497),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_536),
.Y(n_588)
);

OAI221xp5_ASAP7_75t_L g589 ( 
.A1(n_483),
.A2(n_376),
.B1(n_373),
.B2(n_369),
.C(n_383),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_509),
.Y(n_590)
);

A2O1A1Ixp33_ASAP7_75t_L g591 ( 
.A1(n_508),
.A2(n_344),
.B(n_376),
.C(n_383),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_501),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_529),
.B(n_483),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_497),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_491),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_491),
.Y(n_596)
);

INVx1_ASAP7_75t_SL g597 ( 
.A(n_505),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_480),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_480),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_546),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_492),
.B(n_376),
.Y(n_601)
);

AND2x6_ASAP7_75t_L g602 ( 
.A(n_540),
.B(n_376),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_482),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_526),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_543),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_481),
.Y(n_606)
);

OAI221xp5_ASAP7_75t_L g607 ( 
.A1(n_539),
.A2(n_508),
.B1(n_496),
.B2(n_510),
.C(n_503),
.Y(n_607)
);

OAI221xp5_ASAP7_75t_L g608 ( 
.A1(n_507),
.A2(n_376),
.B1(n_383),
.B2(n_398),
.C(n_402),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_541),
.Y(n_609)
);

OR2x2_ASAP7_75t_SL g610 ( 
.A(n_517),
.B(n_405),
.Y(n_610)
);

BUFx8_ASAP7_75t_L g611 ( 
.A(n_495),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_L g612 ( 
.A(n_543),
.B(n_253),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_515),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_526),
.Y(n_614)
);

OAI22xp33_ASAP7_75t_L g615 ( 
.A1(n_499),
.A2(n_383),
.B1(n_258),
.B2(n_8),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_501),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_524),
.Y(n_617)
);

OR2x2_ASAP7_75t_L g618 ( 
.A(n_504),
.B(n_383),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_498),
.B(n_6),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_590),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_573),
.B(n_498),
.Y(n_621)
);

NAND2x1p5_ASAP7_75t_L g622 ( 
.A(n_592),
.B(n_472),
.Y(n_622)
);

A2O1A1Ixp33_ASAP7_75t_L g623 ( 
.A1(n_585),
.A2(n_550),
.B(n_540),
.C(n_548),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_576),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_557),
.A2(n_533),
.B(n_532),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_593),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_607),
.A2(n_580),
.B1(n_574),
.B2(n_606),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_603),
.B(n_501),
.Y(n_628)
);

OR2x6_ASAP7_75t_L g629 ( 
.A(n_592),
.B(n_511),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_562),
.A2(n_533),
.B(n_522),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_577),
.A2(n_477),
.B(n_549),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_592),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_L g633 ( 
.A1(n_591),
.A2(n_528),
.B(n_527),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_601),
.A2(n_535),
.B(n_500),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_L g635 ( 
.A1(n_569),
.A2(n_534),
.B(n_523),
.Y(n_635)
);

NAND3xp33_ASAP7_75t_L g636 ( 
.A(n_572),
.B(n_479),
.C(n_494),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_616),
.Y(n_637)
);

AND2x6_ASAP7_75t_L g638 ( 
.A(n_616),
.B(n_598),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_556),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_589),
.A2(n_518),
.B(n_487),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_583),
.A2(n_487),
.B(n_486),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_597),
.B(n_506),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_609),
.B(n_547),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_582),
.B(n_599),
.Y(n_644)
);

CKINVDCx10_ASAP7_75t_R g645 ( 
.A(n_579),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_559),
.A2(n_486),
.B(n_514),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_560),
.A2(n_520),
.B(n_514),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_588),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_561),
.A2(n_520),
.B(n_514),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_618),
.B(n_600),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_563),
.A2(n_520),
.B(n_538),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_564),
.Y(n_652)
);

OR2x6_ASAP7_75t_L g653 ( 
.A(n_616),
.B(n_511),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_587),
.B(n_476),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_594),
.B(n_507),
.Y(n_655)
);

A2O1A1Ixp33_ASAP7_75t_L g656 ( 
.A1(n_619),
.A2(n_548),
.B(n_490),
.C(n_537),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_565),
.A2(n_538),
.B(n_344),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_568),
.A2(n_543),
.B(n_386),
.Y(n_658)
);

AOI21x1_ASAP7_75t_L g659 ( 
.A1(n_570),
.A2(n_543),
.B(n_258),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_595),
.B(n_545),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_596),
.B(n_517),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_566),
.B(n_553),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_575),
.B(n_578),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_566),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_604),
.A2(n_386),
.B(n_34),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_614),
.A2(n_386),
.B(n_36),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_612),
.A2(n_386),
.B(n_38),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_613),
.Y(n_668)
);

OAI21xp33_ASAP7_75t_L g669 ( 
.A1(n_571),
.A2(n_7),
.B(n_9),
.Y(n_669)
);

CKINVDCx10_ASAP7_75t_R g670 ( 
.A(n_579),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_617),
.A2(n_386),
.B(n_39),
.Y(n_671)
);

OAI22xp5_ASAP7_75t_L g672 ( 
.A1(n_605),
.A2(n_258),
.B1(n_120),
.B2(n_216),
.Y(n_672)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_586),
.A2(n_386),
.B(n_40),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_610),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_608),
.B(n_10),
.Y(n_675)
);

INVx4_ASAP7_75t_L g676 ( 
.A(n_586),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_558),
.B(n_602),
.Y(n_677)
);

O2A1O1Ixp5_ASAP7_75t_L g678 ( 
.A1(n_615),
.A2(n_602),
.B(n_584),
.C(n_567),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_602),
.B(n_10),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_602),
.A2(n_41),
.B(n_31),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_581),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_567),
.A2(n_45),
.B(n_42),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_581),
.A2(n_48),
.B(n_46),
.Y(n_683)
);

O2A1O1Ixp5_ASAP7_75t_L g684 ( 
.A1(n_621),
.A2(n_555),
.B(n_12),
.C(n_13),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_625),
.A2(n_631),
.B(n_635),
.Y(n_685)
);

NAND3xp33_ASAP7_75t_L g686 ( 
.A(n_675),
.B(n_611),
.C(n_555),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_650),
.B(n_611),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_644),
.B(n_11),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_639),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_627),
.B(n_11),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_638),
.Y(n_691)
);

OAI22xp5_ASAP7_75t_L g692 ( 
.A1(n_623),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_652),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_628),
.B(n_15),
.Y(n_694)
);

AOI22x1_ASAP7_75t_L g695 ( 
.A1(n_640),
.A2(n_127),
.B1(n_213),
.B2(n_210),
.Y(n_695)
);

NOR3xp33_ASAP7_75t_L g696 ( 
.A(n_642),
.B(n_16),
.C(n_17),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_630),
.A2(n_51),
.B(n_49),
.Y(n_697)
);

AOI22x1_ASAP7_75t_L g698 ( 
.A1(n_634),
.A2(n_129),
.B1(n_208),
.B2(n_207),
.Y(n_698)
);

OR2x6_ASAP7_75t_L g699 ( 
.A(n_629),
.B(n_653),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_648),
.Y(n_700)
);

BUFx4f_ASAP7_75t_L g701 ( 
.A(n_629),
.Y(n_701)
);

O2A1O1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_656),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_SL g703 ( 
.A(n_620),
.B(n_54),
.Y(n_703)
);

BUFx2_ASAP7_75t_L g704 ( 
.A(n_626),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_643),
.B(n_18),
.Y(n_705)
);

BUFx4f_ASAP7_75t_L g706 ( 
.A(n_653),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_654),
.B(n_20),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_633),
.A2(n_130),
.B(n_206),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_668),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_663),
.B(n_21),
.Y(n_710)
);

O2A1O1Ixp33_ASAP7_75t_L g711 ( 
.A1(n_678),
.A2(n_21),
.B(n_23),
.C(n_24),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_655),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_624),
.B(n_23),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_657),
.A2(n_131),
.B(n_204),
.Y(n_714)
);

A2O1A1Ixp33_ASAP7_75t_L g715 ( 
.A1(n_669),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_715)
);

OAI21xp33_ASAP7_75t_L g716 ( 
.A1(n_660),
.A2(n_26),
.B(n_27),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_664),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_SL g718 ( 
.A(n_676),
.B(n_55),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_636),
.B(n_28),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_662),
.B(n_29),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_651),
.A2(n_136),
.B(n_56),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_622),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_681),
.B(n_29),
.Y(n_723)
);

OAI21xp33_ASAP7_75t_L g724 ( 
.A1(n_661),
.A2(n_57),
.B(n_58),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_647),
.A2(n_62),
.B(n_63),
.Y(n_725)
);

A2O1A1Ixp33_ASAP7_75t_L g726 ( 
.A1(n_682),
.A2(n_683),
.B(n_658),
.C(n_641),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_637),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_637),
.Y(n_728)
);

BUFx2_ASAP7_75t_L g729 ( 
.A(n_632),
.Y(n_729)
);

AND2x6_ASAP7_75t_L g730 ( 
.A(n_637),
.B(n_64),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_632),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_638),
.B(n_65),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_638),
.Y(n_733)
);

A2O1A1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_649),
.A2(n_66),
.B(n_67),
.C(n_68),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_674),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_638),
.B(n_74),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_679),
.B(n_214),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_677),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_646),
.B(n_75),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_SL g740 ( 
.A1(n_672),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_L g741 ( 
.A1(n_680),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_741)
);

O2A1O1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_671),
.A2(n_83),
.B(n_84),
.C(n_86),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_R g743 ( 
.A(n_645),
.B(n_88),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_743),
.Y(n_744)
);

INVxp67_ASAP7_75t_SL g745 ( 
.A(n_689),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_738),
.B(n_659),
.Y(n_746)
);

INVx4_ASAP7_75t_L g747 ( 
.A(n_701),
.Y(n_747)
);

BUFx12f_ASAP7_75t_L g748 ( 
.A(n_699),
.Y(n_748)
);

INVxp67_ASAP7_75t_SL g749 ( 
.A(n_693),
.Y(n_749)
);

BUFx2_ASAP7_75t_SL g750 ( 
.A(n_729),
.Y(n_750)
);

INVx1_ASAP7_75t_SL g751 ( 
.A(n_704),
.Y(n_751)
);

INVxp67_ASAP7_75t_SL g752 ( 
.A(n_709),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_690),
.B(n_673),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_719),
.B(n_670),
.Y(n_754)
);

INVx4_ASAP7_75t_L g755 ( 
.A(n_701),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_691),
.Y(n_756)
);

INVxp67_ASAP7_75t_SL g757 ( 
.A(n_685),
.Y(n_757)
);

INVx5_ASAP7_75t_L g758 ( 
.A(n_730),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_706),
.Y(n_759)
);

BUFx4_ASAP7_75t_SL g760 ( 
.A(n_699),
.Y(n_760)
);

INVx5_ASAP7_75t_SL g761 ( 
.A(n_731),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_696),
.A2(n_716),
.B1(n_692),
.B2(n_688),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_712),
.B(n_722),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_707),
.A2(n_667),
.B1(n_666),
.B2(n_665),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_705),
.B(n_89),
.Y(n_765)
);

BUFx2_ASAP7_75t_SL g766 ( 
.A(n_728),
.Y(n_766)
);

INVx5_ASAP7_75t_L g767 ( 
.A(n_730),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_706),
.Y(n_768)
);

BUFx2_ASAP7_75t_L g769 ( 
.A(n_727),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_717),
.Y(n_770)
);

BUFx8_ASAP7_75t_L g771 ( 
.A(n_730),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_710),
.B(n_90),
.Y(n_772)
);

BUFx12f_ASAP7_75t_L g773 ( 
.A(n_730),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_720),
.B(n_91),
.Y(n_774)
);

INVx1_ASAP7_75t_SL g775 ( 
.A(n_694),
.Y(n_775)
);

BUFx2_ASAP7_75t_L g776 ( 
.A(n_700),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_691),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_687),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_733),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_732),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_723),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_695),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_737),
.B(n_715),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_698),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_736),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_711),
.Y(n_786)
);

INVxp67_ASAP7_75t_SL g787 ( 
.A(n_702),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_713),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_684),
.Y(n_789)
);

BUFx12f_ASAP7_75t_L g790 ( 
.A(n_703),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_739),
.Y(n_791)
);

BUFx3_ASAP7_75t_L g792 ( 
.A(n_686),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_718),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_735),
.Y(n_794)
);

INVxp67_ASAP7_75t_SL g795 ( 
.A(n_708),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_741),
.Y(n_796)
);

AO22x2_ASAP7_75t_L g797 ( 
.A1(n_714),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_734),
.Y(n_798)
);

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_740),
.Y(n_799)
);

BUFx8_ASAP7_75t_L g800 ( 
.A(n_724),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_721),
.Y(n_801)
);

BUFx2_ASAP7_75t_SL g802 ( 
.A(n_725),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_726),
.B(n_96),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_697),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_742),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_738),
.B(n_203),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_701),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_738),
.B(n_98),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_699),
.B(n_99),
.Y(n_809)
);

BUFx8_ASAP7_75t_L g810 ( 
.A(n_729),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_689),
.Y(n_811)
);

BUFx2_ASAP7_75t_L g812 ( 
.A(n_704),
.Y(n_812)
);

OAI21x1_ASAP7_75t_L g813 ( 
.A1(n_784),
.A2(n_102),
.B(n_103),
.Y(n_813)
);

OAI21x1_ASAP7_75t_L g814 ( 
.A1(n_782),
.A2(n_104),
.B(n_106),
.Y(n_814)
);

NAND2x1p5_ASAP7_75t_L g815 ( 
.A(n_758),
.B(n_107),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_762),
.A2(n_202),
.B1(n_111),
.B2(n_113),
.Y(n_816)
);

OAI21x1_ASAP7_75t_L g817 ( 
.A1(n_757),
.A2(n_108),
.B(n_114),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_776),
.B(n_115),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_745),
.B(n_116),
.Y(n_819)
);

OA21x2_ASAP7_75t_L g820 ( 
.A1(n_789),
.A2(n_795),
.B(n_757),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_744),
.Y(n_821)
);

AOI21x1_ASAP7_75t_L g822 ( 
.A1(n_783),
.A2(n_117),
.B(n_122),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_810),
.Y(n_823)
);

BUFx3_ASAP7_75t_L g824 ( 
.A(n_810),
.Y(n_824)
);

OAI22xp33_ASAP7_75t_L g825 ( 
.A1(n_799),
.A2(n_123),
.B1(n_124),
.B2(n_126),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_749),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_783),
.A2(n_128),
.B(n_132),
.C(n_133),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_762),
.A2(n_137),
.B1(n_138),
.B2(n_140),
.Y(n_828)
);

OAI21x1_ASAP7_75t_L g829 ( 
.A1(n_746),
.A2(n_141),
.B(n_142),
.Y(n_829)
);

AOI22x1_ASAP7_75t_L g830 ( 
.A1(n_797),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_830)
);

OA21x2_ASAP7_75t_L g831 ( 
.A1(n_795),
.A2(n_146),
.B(n_147),
.Y(n_831)
);

NOR2x1_ASAP7_75t_SL g832 ( 
.A(n_758),
.B(n_767),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_749),
.B(n_148),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_R g834 ( 
.A(n_758),
.B(n_149),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_752),
.B(n_152),
.Y(n_835)
);

OAI21x1_ASAP7_75t_L g836 ( 
.A1(n_803),
.A2(n_154),
.B(n_155),
.Y(n_836)
);

OAI21xp33_ASAP7_75t_SL g837 ( 
.A1(n_772),
.A2(n_156),
.B(n_157),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_758),
.B(n_160),
.Y(n_838)
);

O2A1O1Ixp33_ASAP7_75t_SL g839 ( 
.A1(n_794),
.A2(n_161),
.B(n_162),
.C(n_163),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_811),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_787),
.A2(n_201),
.B1(n_165),
.B2(n_166),
.Y(n_841)
);

NOR2xp67_ASAP7_75t_L g842 ( 
.A(n_747),
.B(n_164),
.Y(n_842)
);

AO31x2_ASAP7_75t_L g843 ( 
.A1(n_786),
.A2(n_168),
.A3(n_170),
.B(n_171),
.Y(n_843)
);

AOI21x1_ASAP7_75t_L g844 ( 
.A1(n_753),
.A2(n_172),
.B(n_174),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_804),
.A2(n_175),
.B(n_178),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_769),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_791),
.B(n_179),
.Y(n_847)
);

OAI21x1_ASAP7_75t_L g848 ( 
.A1(n_798),
.A2(n_180),
.B(n_181),
.Y(n_848)
);

AO21x2_ASAP7_75t_L g849 ( 
.A1(n_787),
.A2(n_182),
.B(n_183),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_763),
.Y(n_850)
);

AO21x2_ASAP7_75t_L g851 ( 
.A1(n_753),
.A2(n_184),
.B(n_185),
.Y(n_851)
);

INVx6_ASAP7_75t_L g852 ( 
.A(n_771),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_777),
.Y(n_853)
);

NAND2x1p5_ASAP7_75t_L g854 ( 
.A(n_767),
.B(n_793),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_788),
.B(n_186),
.Y(n_855)
);

OAI21x1_ASAP7_75t_L g856 ( 
.A1(n_798),
.A2(n_188),
.B(n_189),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_812),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_775),
.B(n_190),
.Y(n_858)
);

NAND2x1p5_ASAP7_75t_L g859 ( 
.A(n_767),
.B(n_192),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_797),
.A2(n_196),
.B(n_197),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_799),
.A2(n_198),
.B1(n_200),
.B2(n_781),
.Y(n_861)
);

OAI22xp5_ASAP7_75t_L g862 ( 
.A1(n_767),
.A2(n_797),
.B1(n_775),
.B2(n_790),
.Y(n_862)
);

OAI21x1_ASAP7_75t_L g863 ( 
.A1(n_764),
.A2(n_808),
.B(n_806),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_770),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_777),
.Y(n_865)
);

OAI21x1_ASAP7_75t_L g866 ( 
.A1(n_764),
.A2(n_808),
.B(n_806),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_779),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_780),
.B(n_785),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_759),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_840),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_820),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_826),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_826),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_852),
.Y(n_874)
);

OA21x2_ASAP7_75t_L g875 ( 
.A1(n_863),
.A2(n_772),
.B(n_796),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_868),
.B(n_751),
.Y(n_876)
);

CKINVDCx8_ASAP7_75t_R g877 ( 
.A(n_869),
.Y(n_877)
);

INVx3_ASAP7_75t_L g878 ( 
.A(n_854),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_846),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_825),
.A2(n_792),
.B1(n_805),
.B2(n_800),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_866),
.Y(n_881)
);

HB1xp67_ASAP7_75t_L g882 ( 
.A(n_868),
.Y(n_882)
);

INVxp67_ASAP7_75t_L g883 ( 
.A(n_857),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_843),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_854),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_843),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_843),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_825),
.A2(n_805),
.B1(n_800),
.B2(n_793),
.Y(n_888)
);

OAI21x1_ASAP7_75t_L g889 ( 
.A1(n_829),
.A2(n_756),
.B(n_802),
.Y(n_889)
);

NAND2x1p5_ASAP7_75t_L g890 ( 
.A(n_830),
.B(n_801),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_843),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_861),
.A2(n_805),
.B1(n_774),
.B2(n_765),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_852),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_831),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_L g895 ( 
.A1(n_861),
.A2(n_765),
.B1(n_754),
.B2(n_773),
.Y(n_895)
);

INVx1_ASAP7_75t_SL g896 ( 
.A(n_869),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_864),
.Y(n_897)
);

OAI21x1_ASAP7_75t_L g898 ( 
.A1(n_817),
.A2(n_801),
.B(n_785),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_831),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_850),
.B(n_780),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_819),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_852),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_858),
.B(n_751),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_867),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_851),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_862),
.A2(n_754),
.B1(n_748),
.B2(n_809),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_819),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_833),
.Y(n_908)
);

OR2x2_ASAP7_75t_L g909 ( 
.A(n_862),
.B(n_780),
.Y(n_909)
);

INVxp67_ASAP7_75t_L g910 ( 
.A(n_869),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_880),
.A2(n_828),
.B1(n_816),
.B2(n_841),
.Y(n_911)
);

NAND3xp33_ASAP7_75t_SL g912 ( 
.A(n_895),
.B(n_888),
.C(n_860),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_893),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_871),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_870),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_870),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_893),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_882),
.B(n_778),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_R g919 ( 
.A(n_877),
.B(n_771),
.Y(n_919)
);

OR2x6_ASAP7_75t_L g920 ( 
.A(n_909),
.B(n_860),
.Y(n_920)
);

AND2x2_ASAP7_75t_SL g921 ( 
.A(n_875),
.B(n_838),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_879),
.B(n_824),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_897),
.B(n_823),
.Y(n_923)
);

NOR3xp33_ASAP7_75t_SL g924 ( 
.A(n_903),
.B(n_855),
.C(n_847),
.Y(n_924)
);

INVx8_ASAP7_75t_L g925 ( 
.A(n_893),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_872),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_871),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_904),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_892),
.A2(n_828),
.B1(n_816),
.B2(n_841),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_901),
.B(n_785),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_883),
.B(n_855),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_872),
.Y(n_932)
);

OR2x6_ASAP7_75t_L g933 ( 
.A(n_909),
.B(n_815),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_873),
.B(n_835),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_R g935 ( 
.A(n_877),
.B(n_821),
.Y(n_935)
);

OR2x2_ASAP7_75t_L g936 ( 
.A(n_901),
.B(n_833),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_893),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_874),
.Y(n_938)
);

NAND2xp33_ASAP7_75t_L g939 ( 
.A(n_893),
.B(n_834),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_874),
.Y(n_940)
);

BUFx4f_ASAP7_75t_SL g941 ( 
.A(n_896),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_907),
.B(n_858),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_900),
.B(n_832),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_937),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_937),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_921),
.B(n_918),
.Y(n_946)
);

INVx2_ASAP7_75t_SL g947 ( 
.A(n_940),
.Y(n_947)
);

OR2x2_ASAP7_75t_L g948 ( 
.A(n_934),
.B(n_884),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_942),
.B(n_907),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_942),
.B(n_908),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_914),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_936),
.B(n_908),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_914),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_937),
.Y(n_954)
);

OR2x2_ASAP7_75t_L g955 ( 
.A(n_927),
.B(n_884),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_927),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_930),
.B(n_876),
.Y(n_957)
);

AOI211x1_ASAP7_75t_L g958 ( 
.A1(n_912),
.A2(n_845),
.B(n_822),
.C(n_886),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_926),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_932),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_921),
.B(n_875),
.Y(n_961)
);

OR2x2_ASAP7_75t_L g962 ( 
.A(n_916),
.B(n_891),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_928),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_915),
.Y(n_964)
);

OA21x2_ASAP7_75t_L g965 ( 
.A1(n_924),
.A2(n_881),
.B(n_886),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_943),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_922),
.B(n_875),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_962),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_955),
.Y(n_969)
);

CKINVDCx20_ASAP7_75t_R g970 ( 
.A(n_957),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_965),
.A2(n_924),
.B(n_912),
.Y(n_971)
);

OA21x2_ASAP7_75t_L g972 ( 
.A1(n_961),
.A2(n_881),
.B(n_894),
.Y(n_972)
);

AOI21xp33_ASAP7_75t_L g973 ( 
.A1(n_965),
.A2(n_920),
.B(n_929),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_948),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_949),
.A2(n_911),
.B(n_920),
.C(n_939),
.Y(n_975)
);

OAI22xp33_ASAP7_75t_L g976 ( 
.A1(n_946),
.A2(n_906),
.B1(n_920),
.B2(n_933),
.Y(n_976)
);

HB1xp67_ASAP7_75t_L g977 ( 
.A(n_948),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_962),
.Y(n_978)
);

AOI22xp33_ASAP7_75t_L g979 ( 
.A1(n_946),
.A2(n_933),
.B1(n_923),
.B2(n_838),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_945),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_967),
.B(n_940),
.Y(n_981)
);

INVxp67_ASAP7_75t_L g982 ( 
.A(n_950),
.Y(n_982)
);

BUFx3_ASAP7_75t_L g983 ( 
.A(n_945),
.Y(n_983)
);

AOI22xp33_ASAP7_75t_L g984 ( 
.A1(n_965),
.A2(n_933),
.B1(n_931),
.B2(n_849),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_967),
.B(n_913),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_955),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_980),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_972),
.Y(n_988)
);

INVx3_ASAP7_75t_SL g989 ( 
.A(n_980),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_982),
.B(n_960),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_968),
.B(n_960),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_968),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_978),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_980),
.Y(n_994)
);

INVx1_ASAP7_75t_SL g995 ( 
.A(n_970),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_978),
.Y(n_996)
);

OR2x2_ASAP7_75t_L g997 ( 
.A(n_973),
.B(n_952),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_981),
.B(n_966),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_974),
.Y(n_999)
);

INVx2_ASAP7_75t_SL g1000 ( 
.A(n_983),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_999),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_997),
.B(n_971),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_988),
.Y(n_1003)
);

NAND2xp33_ASAP7_75t_R g1004 ( 
.A(n_987),
.B(n_935),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_989),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_989),
.B(n_983),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_999),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_994),
.B(n_981),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_992),
.Y(n_1009)
);

OR2x2_ASAP7_75t_L g1010 ( 
.A(n_990),
.B(n_971),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_1005),
.B(n_1000),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_1006),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_1001),
.B(n_995),
.Y(n_1013)
);

INVx2_ASAP7_75t_SL g1014 ( 
.A(n_1006),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_1008),
.B(n_998),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_1007),
.Y(n_1016)
);

NAND2xp33_ASAP7_75t_L g1017 ( 
.A(n_1010),
.B(n_935),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_1009),
.B(n_993),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_1013),
.B(n_1002),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_1018),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1018),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_1011),
.B(n_983),
.Y(n_1022)
);

BUFx2_ASAP7_75t_L g1023 ( 
.A(n_1014),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_1012),
.Y(n_1024)
);

INVx1_ASAP7_75t_SL g1025 ( 
.A(n_1017),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_1015),
.B(n_996),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1016),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_1012),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1018),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_1023),
.B(n_1028),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_1025),
.B(n_990),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1028),
.B(n_991),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_1024),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_1019),
.B(n_975),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_1022),
.B(n_1026),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1024),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1028),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_1027),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_1034),
.A2(n_1019),
.B1(n_1021),
.B2(n_1020),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1033),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_1030),
.A2(n_1029),
.B1(n_979),
.B2(n_976),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_SL g1042 ( 
.A1(n_1031),
.A2(n_984),
.B(n_1004),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1036),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_1035),
.B(n_991),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1037),
.Y(n_1045)
);

NOR2xp67_ASAP7_75t_SL g1046 ( 
.A(n_1038),
.B(n_768),
.Y(n_1046)
);

INVx2_ASAP7_75t_SL g1047 ( 
.A(n_1040),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1043),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_1039),
.A2(n_1032),
.B(n_1038),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_1045),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_1044),
.B(n_969),
.Y(n_1051)
);

NAND2x1_ASAP7_75t_L g1052 ( 
.A(n_1047),
.B(n_1046),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_1050),
.B(n_1041),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1048),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1051),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_1049),
.B(n_1003),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_1047),
.B(n_1042),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_SL g1058 ( 
.A1(n_1053),
.A2(n_902),
.B(n_1003),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1057),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1056),
.Y(n_1060)
);

NAND2xp33_ASAP7_75t_L g1061 ( 
.A(n_1054),
.B(n_1004),
.Y(n_1061)
);

AOI211x1_ASAP7_75t_L g1062 ( 
.A1(n_1055),
.A2(n_985),
.B(n_961),
.C(n_953),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_1052),
.A2(n_919),
.B1(n_902),
.B2(n_988),
.Y(n_1063)
);

AOI221xp5_ASAP7_75t_L g1064 ( 
.A1(n_1061),
.A2(n_958),
.B1(n_839),
.B2(n_837),
.C(n_938),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_1059),
.A2(n_910),
.B1(n_941),
.B2(n_755),
.Y(n_1065)
);

AOI221x1_ASAP7_75t_L g1066 ( 
.A1(n_1060),
.A2(n_747),
.B1(n_755),
.B2(n_809),
.C(n_845),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1058),
.B(n_969),
.Y(n_1067)
);

O2A1O1Ixp5_ASAP7_75t_L g1068 ( 
.A1(n_1067),
.A2(n_1063),
.B(n_1062),
.C(n_969),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1065),
.Y(n_1069)
);

OAI211xp5_ASAP7_75t_L g1070 ( 
.A1(n_1066),
.A2(n_919),
.B(n_834),
.C(n_807),
.Y(n_1070)
);

INVx1_ASAP7_75t_SL g1071 ( 
.A(n_1064),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_1067),
.A2(n_839),
.B(n_827),
.C(n_859),
.Y(n_1072)
);

OAI221xp5_ASAP7_75t_L g1073 ( 
.A1(n_1067),
.A2(n_859),
.B1(n_815),
.B2(n_750),
.C(n_842),
.Y(n_1073)
);

CKINVDCx20_ASAP7_75t_R g1074 ( 
.A(n_1065),
.Y(n_1074)
);

OAI211xp5_ASAP7_75t_SL g1075 ( 
.A1(n_1067),
.A2(n_760),
.B(n_847),
.C(n_835),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_1069),
.A2(n_954),
.B1(n_945),
.B2(n_941),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1071),
.B(n_986),
.Y(n_1077)
);

INVx1_ASAP7_75t_SL g1078 ( 
.A(n_1074),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_1070),
.A2(n_760),
.B(n_849),
.C(n_977),
.Y(n_1079)
);

OAI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_1073),
.A2(n_986),
.B1(n_954),
.B2(n_944),
.Y(n_1080)
);

OAI211xp5_ASAP7_75t_SL g1081 ( 
.A1(n_1068),
.A2(n_944),
.B(n_986),
.C(n_917),
.Y(n_1081)
);

OR2x2_ASAP7_75t_L g1082 ( 
.A(n_1075),
.B(n_972),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_1072),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1069),
.B(n_944),
.Y(n_1084)
);

AOI311xp33_ASAP7_75t_L g1085 ( 
.A1(n_1069),
.A2(n_951),
.A3(n_956),
.B(n_953),
.C(n_887),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_1078),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1076),
.B(n_944),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1077),
.Y(n_1088)
);

OAI211xp5_ASAP7_75t_L g1089 ( 
.A1(n_1084),
.A2(n_818),
.B(n_958),
.C(n_972),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_1079),
.A2(n_954),
.B(n_947),
.C(n_985),
.Y(n_1090)
);

AND3x2_ASAP7_75t_L g1091 ( 
.A(n_1083),
.B(n_951),
.C(n_956),
.Y(n_1091)
);

NOR2x1_ASAP7_75t_L g1092 ( 
.A(n_1081),
.B(n_766),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_1082),
.Y(n_1093)
);

NOR3xp33_ASAP7_75t_L g1094 ( 
.A(n_1080),
.B(n_844),
.C(n_856),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1085),
.A2(n_947),
.B1(n_972),
.B2(n_937),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_1078),
.B(n_966),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_1078),
.B(n_917),
.Y(n_1097)
);

NOR2x1_ASAP7_75t_L g1098 ( 
.A(n_1078),
.B(n_965),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_1091),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1086),
.Y(n_1100)
);

NOR2x1_ASAP7_75t_L g1101 ( 
.A(n_1088),
.B(n_1093),
.Y(n_1101)
);

XNOR2xp5_ASAP7_75t_L g1102 ( 
.A(n_1097),
.B(n_848),
.Y(n_1102)
);

CKINVDCx20_ASAP7_75t_R g1103 ( 
.A(n_1087),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_1096),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_1095),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_1092),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1099),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1100),
.Y(n_1108)
);

XNOR2x1_ASAP7_75t_L g1109 ( 
.A(n_1104),
.B(n_1098),
.Y(n_1109)
);

NOR3xp33_ASAP7_75t_SL g1110 ( 
.A(n_1106),
.B(n_1090),
.C(n_1089),
.Y(n_1110)
);

OA22x2_ASAP7_75t_L g1111 ( 
.A1(n_1102),
.A2(n_1094),
.B1(n_913),
.B2(n_814),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1105),
.A2(n_761),
.B1(n_959),
.B2(n_925),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1101),
.A2(n_925),
.B(n_836),
.Y(n_1113)
);

OAI221xp5_ASAP7_75t_L g1114 ( 
.A1(n_1107),
.A2(n_1103),
.B1(n_959),
.B2(n_890),
.C(n_878),
.Y(n_1114)
);

OR2x2_ASAP7_75t_L g1115 ( 
.A(n_1108),
.B(n_761),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1112),
.A2(n_925),
.B1(n_761),
.B2(n_885),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1115),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1117),
.Y(n_1118)
);

OAI21xp33_ASAP7_75t_SL g1119 ( 
.A1(n_1118),
.A2(n_1109),
.B(n_1116),
.Y(n_1119)
);

OAI322xp33_ASAP7_75t_L g1120 ( 
.A1(n_1119),
.A2(n_1114),
.A3(n_1110),
.B1(n_1111),
.B2(n_1113),
.C1(n_777),
.C2(n_887),
.Y(n_1120)
);

OAI322xp33_ASAP7_75t_L g1121 ( 
.A1(n_1119),
.A2(n_891),
.A3(n_865),
.B1(n_853),
.B2(n_964),
.C1(n_963),
.C2(n_894),
.Y(n_1121)
);

XNOR2xp5_ASAP7_75t_L g1122 ( 
.A(n_1119),
.B(n_813),
.Y(n_1122)
);

AOI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_1122),
.A2(n_1120),
.B1(n_1121),
.B2(n_905),
.Y(n_1123)
);

OAI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1120),
.A2(n_885),
.B1(n_878),
.B2(n_865),
.Y(n_1124)
);

OR2x2_ASAP7_75t_L g1125 ( 
.A(n_1122),
.B(n_964),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_1125),
.A2(n_1123),
.B1(n_1124),
.B2(n_904),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1125),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1124),
.A2(n_885),
.B1(n_878),
.B2(n_963),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1127),
.A2(n_889),
.B(n_898),
.Y(n_1129)
);

AO21x2_ASAP7_75t_L g1130 ( 
.A1(n_1128),
.A2(n_899),
.B(n_889),
.Y(n_1130)
);

OAI211xp5_ASAP7_75t_L g1131 ( 
.A1(n_1129),
.A2(n_1126),
.B(n_853),
.C(n_905),
.Y(n_1131)
);

AOI211xp5_ASAP7_75t_L g1132 ( 
.A1(n_1131),
.A2(n_1130),
.B(n_779),
.C(n_899),
.Y(n_1132)
);


endmodule