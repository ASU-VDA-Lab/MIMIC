module fake_jpeg_29915_n_194 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_194);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_194;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx10_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_1),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_20),
.B(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_2),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_43),
.Y(n_51)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_15),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_15),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_55),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_28),
.B1(n_24),
.B2(n_23),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_58),
.B1(n_61),
.B2(n_14),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_12),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_25),
.B1(n_27),
.B2(n_18),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_18),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_66),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_29),
.A2(n_25),
.B1(n_17),
.B2(n_14),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_34),
.A2(n_23),
.B1(n_21),
.B2(n_19),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_29),
.A2(n_21),
.B1(n_19),
.B2(n_16),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_64),
.A2(n_13),
.B1(n_16),
.B2(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_17),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_69),
.A2(n_93),
.B(n_36),
.C(n_65),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_40),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_80),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_43),
.B1(n_35),
.B2(n_33),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_75),
.A2(n_31),
.B1(n_33),
.B2(n_65),
.Y(n_104)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_48),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_77),
.B(n_78),
.Y(n_106)
);

NOR2x1_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_13),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_46),
.B(n_12),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_84),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_31),
.Y(n_80)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_37),
.Y(n_84)
);

BUFx8_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_37),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_87),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_48),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_49),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_92),
.Y(n_115)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_94),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_12),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_SL g93 ( 
.A1(n_44),
.A2(n_12),
.B(n_43),
.C(n_35),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_4),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_44),
.B(n_65),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_97),
.Y(n_118)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_12),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

HAxp5_ASAP7_75t_SL g99 ( 
.A(n_60),
.B(n_5),
.CON(n_99),
.SN(n_99)
);

XNOR2x1_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_6),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_54),
.B(n_31),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_54),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_102),
.A2(n_109),
.B1(n_80),
.B2(n_74),
.Y(n_135)
);

AO22x1_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_69),
.B1(n_99),
.B2(n_72),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_91),
.A2(n_54),
.B1(n_36),
.B2(n_8),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_88),
.A2(n_91),
.B1(n_69),
.B2(n_93),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_113),
.A2(n_88),
.B1(n_72),
.B2(n_94),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_70),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_116),
.B(n_122),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_119),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_6),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_82),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_130),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_127),
.A2(n_131),
.B(n_102),
.Y(n_153)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

AND2x6_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_78),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_140),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_101),
.A2(n_81),
.B1(n_80),
.B2(n_71),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_133),
.A2(n_135),
.B1(n_124),
.B2(n_101),
.Y(n_144)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_136),
.B(n_137),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_122),
.B(n_7),
.Y(n_137)
);

A2O1A1O1Ixp25_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_97),
.B(n_95),
.C(n_69),
.D(n_100),
.Y(n_138)
);

OAI21x1_ASAP7_75t_L g154 ( 
.A1(n_138),
.A2(n_103),
.B(n_114),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_111),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_118),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_146),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_115),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_148),
.C(n_152),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_144),
.A2(n_129),
.B1(n_138),
.B2(n_130),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_118),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_120),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_120),
.C(n_119),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_153),
.B(n_135),
.Y(n_156)
);

FAx1_ASAP7_75t_SL g161 ( 
.A(n_154),
.B(n_148),
.CI(n_141),
.CON(n_161),
.SN(n_161)
);

XNOR2x1_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_163),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_158),
.A2(n_129),
.B1(n_142),
.B2(n_100),
.Y(n_171)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_159),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_136),
.C(n_114),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_164),
.C(n_166),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_123),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

OAI21xp33_ASAP7_75t_L g163 ( 
.A1(n_146),
.A2(n_105),
.B(n_123),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_121),
.C(n_117),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_121),
.C(n_105),
.Y(n_166)
);

AOI321xp33_ASAP7_75t_L g168 ( 
.A1(n_155),
.A2(n_132),
.A3(n_150),
.B1(n_145),
.B2(n_151),
.C(n_147),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_165),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_171),
.A2(n_166),
.B1(n_164),
.B2(n_170),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_90),
.B1(n_108),
.B2(n_83),
.Y(n_174)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_174),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_155),
.B(n_108),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_85),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_178),
.C(n_181),
.Y(n_182)
);

AOI31xp67_ASAP7_75t_L g177 ( 
.A1(n_172),
.A2(n_161),
.A3(n_163),
.B(n_160),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_177),
.A2(n_180),
.B(n_173),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_173),
.A2(n_165),
.B(n_8),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_181),
.B(n_167),
.C(n_175),
.Y(n_183)
);

OAI221xp5_ASAP7_75t_L g188 ( 
.A1(n_183),
.A2(n_85),
.B1(n_10),
.B2(n_11),
.C(n_7),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_184),
.A2(n_185),
.B1(n_7),
.B2(n_10),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_169),
.B(n_172),
.Y(n_185)
);

NAND3xp33_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_179),
.C(n_9),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_186),
.B(n_188),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_187),
.B(n_10),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_189),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_11),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_190),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_193),
.A2(n_192),
.B(n_11),
.Y(n_194)
);


endmodule