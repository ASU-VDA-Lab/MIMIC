module fake_jpeg_25710_n_83 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_83);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_83;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

HB1xp67_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_19),
.Y(n_22)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_20),
.A2(n_13),
.B1(n_14),
.B2(n_12),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_23),
.B1(n_24),
.B2(n_19),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_20),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_27),
.B(n_33),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

OAI21xp33_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_30),
.B(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_10),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_9),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_40),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_38),
.A2(n_39),
.B1(n_32),
.B2(n_18),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_25),
.Y(n_54)
);

BUFx24_ASAP7_75t_SL g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_54),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_53),
.B1(n_35),
.B2(n_43),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_18),
.C(n_17),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_51),
.C(n_52),
.Y(n_57)
);

AO22x1_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_34),
.B1(n_25),
.B2(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_17),
.C(n_16),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_17),
.C(n_26),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_25),
.B1(n_15),
.B2(n_0),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_59),
.B1(n_55),
.B2(n_57),
.Y(n_64)
);

XOR2x2_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_42),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_61),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_48),
.A2(n_44),
.B1(n_25),
.B2(n_26),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_50),
.B(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_66),
.Y(n_70)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_56),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_26),
.C(n_4),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

AO22x1_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_58),
.B1(n_63),
.B2(n_66),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_69),
.A2(n_71),
.B1(n_4),
.B2(n_7),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_63),
.A2(n_60),
.B(n_5),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_26),
.C(n_4),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_3),
.C(n_6),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_74),
.A2(n_68),
.B1(n_6),
.B2(n_2),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_76),
.C(n_77),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_26),
.C(n_3),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_26),
.C(n_3),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_79),
.A2(n_6),
.B1(n_7),
.B2(n_0),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_78),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_7),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_1),
.Y(n_83)
);


endmodule