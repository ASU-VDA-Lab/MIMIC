module fake_jpeg_21097_n_283 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_283);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_283;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_23),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_23),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_42),
.B(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_43),
.B(n_44),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_41),
.B(n_18),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_45),
.B(n_52),
.Y(n_90)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_28),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_19),
.B1(n_33),
.B2(n_16),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_54),
.B1(n_22),
.B2(n_32),
.Y(n_71)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_19),
.B1(n_33),
.B2(n_16),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_53),
.A2(n_32),
.B1(n_21),
.B2(n_30),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_19),
.B1(n_33),
.B2(n_16),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_63),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_18),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_64),
.B(n_21),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_65),
.Y(n_69)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_67),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_62),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_71),
.A2(n_87),
.B1(n_57),
.B2(n_61),
.Y(n_103)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_74),
.B(n_86),
.Y(n_92)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_78),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_46),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_80),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_27),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_21),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_83),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_44),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_82)
);

AO21x1_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_31),
.B(n_24),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_44),
.B(n_27),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_26),
.Y(n_86)
);

AOI211xp5_ASAP7_75t_SL g91 ( 
.A1(n_71),
.A2(n_50),
.B(n_39),
.C(n_34),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_91),
.A2(n_104),
.B(n_106),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_85),
.B(n_25),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_93),
.B(n_90),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_56),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_95),
.B(n_113),
.Y(n_133)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_64),
.B1(n_51),
.B2(n_55),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_109),
.B1(n_89),
.B2(n_75),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_103),
.A2(n_89),
.B1(n_75),
.B2(n_77),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_68),
.B(n_78),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_114),
.Y(n_128)
);

O2A1O1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_69),
.A2(n_47),
.B(n_48),
.C(n_52),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_82),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_111),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_66),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_84),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_88),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_88),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_84),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_116),
.B(n_122),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_102),
.Y(n_117)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_69),
.C(n_70),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_119),
.B(n_142),
.Y(n_165)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_131),
.Y(n_155)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_96),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_73),
.B(n_72),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_123),
.A2(n_134),
.B(n_135),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_108),
.B1(n_94),
.B2(n_32),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_130),
.A2(n_139),
.B1(n_109),
.B2(n_106),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_96),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_100),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_91),
.B(n_34),
.Y(n_135)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_92),
.B(n_2),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_140),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_34),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_138),
.A2(n_62),
.B(n_30),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_107),
.A2(n_84),
.B1(n_77),
.B2(n_21),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_99),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_97),
.B(n_34),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_105),
.B(n_113),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_143),
.A2(n_145),
.B(n_147),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_104),
.B(n_111),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_146),
.A2(n_153),
.B1(n_130),
.B2(n_141),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_111),
.B(n_114),
.Y(n_147)
);

AO22x1_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_97),
.B1(n_106),
.B2(n_115),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_SL g176 ( 
.A1(n_149),
.A2(n_157),
.B(n_138),
.C(n_139),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_92),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_158),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_102),
.B1(n_108),
.B2(n_93),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_156),
.B1(n_168),
.B2(n_138),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_123),
.A2(n_30),
.B1(n_94),
.B2(n_29),
.Y(n_156)
);

NAND2x1_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_94),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_29),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_167),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_128),
.A2(n_29),
.B(n_3),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_161),
.A2(n_4),
.B(n_6),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_118),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_162),
.B(n_125),
.Y(n_179)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_62),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_157),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_119),
.B(n_30),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_126),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_155),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_171),
.B(n_185),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_134),
.C(n_118),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_180),
.C(n_189),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_175),
.A2(n_176),
.B(n_151),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_167),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_151),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_178),
.A2(n_181),
.B1(n_191),
.B2(n_193),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_132),
.C(n_125),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_120),
.Y(n_182)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_184),
.Y(n_200)
);

NAND3xp33_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_4),
.C(n_7),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_127),
.Y(n_186)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_149),
.B(n_127),
.Y(n_187)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_144),
.Y(n_188)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_145),
.B(n_117),
.C(n_8),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_190),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_117),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_163),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_181),
.A2(n_143),
.B1(n_170),
.B2(n_147),
.Y(n_196)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_204),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_194),
.B(n_157),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_194),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_208),
.Y(n_227)
);

NAND2xp67_ASAP7_75t_SL g231 ( 
.A(n_206),
.B(n_9),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_172),
.Y(n_208)
);

A2O1A1O1Ixp25_ASAP7_75t_L g209 ( 
.A1(n_172),
.A2(n_161),
.B(n_166),
.C(n_153),
.D(n_158),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_209),
.B(n_189),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_180),
.B(n_169),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_215),
.C(n_192),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_191),
.A2(n_146),
.B1(n_163),
.B2(n_150),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_212),
.A2(n_216),
.B1(n_184),
.B2(n_186),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_175),
.A2(n_164),
.B(n_150),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_190),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_174),
.B(n_7),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_187),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_217),
.A2(n_218),
.B1(n_226),
.B2(n_220),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_197),
.A2(n_178),
.B1(n_174),
.B2(n_176),
.Y(n_219)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_215),
.Y(n_246)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_203),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_225),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_176),
.C(n_183),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_232),
.C(n_207),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_210),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_212),
.A2(n_176),
.B1(n_10),
.B2(n_11),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_230),
.Y(n_242)
);

BUFx12_ASAP7_75t_L g229 ( 
.A(n_198),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_213),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_199),
.B(n_9),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_231),
.A2(n_206),
.B(n_12),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_10),
.C(n_11),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_15),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_216),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_240),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_232),
.B(n_195),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_237),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_209),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_211),
.C(n_208),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_227),
.C(n_223),
.Y(n_247)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_243),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_11),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_245),
.A2(n_228),
.B1(n_204),
.B2(n_218),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_238),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_247),
.B(n_253),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_237),
.A2(n_224),
.B(n_233),
.Y(n_248)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_250),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_229),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_254),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_223),
.C(n_229),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_234),
.Y(n_254)
);

NOR2x1_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_246),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_R g259 ( 
.A(n_255),
.B(n_251),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_259),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_13),
.Y(n_273)
);

BUFx4f_ASAP7_75t_SL g263 ( 
.A(n_254),
.Y(n_263)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_263),
.Y(n_269)
);

AOI21x1_ASAP7_75t_L g264 ( 
.A1(n_256),
.A2(n_239),
.B(n_244),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_264),
.Y(n_267)
);

NOR2x1_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_241),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_247),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_261),
.B(n_257),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_270),
.C(n_271),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_261),
.B(n_253),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_262),
.C(n_258),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_267),
.A2(n_262),
.B1(n_265),
.B2(n_263),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_274),
.Y(n_280)
);

AOI322xp5_ASAP7_75t_L g279 ( 
.A1(n_276),
.A2(n_277),
.A3(n_278),
.B1(n_14),
.B2(n_272),
.C1(n_273),
.C2(n_275),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_15),
.C(n_13),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_269),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_279),
.Y(n_281)
);

NOR3xp33_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_280),
.C(n_14),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_14),
.Y(n_283)
);


endmodule