module real_aes_15724_n_4 (n_0, n_3, n_2, n_1, n_4);
input n_0;
input n_3;
input n_2;
input n_1;
output n_4;
wire n_17;
wire n_22;
wire n_24;
wire n_13;
wire n_6;
wire n_12;
wire n_19;
wire n_25;
wire n_14;
wire n_11;
wire n_16;
wire n_5;
wire n_15;
wire n_9;
wire n_23;
wire n_20;
wire n_26;
wire n_18;
wire n_21;
wire n_7;
wire n_8;
wire n_10;
HB1xp67_ASAP7_75t_L g7 ( .A(n_0), .Y(n_7) );
AND2x4_ASAP7_75t_L g17 ( .A(n_0), .B(n_9), .Y(n_17) );
INVx2_ASAP7_75t_L g13 ( .A(n_1), .Y(n_13) );
INVx1_ASAP7_75t_L g9 ( .A(n_2), .Y(n_9) );
BUFx6f_ASAP7_75t_L g23 ( .A(n_3), .Y(n_23) );
AOI211xp5_ASAP7_75t_L g4 ( .A1(n_5), .A2(n_10), .B(n_14), .C(n_24), .Y(n_4) );
AND2x2_ASAP7_75t_L g5 ( .A(n_6), .B(n_8), .Y(n_5) );
INVx1_ASAP7_75t_L g6 ( .A(n_7), .Y(n_6) );
HB1xp67_ASAP7_75t_L g8 ( .A(n_9), .Y(n_8) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_10), .B(n_19), .Y(n_18) );
HB1xp67_ASAP7_75t_L g10 ( .A(n_11), .Y(n_10) );
INVx6_ASAP7_75t_L g11 ( .A(n_12), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_12), .B(n_26), .Y(n_25) );
BUFx8_ASAP7_75t_L g12 ( .A(n_13), .Y(n_12) );
NOR2xp33_ASAP7_75t_L g14 ( .A(n_15), .B(n_18), .Y(n_14) );
NOR2xp33_ASAP7_75t_L g24 ( .A(n_15), .B(n_25), .Y(n_24) );
INVx2_ASAP7_75t_L g15 ( .A(n_16), .Y(n_15) );
BUFx10_ASAP7_75t_L g16 ( .A(n_17), .Y(n_16) );
INVx1_ASAP7_75t_L g26 ( .A(n_19), .Y(n_26) );
HB1xp67_ASAP7_75t_L g19 ( .A(n_20), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_21), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_22), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_23), .Y(n_22) );
endmodule