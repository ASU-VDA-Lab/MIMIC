module fake_jpeg_8108_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_10),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

AND2x2_ASAP7_75t_SL g45 ( 
.A(n_16),
.B(n_0),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_34),
.C(n_20),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_26),
.B(n_7),
.Y(n_46)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_30),
.Y(n_47)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_29),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_51),
.B(n_63),
.Y(n_101)
);

NAND2xp33_ASAP7_75t_SL g55 ( 
.A(n_45),
.B(n_0),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_55),
.A2(n_34),
.B1(n_44),
.B2(n_37),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_59),
.B(n_39),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_29),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_29),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_36),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_22),
.B1(n_35),
.B2(n_19),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_65),
.A2(n_54),
.B1(n_20),
.B2(n_21),
.Y(n_74)
);

CKINVDCx12_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_26),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_34),
.C(n_20),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_18),
.Y(n_70)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_40),
.A2(n_22),
.B1(n_19),
.B2(n_28),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_24),
.B1(n_33),
.B2(n_32),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_73),
.B(n_108),
.C(n_31),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_74),
.B(n_102),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_75),
.B(n_106),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_21),
.B1(n_22),
.B2(n_44),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_51),
.A2(n_41),
.B1(n_39),
.B2(n_21),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_77),
.A2(n_83),
.B1(n_97),
.B2(n_27),
.Y(n_129)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_79),
.B(n_86),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_41),
.B1(n_28),
.B2(n_18),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_82),
.A2(n_104),
.B1(n_60),
.B2(n_17),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_64),
.B(n_24),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_85),
.B(n_98),
.Y(n_113)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_48),
.A2(n_44),
.B1(n_36),
.B2(n_37),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_65),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_91),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_67),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVxp33_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_59),
.A2(n_41),
.B1(n_42),
.B2(n_37),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_94),
.A2(n_99),
.B1(n_105),
.B2(n_39),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_53),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_100),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_96),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_71),
.A2(n_44),
.B1(n_36),
.B2(n_37),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_53),
.B(n_33),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_55),
.A2(n_42),
.B1(n_39),
.B2(n_36),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_52),
.A2(n_41),
.B1(n_27),
.B2(n_32),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_62),
.A2(n_42),
.B1(n_39),
.B2(n_17),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_109),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_38),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_57),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_110),
.B(n_58),
.Y(n_128)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_90),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_121),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_116),
.A2(n_120),
.B1(n_137),
.B2(n_92),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_89),
.A2(n_39),
.B1(n_58),
.B2(n_60),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_124),
.Y(n_152)
);

BUFx24_ASAP7_75t_SL g124 ( 
.A(n_78),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_126),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_90),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_128),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_129),
.A2(n_134),
.B1(n_88),
.B2(n_103),
.Y(n_161)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_139),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_43),
.C(n_38),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_137),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_102),
.A2(n_38),
.B1(n_43),
.B2(n_17),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_73),
.Y(n_148)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_90),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_111),
.Y(n_165)
);

OR2x4_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_75),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_142),
.A2(n_156),
.B(n_164),
.Y(n_196)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_140),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_143),
.B(n_144),
.Y(n_188)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_140),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_112),
.A2(n_99),
.B(n_106),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_145),
.A2(n_157),
.B(n_160),
.Y(n_181)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_146),
.B(n_149),
.Y(n_192)
);

OAI21xp33_ASAP7_75t_SL g204 ( 
.A1(n_147),
.A2(n_38),
.B(n_126),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_148),
.B(n_43),
.Y(n_195)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_138),
.C(n_132),
.Y(n_186)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_153),
.B(n_159),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_101),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_155),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_101),
.Y(n_155)
);

AND2x2_ASAP7_75t_SL g156 ( 
.A(n_123),
.B(n_88),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

INVxp33_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_119),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_161),
.A2(n_163),
.B1(n_174),
.B2(n_139),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_74),
.B1(n_85),
.B2(n_100),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_127),
.A2(n_78),
.B(n_80),
.Y(n_164)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_169),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_84),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_167),
.B(n_143),
.Y(n_187)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_121),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_118),
.B(n_80),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_171),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_118),
.B(n_83),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_117),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_173),
.Y(n_203)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_117),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_116),
.A2(n_96),
.B1(n_103),
.B2(n_109),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_127),
.B(n_84),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_43),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_176),
.A2(n_197),
.B1(n_204),
.B2(n_107),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_166),
.A2(n_131),
.B1(n_127),
.B2(n_129),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_177),
.A2(n_190),
.B1(n_164),
.B2(n_163),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_158),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_178),
.B(n_179),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_150),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_SL g180 ( 
.A1(n_142),
.A2(n_145),
.B(n_162),
.C(n_147),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_180),
.A2(n_199),
.B(n_31),
.Y(n_232)
);

XNOR2x2_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_136),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_182),
.A2(n_185),
.B(n_189),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_169),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_187),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_157),
.A2(n_133),
.B1(n_134),
.B2(n_136),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_191),
.C(n_195),
.Y(n_213)
);

AND2x2_ASAP7_75t_SL g189 ( 
.A(n_146),
.B(n_149),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_174),
.A2(n_113),
.B1(n_125),
.B2(n_132),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_113),
.Y(n_191)
);

CKINVDCx12_ASAP7_75t_R g193 ( 
.A(n_170),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_208),
.Y(n_219)
);

AO21x2_ASAP7_75t_L g197 ( 
.A1(n_153),
.A2(n_103),
.B(n_38),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_151),
.B(n_0),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_200),
.A2(n_201),
.B1(n_205),
.B2(n_114),
.Y(n_233)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_173),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_156),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_207),
.B(n_144),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_156),
.Y(n_208)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_209),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_206),
.B(n_168),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_211),
.B(n_214),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_212),
.A2(n_234),
.B1(n_205),
.B2(n_185),
.Y(n_238)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_203),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_206),
.B(n_171),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_215),
.B(n_217),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_186),
.C(n_182),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_216),
.B(n_199),
.C(n_25),
.Y(n_259)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_226),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_155),
.Y(n_221)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_153),
.Y(n_222)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_154),
.C(n_156),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_231),
.C(n_207),
.Y(n_244)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_188),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_224),
.B(n_227),
.Y(n_256)
);

BUFx24_ASAP7_75t_SL g226 ( 
.A(n_194),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_141),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_183),
.B(n_160),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_229),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_189),
.Y(n_229)
);

OAI21xp33_ASAP7_75t_L g230 ( 
.A1(n_208),
.A2(n_152),
.B(n_13),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_11),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_43),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_236),
.Y(n_254)
);

OA22x2_ASAP7_75t_L g246 ( 
.A1(n_233),
.A2(n_197),
.B1(n_181),
.B2(n_180),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_196),
.A2(n_26),
.B(n_25),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_235),
.A2(n_197),
.B(n_200),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_189),
.B(n_26),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_234),
.A2(n_190),
.B1(n_202),
.B2(n_177),
.Y(n_237)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_238),
.A2(n_215),
.B1(n_224),
.B2(n_217),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_210),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_239),
.B(n_240),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_218),
.A2(n_176),
.B1(n_180),
.B2(n_181),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_243),
.A2(n_258),
.B1(n_236),
.B2(n_209),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_248),
.C(n_255),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_246),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_180),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_228),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_213),
.B(n_223),
.C(n_220),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_249),
.B(n_235),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_253),
.B(n_9),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_213),
.B(n_220),
.C(n_231),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_229),
.A2(n_197),
.B1(n_201),
.B2(n_199),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_25),
.C(n_17),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_212),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_263),
.C(n_274),
.Y(n_283)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_261),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_214),
.Y(n_262)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_262),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_232),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_268),
.Y(n_289)
);

INVxp33_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_271),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_240),
.A2(n_219),
.B(n_211),
.Y(n_268)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_275),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_267),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_221),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_277),
.C(n_259),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_81),
.C(n_2),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_251),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_239),
.Y(n_290)
);

XNOR2x1_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_246),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_280),
.A2(n_254),
.B(n_253),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_263),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_266),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_265),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_284),
.B(n_285),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_271),
.B(n_241),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_260),
.C(n_274),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_288),
.C(n_276),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_252),
.C(n_258),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_290),
.B(n_292),
.Y(n_307)
);

A2O1A1Ixp33_ASAP7_75t_SL g291 ( 
.A1(n_269),
.A2(n_246),
.B(n_242),
.C(n_243),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_291),
.A2(n_246),
.B(n_264),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_270),
.B(n_245),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_298),
.C(n_303),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_297),
.Y(n_313)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_280),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_6),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_300),
.B(n_301),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_279),
.A2(n_254),
.B1(n_81),
.B2(n_3),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_304),
.B1(n_6),
.B2(n_9),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_293),
.C(n_289),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_293),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_8),
.C(n_13),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_1),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_287),
.A2(n_7),
.B(n_12),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_306),
.A2(n_7),
.B(n_15),
.Y(n_310)
);

AOI21x1_ASAP7_75t_SL g308 ( 
.A1(n_300),
.A2(n_291),
.B(n_282),
.Y(n_308)
);

AOI322xp5_ASAP7_75t_L g318 ( 
.A1(n_308),
.A2(n_311),
.A3(n_296),
.B1(n_295),
.B2(n_298),
.C1(n_305),
.C2(n_11),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_2),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_291),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_316),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_315),
.A2(n_317),
.B1(n_15),
.B2(n_4),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_11),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_299),
.A2(n_304),
.B1(n_307),
.B2(n_302),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_320),
.C(n_309),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_321),
.Y(n_325)
);

AOI32xp33_ASAP7_75t_SL g320 ( 
.A1(n_309),
.A2(n_2),
.A3(n_4),
.B1(n_5),
.B2(n_9),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_311),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_323),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_5),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_327),
.A2(n_325),
.B(n_326),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_328),
.A2(n_322),
.B(n_320),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_329),
.B(n_330),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_327),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_312),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_5),
.Y(n_334)
);


endmodule