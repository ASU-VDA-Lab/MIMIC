module fake_jpeg_1337_n_213 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_213);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_213;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_27),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_14),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_12),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_33),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_22),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_14),
.Y(n_64)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_6),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_28),
.B(n_3),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_74),
.Y(n_89)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

BUFx4f_ASAP7_75t_SL g85 ( 
.A(n_75),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_81),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_74),
.A2(n_61),
.B1(n_72),
.B2(n_70),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_83),
.A2(n_87),
.B1(n_85),
.B2(n_75),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_63),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_91),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_61),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g110 ( 
.A(n_86),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_56),
.B1(n_57),
.B2(n_52),
.Y(n_87)
);

NAND2x1p5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_71),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_75),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_64),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_69),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_92),
.B(n_94),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_67),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_91),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_96),
.B(n_105),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_86),
.A2(n_50),
.B1(n_54),
.B2(n_60),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_106),
.B1(n_89),
.B2(n_95),
.Y(n_115)
);

INVxp33_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_57),
.B1(n_52),
.B2(n_51),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_101),
.A2(n_84),
.B1(n_93),
.B2(n_94),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_50),
.C(n_54),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_65),
.Y(n_131)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

BUFx2_ASAP7_75t_SL g104 ( 
.A(n_85),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

AOI21xp33_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_73),
.B(n_55),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_82),
.A2(n_65),
.B1(n_53),
.B2(n_55),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_65),
.B(n_58),
.C(n_90),
.Y(n_132)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_113),
.Y(n_127)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_112),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_92),
.B(n_62),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_131),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_88),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_119),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_108),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_120),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_108),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_124),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_88),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_103),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_133),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_95),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_129),
.B(n_0),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_98),
.A2(n_101),
.B1(n_107),
.B2(n_109),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_130),
.A2(n_51),
.B1(n_58),
.B2(n_66),
.Y(n_141)
);

NOR3xp33_ASAP7_75t_SL g150 ( 
.A(n_132),
.B(n_1),
.C(n_2),
.Y(n_150)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_90),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_134),
.B(n_100),
.Y(n_139)
);

INVxp33_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_138),
.Y(n_163)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_9),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_8),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_150),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_124),
.A2(n_72),
.B1(n_70),
.B2(n_66),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_154),
.B1(n_155),
.B2(n_157),
.Y(n_164)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_146),
.B(n_149),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_72),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_158),
.C(n_125),
.Y(n_162)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_151),
.B(n_152),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_123),
.B(n_122),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_121),
.A2(n_1),
.B(n_2),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_153),
.A2(n_6),
.B(n_7),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_48),
.B1(n_46),
.B2(n_45),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_116),
.A2(n_44),
.B1(n_42),
.B2(n_41),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_38),
.C(n_37),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_147),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_160),
.B(n_162),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_156),
.A2(n_120),
.B1(n_115),
.B2(n_131),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_161),
.A2(n_135),
.B1(n_155),
.B2(n_142),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_132),
.B1(n_125),
.B2(n_8),
.Y(n_165)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

AOI21xp33_ASAP7_75t_L g183 ( 
.A1(n_168),
.A2(n_174),
.B(n_176),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_35),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_171),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_34),
.C(n_32),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_173),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_31),
.C(n_30),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_157),
.Y(n_177)
);

AOI322xp5_ASAP7_75t_L g182 ( 
.A1(n_177),
.A2(n_10),
.A3(n_15),
.B1(n_16),
.B2(n_17),
.C1(n_18),
.C2(n_19),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_180),
.B(n_182),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_161),
.A2(n_150),
.B1(n_11),
.B2(n_13),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_181),
.A2(n_185),
.B1(n_188),
.B2(n_168),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_159),
.A2(n_29),
.B(n_26),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_175),
.Y(n_186)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_186),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_167),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_162),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_193),
.C(n_194),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_192),
.A2(n_195),
.B1(n_164),
.B2(n_187),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_169),
.C(n_178),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_163),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_186),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_179),
.A2(n_167),
.B1(n_173),
.B2(n_166),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_197),
.A2(n_179),
.B1(n_188),
.B2(n_181),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_198),
.B(n_200),
.Y(n_204)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_194),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_199),
.A2(n_202),
.B1(n_197),
.B2(n_193),
.Y(n_205)
);

NOR3xp33_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_167),
.C(n_185),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_190),
.C(n_172),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_176),
.C(n_183),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_205),
.A2(n_191),
.B1(n_200),
.B2(n_189),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_206),
.A2(n_207),
.B1(n_204),
.B2(n_19),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_18),
.C(n_21),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_23),
.C(n_24),
.Y(n_210)
);

INVxp33_ASAP7_75t_L g211 ( 
.A(n_210),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_211),
.A2(n_23),
.B(n_25),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_25),
.Y(n_213)
);


endmodule