module fake_aes_5641_n_291 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_93, n_51, n_96, n_39, n_291);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_93;
input n_51;
input n_96;
input n_39;
output n_291;
wire n_117;
wire n_219;
wire n_133;
wire n_149;
wire n_289;
wire n_220;
wire n_214;
wire n_267;
wire n_204;
wire n_221;
wire n_249;
wire n_185;
wire n_203;
wire n_244;
wire n_102;
wire n_119;
wire n_141;
wire n_115;
wire n_167;
wire n_284;
wire n_107;
wire n_158;
wire n_278;
wire n_114;
wire n_121;
wire n_171;
wire n_196;
wire n_125;
wire n_192;
wire n_240;
wire n_254;
wire n_161;
wire n_262;
wire n_177;
wire n_130;
wire n_189;
wire n_103;
wire n_239;
wire n_137;
wire n_180;
wire n_104;
wire n_277;
wire n_160;
wire n_276;
wire n_154;
wire n_272;
wire n_285;
wire n_195;
wire n_165;
wire n_146;
wire n_250;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_215;
wire n_155;
wire n_108;
wire n_116;
wire n_229;
wire n_209;
wire n_217;
wire n_139;
wire n_230;
wire n_274;
wire n_198;
wire n_169;
wire n_193;
wire n_273;
wire n_282;
wire n_252;
wire n_152;
wire n_113;
wire n_241;
wire n_124;
wire n_156;
wire n_238;
wire n_128;
wire n_120;
wire n_129;
wire n_206;
wire n_245;
wire n_135;
wire n_188;
wire n_260;
wire n_201;
wire n_197;
wire n_242;
wire n_247;
wire n_127;
wire n_170;
wire n_111;
wire n_157;
wire n_202;
wire n_210;
wire n_142;
wire n_184;
wire n_265;
wire n_191;
wire n_264;
wire n_281;
wire n_232;
wire n_200;
wire n_208;
wire n_211;
wire n_122;
wire n_187;
wire n_138;
wire n_126;
wire n_275;
wire n_178;
wire n_118;
wire n_258;
wire n_253;
wire n_179;
wire n_131;
wire n_112;
wire n_266;
wire n_205;
wire n_213;
wire n_143;
wire n_235;
wire n_243;
wire n_182;
wire n_263;
wire n_166;
wire n_186;
wire n_162;
wire n_163;
wire n_226;
wire n_105;
wire n_227;
wire n_174;
wire n_159;
wire n_248;
wire n_268;
wire n_231;
wire n_136;
wire n_283;
wire n_176;
wire n_144;
wire n_183;
wire n_256;
wire n_216;
wire n_147;
wire n_199;
wire n_148;
wire n_123;
wire n_172;
wire n_100;
wire n_212;
wire n_228;
wire n_223;
wire n_251;
wire n_236;
wire n_150;
wire n_218;
wire n_168;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_134;
wire n_222;
wire n_234;
wire n_164;
wire n_233;
wire n_271;
wire n_106;
wire n_175;
wire n_173;
wire n_190;
wire n_286;
wire n_145;
wire n_270;
wire n_246;
wire n_153;
wire n_259;
wire n_290;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_288;
wire n_151;
wire n_140;
wire n_207;
wire n_257;
wire n_224;
wire n_269;
wire n_225;
wire n_279;
INVx1_ASAP7_75t_L g99 ( .A(n_95), .Y(n_99) );
INVxp67_ASAP7_75t_L g100 ( .A(n_74), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_5), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_53), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_80), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_67), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_51), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_60), .Y(n_106) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_54), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_86), .Y(n_108) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_46), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_19), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_92), .Y(n_111) );
BUFx3_ASAP7_75t_L g112 ( .A(n_30), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_66), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_71), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_24), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_69), .B(n_90), .Y(n_116) );
BUFx3_ASAP7_75t_L g117 ( .A(n_40), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_17), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_32), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_96), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_29), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_27), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_47), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_88), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_70), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_31), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_83), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_3), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_41), .Y(n_129) );
INVx2_ASAP7_75t_SL g130 ( .A(n_91), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_37), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_36), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_93), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_78), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_87), .Y(n_135) );
CKINVDCx16_ASAP7_75t_R g136 ( .A(n_77), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_1), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_34), .Y(n_138) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_75), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_79), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_33), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_39), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_89), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_14), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_3), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_55), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_28), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_18), .Y(n_148) );
INVxp67_ASAP7_75t_SL g149 ( .A(n_81), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_11), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_43), .Y(n_151) );
INVxp67_ASAP7_75t_SL g152 ( .A(n_35), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_15), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_82), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_1), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_73), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_42), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_20), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_72), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_85), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_94), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_13), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_26), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_68), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_38), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_76), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_84), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_111), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_139), .Y(n_169) );
NOR2xp33_ASAP7_75t_SL g170 ( .A(n_107), .B(n_6), .Y(n_170) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_101), .Y(n_171) );
CKINVDCx16_ASAP7_75t_R g172 ( .A(n_136), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_130), .B(n_0), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_109), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_145), .Y(n_175) );
AND2x4_ASAP7_75t_L g176 ( .A(n_128), .B(n_2), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_137), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_109), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_155), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_132), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_99), .Y(n_181) );
OAI22x1_ASAP7_75t_L g182 ( .A1(n_168), .A2(n_152), .B1(n_149), .B2(n_102), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_176), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_180), .Y(n_184) );
INVx4_ASAP7_75t_L g185 ( .A(n_172), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_181), .Y(n_186) );
NOR2x1p5_ASAP7_75t_L g187 ( .A(n_169), .B(n_103), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_171), .B(n_100), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_186), .B(n_177), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_187), .A2(n_179), .B1(n_173), .B2(n_170), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_184), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_186), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_188), .B(n_175), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_183), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_183), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_187), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_196), .B(n_185), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_192), .A2(n_122), .B1(n_125), .B2(n_114), .Y(n_198) );
OAI21xp33_ASAP7_75t_L g199 ( .A1(n_194), .A2(n_182), .B(n_113), .Y(n_199) );
OAI21xp33_ASAP7_75t_L g200 ( .A1(n_195), .A2(n_118), .B(n_108), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_189), .A2(n_116), .B(n_104), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_190), .B(n_119), .Y(n_202) );
BUFx2_ASAP7_75t_SL g203 ( .A(n_193), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_191), .Y(n_204) );
AOI221x1_ASAP7_75t_L g205 ( .A1(n_199), .A2(n_141), .B1(n_105), .B2(n_106), .C(n_110), .Y(n_205) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_201), .A2(n_115), .B(n_121), .C(n_120), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_202), .A2(n_126), .B(n_124), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_204), .Y(n_208) );
AO31x2_ASAP7_75t_L g209 ( .A1(n_197), .A2(n_150), .A3(n_127), .B(n_129), .Y(n_209) );
OR2x2_ASAP7_75t_L g210 ( .A(n_198), .B(n_4), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_200), .A2(n_133), .B(n_131), .Y(n_211) );
INVxp67_ASAP7_75t_L g212 ( .A(n_198), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_203), .B(n_135), .Y(n_213) );
OAI21x1_ASAP7_75t_SL g214 ( .A1(n_201), .A2(n_140), .B(n_138), .Y(n_214) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_204), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_215), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_213), .B(n_123), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_210), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_209), .Y(n_219) );
AOI21x1_ASAP7_75t_L g220 ( .A1(n_214), .A2(n_144), .B(n_142), .Y(n_220) );
OA21x2_ASAP7_75t_L g221 ( .A1(n_205), .A2(n_147), .B(n_146), .Y(n_221) );
AO22x2_ASAP7_75t_L g222 ( .A1(n_207), .A2(n_167), .B1(n_148), .B2(n_165), .Y(n_222) );
AO31x2_ASAP7_75t_L g223 ( .A1(n_211), .A2(n_160), .A3(n_151), .B(n_153), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_208), .Y(n_224) );
AO31x2_ASAP7_75t_L g225 ( .A1(n_205), .A2(n_162), .A3(n_154), .B(n_156), .Y(n_225) );
OAI21xp5_ASAP7_75t_L g226 ( .A1(n_206), .A2(n_161), .B(n_158), .Y(n_226) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_215), .Y(n_227) );
INVx6_ASAP7_75t_L g228 ( .A(n_215), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_212), .A2(n_112), .B1(n_117), .B2(n_134), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_224), .Y(n_230) );
INVx2_ASAP7_75t_SL g231 ( .A(n_228), .Y(n_231) );
INVx3_ASAP7_75t_L g232 ( .A(n_216), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_227), .Y(n_233) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_220), .A2(n_178), .B(n_174), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_223), .Y(n_235) );
INVx2_ASAP7_75t_SL g236 ( .A(n_217), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_222), .B(n_157), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_225), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_221), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_226), .B(n_159), .Y(n_240) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_229), .A2(n_166), .B(n_164), .Y(n_241) );
AND2x4_ASAP7_75t_L g242 ( .A(n_216), .B(n_143), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_218), .B(n_163), .Y(n_243) );
OA21x2_ASAP7_75t_L g244 ( .A1(n_219), .A2(n_7), .B(n_8), .Y(n_244) );
INVx3_ASAP7_75t_L g245 ( .A(n_216), .Y(n_245) );
AO21x2_ASAP7_75t_L g246 ( .A1(n_219), .A2(n_9), .B(n_10), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_230), .B(n_12), .Y(n_247) );
BUFx2_ASAP7_75t_L g248 ( .A(n_232), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_237), .B(n_16), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_238), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_233), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_231), .B(n_21), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_245), .B(n_22), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_242), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_238), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_236), .B(n_98), .Y(n_256) );
INVxp67_ASAP7_75t_SL g257 ( .A(n_239), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_235), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_243), .B(n_23), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_251), .B(n_246), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_248), .B(n_241), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_250), .B(n_234), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_250), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_255), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_255), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_249), .B(n_244), .Y(n_266) );
OR2x2_ASAP7_75t_L g267 ( .A(n_257), .B(n_240), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_254), .B(n_25), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_258), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_263), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_264), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_265), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_269), .Y(n_273) );
OR2x2_ASAP7_75t_L g274 ( .A(n_273), .B(n_267), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_270), .Y(n_275) );
OAI221xp5_ASAP7_75t_SL g276 ( .A1(n_274), .A2(n_266), .B1(n_261), .B2(n_272), .C(n_271), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_275), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_275), .Y(n_278) );
AOI221xp5_ASAP7_75t_L g279 ( .A1(n_276), .A2(n_256), .B1(n_259), .B2(n_262), .C(n_260), .Y(n_279) );
NOR4xp25_ASAP7_75t_L g280 ( .A(n_277), .B(n_268), .C(n_247), .D(n_252), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_278), .B(n_253), .Y(n_281) );
NAND3xp33_ASAP7_75t_L g282 ( .A(n_279), .B(n_280), .C(n_281), .Y(n_282) );
NOR2x1_ASAP7_75t_L g283 ( .A(n_282), .B(n_44), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_283), .B(n_97), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_284), .Y(n_285) );
OAI22xp5_ASAP7_75t_SL g286 ( .A1(n_285), .A2(n_45), .B1(n_48), .B2(n_49), .Y(n_286) );
AND2x4_ASAP7_75t_L g287 ( .A(n_286), .B(n_50), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_287), .A2(n_52), .B1(n_56), .B2(n_57), .Y(n_288) );
NAND2x1p5_ASAP7_75t_L g289 ( .A(n_288), .B(n_58), .Y(n_289) );
XNOR2xp5_ASAP7_75t_L g290 ( .A(n_289), .B(n_59), .Y(n_290) );
AOI222xp33_ASAP7_75t_L g291 ( .A1(n_290), .A2(n_61), .B1(n_62), .B2(n_63), .C1(n_64), .C2(n_65), .Y(n_291) );
endmodule