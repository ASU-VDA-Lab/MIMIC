module fake_jpeg_24492_n_343 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_0),
.B(n_5),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_8),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

CKINVDCx6p67_ASAP7_75t_R g70 ( 
.A(n_40),
.Y(n_70)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_44),
.Y(n_58)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_8),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_37),
.B(n_18),
.C(n_23),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_32),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_47),
.A2(n_19),
.B1(n_17),
.B2(n_31),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_19),
.B1(n_25),
.B2(n_29),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_51),
.A2(n_64),
.B1(n_42),
.B2(n_26),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_52),
.Y(n_88)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_55),
.B(n_61),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_56),
.A2(n_17),
.B1(n_31),
.B2(n_27),
.Y(n_94)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_62),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_46),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_18),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_25),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_69),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_36),
.B1(n_34),
.B2(n_19),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_27),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_72),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_69),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_76),
.Y(n_115)
);

AO22x1_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_47),
.B1(n_48),
.B2(n_38),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_75),
.A2(n_101),
.B(n_39),
.Y(n_122)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_61),
.B(n_34),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_L g111 ( 
.A1(n_77),
.A2(n_84),
.B(n_85),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_79),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_86),
.Y(n_116)
);

NOR2x1_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_34),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_82),
.A2(n_94),
.B1(n_17),
.B2(n_31),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_36),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_52),
.B(n_36),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_70),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_90),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_89),
.A2(n_59),
.B1(n_60),
.B2(n_50),
.Y(n_105)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_52),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_92),
.B(n_93),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_29),
.B(n_23),
.C(n_26),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_70),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_97),
.A2(n_98),
.B1(n_59),
.B2(n_49),
.Y(n_108)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

OA22x2_ASAP7_75t_SL g101 ( 
.A1(n_54),
.A2(n_48),
.B1(n_38),
.B2(n_40),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_80),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_104),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_53),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_105),
.A2(n_122),
.B1(n_126),
.B2(n_97),
.Y(n_158)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_113),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_80),
.B1(n_71),
.B2(n_82),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_119),
.B1(n_121),
.B2(n_123),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_75),
.A2(n_49),
.B1(n_59),
.B2(n_65),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_86),
.B(n_96),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_79),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_117),
.B(n_120),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_130),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_67),
.B1(n_57),
.B2(n_50),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_84),
.A2(n_26),
.B1(n_30),
.B2(n_33),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_101),
.A2(n_66),
.B1(n_30),
.B2(n_33),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_73),
.A2(n_66),
.B1(n_30),
.B2(n_33),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_91),
.B1(n_95),
.B2(n_83),
.Y(n_159)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_128),
.B(n_55),
.Y(n_154)
);

INVxp33_ASAP7_75t_SL g129 ( 
.A(n_101),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_126),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_131),
.A2(n_142),
.B(n_117),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_129),
.A2(n_128),
.B1(n_120),
.B2(n_121),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_151),
.B1(n_159),
.B2(n_110),
.Y(n_163)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_139),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_80),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_137),
.B(n_149),
.Y(n_189)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_138),
.B(n_145),
.Y(n_194)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_147),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_77),
.B(n_78),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_143),
.Y(n_185)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_152),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_104),
.B(n_77),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_103),
.B(n_125),
.Y(n_150)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_122),
.A2(n_78),
.B1(n_90),
.B2(n_87),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_103),
.B(n_85),
.Y(n_153)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_154),
.A2(n_158),
.B1(n_123),
.B2(n_109),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_112),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_155),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_98),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_156),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_108),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_79),
.Y(n_181)
);

AO22x1_ASAP7_75t_L g169 ( 
.A1(n_160),
.A2(n_127),
.B1(n_105),
.B2(n_48),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_116),
.B(n_85),
.Y(n_161)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_163),
.A2(n_179),
.B1(n_181),
.B2(n_153),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_164),
.B(n_175),
.Y(n_211)
);

NAND2x1_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_111),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_L g218 ( 
.A1(n_165),
.A2(n_169),
.B(n_173),
.Y(n_218)
);

AND2x6_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_112),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_172),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_R g170 ( 
.A(n_142),
.B(n_21),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_170),
.B(n_135),
.Y(n_198)
);

INVx3_ASAP7_75t_SL g172 ( 
.A(n_143),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_83),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_193),
.C(n_144),
.Y(n_195)
);

NOR2x1_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_107),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_132),
.A2(n_107),
.B1(n_95),
.B2(n_74),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_131),
.A2(n_74),
.B(n_88),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_91),
.Y(n_182)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_24),
.Y(n_184)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_184),
.Y(n_203)
);

INVx13_ASAP7_75t_L g186 ( 
.A(n_143),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_187),
.Y(n_210)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

AO22x2_ASAP7_75t_L g188 ( 
.A1(n_160),
.A2(n_33),
.B1(n_26),
.B2(n_40),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_188),
.A2(n_159),
.B1(n_157),
.B2(n_146),
.Y(n_196)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_134),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_3),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_139),
.B(n_24),
.Y(n_191)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_152),
.B(n_28),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_192),
.B(n_21),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_133),
.B(n_24),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_212),
.C(n_214),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_196),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_242)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_199),
.B(n_209),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_163),
.A2(n_146),
.B1(n_151),
.B2(n_141),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_200),
.A2(n_201),
.B1(n_207),
.B2(n_208),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_167),
.B(n_133),
.Y(n_206)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_206),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_179),
.A2(n_160),
.B1(n_148),
.B2(n_147),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_166),
.A2(n_132),
.B1(n_138),
.B2(n_145),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_168),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_136),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_24),
.Y(n_213)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_213),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_28),
.C(n_24),
.Y(n_214)
);

OAI22x1_ASAP7_75t_L g215 ( 
.A1(n_188),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_188),
.A2(n_20),
.B1(n_3),
.B2(n_2),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_188),
.A2(n_20),
.B1(n_3),
.B2(n_2),
.Y(n_217)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_220),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_4),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_165),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_171),
.B(n_4),
.Y(n_222)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_222),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_4),
.C(n_5),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_192),
.C(n_9),
.Y(n_250)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_162),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_224),
.B(n_190),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_210),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_234),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_185),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_227),
.B(n_216),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_205),
.A2(n_173),
.B(n_180),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_228),
.A2(n_229),
.B1(n_245),
.B2(n_217),
.Y(n_271)
);

OA22x2_ASAP7_75t_L g229 ( 
.A1(n_215),
.A2(n_175),
.B1(n_169),
.B2(n_176),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_233),
.C(n_238),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_195),
.C(n_165),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_197),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_236),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_207),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_177),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_239),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_178),
.C(n_183),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_178),
.C(n_183),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_200),
.B(n_167),
.C(n_194),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_244),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_202),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_243),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_170),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_205),
.A2(n_176),
.B(n_169),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_250),
.B(n_223),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_238),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_248),
.B(n_218),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_253),
.B(n_258),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_226),
.Y(n_257)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_257),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_248),
.B(n_196),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_221),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_231),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_211),
.Y(n_261)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_251),
.Y(n_262)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_262),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_186),
.Y(n_263)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_185),
.Y(n_264)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_264),
.Y(n_285)
);

INVxp67_ASAP7_75t_SL g265 ( 
.A(n_246),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_265),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_241),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_267),
.Y(n_289)
);

MAJx2_ASAP7_75t_L g269 ( 
.A(n_225),
.B(n_203),
.C(n_204),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_269),
.B(n_271),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_237),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_272),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_233),
.B(n_172),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_239),
.C(n_228),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_232),
.Y(n_274)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_274),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_276),
.B(n_279),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_280),
.C(n_282),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_230),
.C(n_245),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_235),
.C(n_242),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_255),
.B(n_247),
.C(n_250),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_256),
.C(n_268),
.Y(n_300)
);

NOR3xp33_ASAP7_75t_SL g291 ( 
.A(n_289),
.B(n_269),
.C(n_261),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_295),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_282),
.A2(n_285),
.B(n_284),
.Y(n_292)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_292),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_266),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_293),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_286),
.B(n_253),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_268),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_187),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_274),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_296),
.A2(n_304),
.B(n_290),
.Y(n_318)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_287),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_302),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_277),
.C(n_280),
.Y(n_308)
);

OAI21x1_ASAP7_75t_L g301 ( 
.A1(n_287),
.A2(n_265),
.B(n_263),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_286),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_283),
.B(n_249),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_275),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_303),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_278),
.A2(n_254),
.B(n_258),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_229),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_294),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_308),
.C(n_314),
.Y(n_322)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_312),
.Y(n_321)
);

INVx6_ASAP7_75t_L g313 ( 
.A(n_291),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_313),
.A2(n_318),
.B1(n_16),
.B2(n_11),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_296),
.B(n_276),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_229),
.Y(n_317)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_317),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_319),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_305),
.Y(n_320)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_320),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_316),
.B(n_298),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_309),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_300),
.C(n_172),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_324),
.A2(n_327),
.B(n_312),
.Y(n_335)
);

AOI322xp5_ASAP7_75t_L g325 ( 
.A1(n_310),
.A2(n_7),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_14),
.C2(n_15),
.Y(n_325)
);

OAI21x1_ASAP7_75t_L g332 ( 
.A1(n_325),
.A2(n_7),
.B(n_11),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_7),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_326),
.B(n_315),
.Y(n_331)
);

OA21x2_ASAP7_75t_SL g330 ( 
.A1(n_324),
.A2(n_311),
.B(n_306),
.Y(n_330)
);

OAI31xp33_ASAP7_75t_L g337 ( 
.A1(n_330),
.A2(n_332),
.A3(n_327),
.B(n_328),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_331),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_334),
.A2(n_335),
.B(n_16),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_333),
.A2(n_322),
.B(n_321),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_336),
.A2(n_337),
.B(n_339),
.Y(n_340)
);

AOI322xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_329),
.A3(n_338),
.B1(n_14),
.B2(n_15),
.C1(n_16),
.C2(n_12),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_13),
.B(n_14),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_13),
.Y(n_343)
);


endmodule