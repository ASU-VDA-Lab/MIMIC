module fake_jpeg_21835_n_317 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_19),
.B(n_9),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_43),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_42),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_39),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_28),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_33),
.B1(n_32),
.B2(n_29),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_20),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_30),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_28),
.B1(n_23),
.B2(n_30),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_49),
.A2(n_42),
.B1(n_23),
.B2(n_25),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_21),
.Y(n_51)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_34),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_21),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_53),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_SL g69 ( 
.A1(n_55),
.A2(n_40),
.B(n_30),
.C(n_24),
.Y(n_69)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_27),
.B1(n_25),
.B2(n_24),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_25),
.B1(n_24),
.B2(n_27),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_20),
.B(n_27),
.C(n_23),
.Y(n_87)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_34),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_21),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_66),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_69),
.A2(n_83),
.B1(n_54),
.B2(n_18),
.Y(n_122)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_39),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_75),
.B(n_84),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_78),
.B(n_81),
.Y(n_117)
);

NOR2x1_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_39),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_79),
.B(n_49),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_43),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_91),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_64),
.B(n_19),
.Y(n_84)
);

OR2x2_ASAP7_75t_SL g86 ( 
.A(n_48),
.B(n_52),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_95),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_87),
.A2(n_94),
.B1(n_54),
.B2(n_65),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_19),
.Y(n_88)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_48),
.B(n_22),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_89),
.B(n_17),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_43),
.Y(n_91)
);

AO22x1_ASAP7_75t_SL g94 ( 
.A1(n_55),
.A2(n_42),
.B1(n_36),
.B2(n_20),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_31),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_22),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_97),
.B(n_98),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_22),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_99),
.A2(n_69),
.B(n_89),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_26),
.Y(n_100)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_70),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_102),
.Y(n_124)
);

INVx4_ASAP7_75t_SL g102 ( 
.A(n_70),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_50),
.C(n_57),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_109),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_26),
.Y(n_104)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_75),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_114),
.Y(n_126)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_108),
.A2(n_72),
.B1(n_71),
.B2(n_92),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_57),
.C(n_59),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_26),
.Y(n_111)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_113),
.B(n_32),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_75),
.Y(n_114)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_34),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_33),
.Y(n_116)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_31),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_63),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_119),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_79),
.B(n_33),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_121),
.A2(n_122),
.B1(n_94),
.B2(n_76),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_79),
.B(n_29),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_29),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_131),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_129),
.A2(n_96),
.B1(n_106),
.B2(n_110),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_SL g132 ( 
.A1(n_117),
.A2(n_94),
.B(n_69),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_107),
.C(n_100),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_119),
.A2(n_94),
.B(n_76),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_133),
.A2(n_106),
.B(n_104),
.Y(n_156)
);

OA21x2_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_69),
.B(n_87),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_134),
.A2(n_144),
.B(n_18),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_69),
.B1(n_83),
.B2(n_68),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_135),
.A2(n_138),
.B1(n_143),
.B2(n_145),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_96),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_99),
.A2(n_84),
.B1(n_93),
.B2(n_71),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_92),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_149),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_57),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_148),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_109),
.A2(n_93),
.B1(n_72),
.B2(n_77),
.Y(n_143)
);

AO21x1_ASAP7_75t_L g144 ( 
.A1(n_110),
.A2(n_118),
.B(n_123),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_103),
.A2(n_72),
.B1(n_62),
.B2(n_61),
.Y(n_145)
);

XOR2x2_ASAP7_75t_SL g160 ( 
.A(n_146),
.B(n_98),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_147),
.B(n_150),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_62),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_80),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_67),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_108),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_153),
.B(n_144),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_154),
.A2(n_176),
.B1(n_179),
.B2(n_182),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_156),
.A2(n_163),
.B(n_173),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_139),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_157),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_159),
.C(n_175),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_107),
.C(n_101),
.Y(n_159)
);

AO21x1_ASAP7_75t_L g199 ( 
.A1(n_160),
.A2(n_133),
.B(n_142),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_125),
.A2(n_108),
.B1(n_113),
.B2(n_97),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_161),
.B(n_167),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_111),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_162),
.Y(n_211)
);

OA21x2_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_61),
.B(n_67),
.Y(n_163)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_170),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_126),
.B(n_116),
.Y(n_170)
);

OAI32xp33_ASAP7_75t_L g171 ( 
.A1(n_137),
.A2(n_32),
.A3(n_20),
.B1(n_34),
.B2(n_47),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_141),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_124),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_172),
.B(n_174),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_149),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_148),
.A2(n_101),
.B(n_34),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_135),
.A2(n_102),
.B1(n_112),
.B2(n_115),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_151),
.A2(n_34),
.B(n_20),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_145),
.C(n_147),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_47),
.Y(n_178)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_129),
.A2(n_102),
.B1(n_112),
.B2(n_115),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_20),
.Y(n_180)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_134),
.A2(n_112),
.B(n_90),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_181),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_134),
.A2(n_20),
.B1(n_80),
.B2(n_90),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_80),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_183),
.B(n_131),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_184),
.B(n_10),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_190),
.A2(n_182),
.B1(n_166),
.B2(n_156),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_125),
.Y(n_193)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_162),
.B(n_142),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_195),
.B(n_152),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_210),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_168),
.A2(n_176),
.B1(n_179),
.B2(n_154),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_197),
.A2(n_205),
.B1(n_206),
.B2(n_171),
.Y(n_229)
);

FAx1_ASAP7_75t_SL g198 ( 
.A(n_158),
.B(n_137),
.CI(n_144),
.CON(n_198),
.SN(n_198)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_201),
.Y(n_212)
);

FAx1_ASAP7_75t_SL g216 ( 
.A(n_199),
.B(n_209),
.CI(n_180),
.CON(n_216),
.SN(n_216)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_130),
.Y(n_200)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

BUFx12_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

NAND3xp33_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_130),
.C(n_152),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_208),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_126),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_164),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_168),
.A2(n_163),
.B1(n_166),
.B2(n_181),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_163),
.A2(n_143),
.B1(n_138),
.B2(n_128),
.Y(n_206)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_167),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_155),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_191),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_213),
.A2(n_223),
.B1(n_232),
.B2(n_236),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_224),
.Y(n_250)
);

OA22x2_ASAP7_75t_SL g215 ( 
.A1(n_190),
.A2(n_163),
.B1(n_173),
.B2(n_175),
.Y(n_215)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_233),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_192),
.A2(n_172),
.B1(n_165),
.B2(n_157),
.Y(n_218)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_177),
.C(n_153),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_221),
.C(n_234),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_160),
.C(n_155),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_192),
.A2(n_194),
.B1(n_202),
.B2(n_197),
.Y(n_222)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_222),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_185),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_187),
.A2(n_141),
.B(n_170),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_225),
.A2(n_226),
.B(n_229),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_228),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_194),
.A2(n_164),
.B1(n_150),
.B2(n_80),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_230),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_187),
.A2(n_10),
.B(n_15),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_231),
.A2(n_211),
.B(n_188),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_208),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_0),
.C(n_1),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_207),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_232),
.Y(n_237)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_239),
.B(n_244),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_201),
.C(n_202),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_253),
.C(n_233),
.Y(n_260)
);

INVxp67_ASAP7_75t_SL g244 ( 
.A(n_215),
.Y(n_244)
);

NOR3xp33_ASAP7_75t_SL g246 ( 
.A(n_215),
.B(n_207),
.C(n_199),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_231),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_184),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_249),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_225),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_222),
.A2(n_226),
.B(n_223),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_1),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_206),
.C(n_209),
.Y(n_253)
);

NAND2xp33_ASAP7_75t_SL g255 ( 
.A(n_218),
.B(n_210),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_255),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_235),
.A2(n_219),
.B1(n_227),
.B2(n_217),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_257),
.A2(n_189),
.B1(n_216),
.B2(n_198),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_263),
.C(n_265),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_204),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_262),
.A2(n_243),
.B(n_251),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_188),
.C(n_228),
.Y(n_263)
);

AOI21xp33_ASAP7_75t_L g264 ( 
.A1(n_250),
.A2(n_216),
.B(n_198),
.Y(n_264)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_264),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_253),
.C(n_252),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_256),
.A2(n_189),
.B1(n_230),
.B2(n_229),
.Y(n_266)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_266),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_267),
.B(n_269),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_12),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_11),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_270),
.B(n_245),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_254),
.B1(n_243),
.B2(n_240),
.Y(n_275)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

HAxp5_ASAP7_75t_SL g274 ( 
.A(n_270),
.B(n_247),
.CON(n_274),
.SN(n_274)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_274),
.A2(n_276),
.B1(n_277),
.B2(n_7),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_275),
.B(n_282),
.Y(n_292)
);

OAI21xp33_ASAP7_75t_L g277 ( 
.A1(n_258),
.A2(n_246),
.B(n_251),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_261),
.A2(n_241),
.B(n_237),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_284),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_263),
.A2(n_245),
.B(n_248),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_283),
.C(n_260),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_265),
.A2(n_12),
.B(n_15),
.Y(n_284)
);

NOR2xp67_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_259),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_285),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_279),
.A2(n_268),
.B1(n_276),
.B2(n_262),
.Y(n_286)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_286),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_288),
.C(n_281),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_259),
.C(n_262),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_6),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_291),
.B(n_295),
.Y(n_296)
);

AOI21xp33_ASAP7_75t_L g293 ( 
.A1(n_277),
.A2(n_7),
.B(n_14),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_293),
.A2(n_7),
.B(n_14),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_272),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_295),
.B(n_273),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_297),
.B(n_301),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_288),
.C(n_287),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_294),
.A2(n_6),
.B(n_12),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_302),
.A2(n_13),
.B(n_16),
.Y(n_308)
);

AOI322xp5_ASAP7_75t_L g310 ( 
.A1(n_303),
.A2(n_4),
.A3(n_5),
.B1(n_237),
.B2(n_262),
.C1(n_277),
.C2(n_272),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_308),
.Y(n_312)
);

NAND3xp33_ASAP7_75t_SL g306 ( 
.A(n_299),
.B(n_286),
.C(n_290),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_307),
.B(n_309),
.Y(n_313)
);

AOI322xp5_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_292),
.A3(n_13),
.B1(n_16),
.B2(n_4),
.C1(n_5),
.C2(n_3),
.Y(n_307)
);

NOR2x1_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_13),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_310),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_304),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_296),
.Y(n_315)
);

OAI21x1_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_313),
.B(n_311),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_312),
.Y(n_317)
);


endmodule