module fake_jpeg_13924_n_61 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_61);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_61;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_22),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_31),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_28),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_33),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_4),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_25),
.C(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_36),
.B(n_37),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_28),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_5),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_40),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_44),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_45),
.A2(n_47),
.B1(n_15),
.B2(n_17),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_8),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_18),
.Y(n_53)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_49),
.B(n_55),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_48),
.C(n_52),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_53),
.B(n_51),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_19),
.B(n_20),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_21),
.Y(n_61)
);


endmodule