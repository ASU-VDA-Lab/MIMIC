module fake_jpeg_18975_n_212 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_212);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_212;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_19),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_0),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_28),
.C(n_34),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_18),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_52),
.B(n_53),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_25),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_26),
.B1(n_22),
.B2(n_21),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_55),
.A2(n_61),
.B1(n_18),
.B2(n_1),
.Y(n_87)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_62),
.Y(n_105)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_26),
.B1(n_20),
.B2(n_28),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_22),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_21),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_34),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_23),
.Y(n_100)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_39),
.A2(n_20),
.B1(n_29),
.B2(n_32),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_71),
.A2(n_73),
.B1(n_78),
.B2(n_42),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_38),
.B(n_32),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_72),
.B(n_74),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_20),
.B1(n_31),
.B2(n_29),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_31),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_19),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_75),
.B(n_30),
.Y(n_89)
);

BUFx10_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_44),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_86),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_54),
.B(n_30),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_83),
.A2(n_100),
.B(n_104),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_71),
.A2(n_46),
.B1(n_43),
.B2(n_33),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_84),
.A2(n_94),
.B1(n_95),
.B2(n_98),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_46),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_66),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_46),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_107),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_58),
.A2(n_43),
.B1(n_27),
.B2(n_24),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_27),
.B1(n_24),
.B2(n_18),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_61),
.A2(n_27),
.B1(n_24),
.B2(n_30),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_76),
.A2(n_42),
.B(n_23),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_76),
.A2(n_0),
.B(n_1),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_56),
.B(n_59),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_95),
.B1(n_83),
.B2(n_99),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_100),
.A2(n_106),
.B1(n_89),
.B2(n_87),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_111),
.A2(n_124),
.B1(n_125),
.B2(n_102),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_104),
.A2(n_63),
.B(n_54),
.C(n_79),
.Y(n_113)
);

O2A1O1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_113),
.A2(n_77),
.B(n_96),
.C(n_6),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_97),
.A2(n_70),
.B1(n_63),
.B2(n_48),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_121),
.B1(n_114),
.B2(n_96),
.Y(n_145)
);

XNOR2x1_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_86),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_118),
.B(n_83),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_97),
.A2(n_51),
.B1(n_2),
.B2(n_4),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_14),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_123),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_14),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_77),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_77),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_80),
.B(n_51),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_103),
.Y(n_144)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_130),
.Y(n_153)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_129),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_1),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_85),
.B(n_2),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_131),
.Y(n_148)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_132),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_140),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_136),
.A2(n_137),
.B(n_149),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_85),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_108),
.A2(n_83),
.B1(n_88),
.B2(n_93),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_139),
.A2(n_151),
.B1(n_119),
.B2(n_113),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_92),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_102),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_120),
.C(n_127),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_147),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_117),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_146),
.A2(n_150),
.B(n_132),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_111),
.A2(n_99),
.B1(n_102),
.B2(n_103),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_110),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_108),
.A2(n_96),
.B1(n_5),
.B2(n_7),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_4),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_109),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_154),
.A2(n_171),
.B1(n_167),
.B2(n_151),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_149),
.A2(n_114),
.B(n_119),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_137),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_157),
.A2(n_150),
.B1(n_153),
.B2(n_133),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_152),
.B(n_125),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_159),
.B(n_168),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_140),
.C(n_141),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_165),
.C(n_146),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_125),
.B(n_124),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_161),
.A2(n_139),
.B(n_136),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_144),
.B(n_115),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_166),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_126),
.C(n_124),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_117),
.Y(n_167)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_142),
.Y(n_170)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_170),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_182),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_169),
.C(n_156),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_180),
.C(n_128),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_176),
.A2(n_159),
.B(n_163),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_177),
.B(n_157),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_158),
.C(n_165),
.Y(n_180)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_184),
.A2(n_162),
.B1(n_161),
.B2(n_164),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_R g187 ( 
.A1(n_184),
.A2(n_171),
.B1(n_155),
.B2(n_158),
.Y(n_187)
);

AOI31xp67_ASAP7_75t_L g199 ( 
.A1(n_187),
.A2(n_181),
.A3(n_178),
.B(n_8),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_174),
.A2(n_170),
.B1(n_133),
.B2(n_134),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_190),
.A2(n_191),
.B(n_179),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_181),
.A2(n_142),
.B(n_129),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_183),
.A2(n_148),
.B1(n_138),
.B2(n_128),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_192),
.A2(n_176),
.B1(n_179),
.B2(n_175),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_182),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_173),
.C(n_172),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_195),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_196),
.A2(n_190),
.B(n_189),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_180),
.Y(n_197)
);

AO21x1_ASAP7_75t_L g202 ( 
.A1(n_199),
.A2(n_200),
.B(n_186),
.Y(n_202)
);

OA21x2_ASAP7_75t_SL g200 ( 
.A1(n_185),
.A2(n_178),
.B(n_7),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_203),
.Y(n_206)
);

FAx1_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_192),
.CI(n_188),
.CON(n_203),
.SN(n_203)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_198),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_205),
.B(n_207),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_201),
.A2(n_194),
.B1(n_197),
.B2(n_9),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_5),
.C(n_8),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_9),
.C(n_10),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_208),
.C(n_13),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_211),
.Y(n_212)
);


endmodule