module fake_jpeg_9464_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_45),
.Y(n_53)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_46),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_15),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_42),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_49),
.B(n_25),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_50),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_18),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_68),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_31),
.B1(n_27),
.B2(n_18),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_65),
.B1(n_48),
.B2(n_24),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_74),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_43),
.A2(n_31),
.B1(n_27),
.B2(n_18),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_64),
.A2(n_70),
.B1(n_72),
.B2(n_24),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_46),
.A2(n_31),
.B1(n_18),
.B2(n_29),
.Y(n_65)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_39),
.B(n_19),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_31),
.B1(n_19),
.B2(n_29),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_48),
.A2(n_19),
.B1(n_29),
.B2(n_35),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_36),
.B(n_26),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_73),
.B(n_22),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_34),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_36),
.B(n_35),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_47),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_SL g142 ( 
.A1(n_78),
.A2(n_104),
.B(n_115),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_89),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_SL g82 ( 
.A(n_51),
.B(n_22),
.C(n_25),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_82),
.A2(n_88),
.B(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_83),
.B(n_92),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_74),
.A2(n_72),
.B1(n_70),
.B2(n_69),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_84),
.A2(n_87),
.B1(n_96),
.B2(n_30),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_91),
.Y(n_127)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_53),
.B(n_21),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_62),
.A2(n_21),
.B(n_26),
.C(n_28),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_95),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_59),
.A2(n_35),
.B(n_28),
.C(n_22),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_69),
.A2(n_28),
.B1(n_34),
.B2(n_32),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_24),
.Y(n_97)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_114),
.B(n_47),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_53),
.A2(n_22),
.B(n_25),
.C(n_13),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_103),
.B(n_106),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_66),
.A2(n_34),
.B1(n_32),
.B2(n_30),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_14),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_50),
.B(n_40),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_109),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_58),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_52),
.B(n_40),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_113),
.Y(n_137)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_58),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_91),
.A2(n_61),
.B1(n_67),
.B2(n_52),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_116),
.A2(n_125),
.B1(n_132),
.B2(n_144),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_61),
.B1(n_55),
.B2(n_30),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_118),
.A2(n_133),
.B1(n_143),
.B2(n_109),
.Y(n_157)
);

NAND3xp33_ASAP7_75t_SL g119 ( 
.A(n_82),
.B(n_100),
.C(n_94),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_119),
.B(n_85),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_37),
.C(n_38),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_131),
.C(n_140),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_122),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_87),
.A2(n_55),
.B1(n_32),
.B2(n_38),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_126),
.A2(n_134),
.B(n_112),
.Y(n_155)
);

AND2x2_ASAP7_75t_SL g131 ( 
.A(n_89),
.B(n_38),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_90),
.A2(n_40),
.B1(n_16),
.B2(n_33),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_33),
.B1(n_23),
.B2(n_22),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_97),
.A2(n_20),
.B(n_25),
.Y(n_134)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_77),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_85),
.A2(n_23),
.B1(n_33),
.B2(n_20),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_138),
.A2(n_133),
.B1(n_127),
.B2(n_115),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_85),
.B(n_33),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_103),
.A2(n_23),
.B1(n_57),
.B2(n_56),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_95),
.A2(n_23),
.B1(n_25),
.B2(n_56),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_147),
.A2(n_129),
.B(n_14),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_97),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_149),
.B(n_161),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_150),
.A2(n_169),
.B1(n_170),
.B2(n_121),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_128),
.B(n_106),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_151),
.B(n_157),
.Y(n_187)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_176),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_142),
.A2(n_88),
.B1(n_113),
.B2(n_114),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_153),
.A2(n_165),
.B1(n_135),
.B2(n_146),
.Y(n_200)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_154),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_155),
.B(n_4),
.Y(n_208)
);

BUFx24_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_158),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_126),
.A2(n_88),
.B(n_110),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_160),
.A2(n_155),
.B(n_134),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_137),
.B(n_101),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_101),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_162),
.B(n_163),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_130),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_120),
.B(n_57),
.C(n_76),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_168),
.C(n_171),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_142),
.A2(n_107),
.B1(n_99),
.B2(n_81),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_130),
.B(n_93),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_174),
.Y(n_198)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_167),
.B(n_172),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_105),
.C(n_98),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_122),
.A2(n_98),
.B1(n_102),
.B2(n_80),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_128),
.A2(n_102),
.B1(n_80),
.B2(n_111),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_111),
.C(n_2),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_14),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_173),
.B(n_175),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_1),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_124),
.B(n_1),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_116),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_1),
.Y(n_177)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_2),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_178),
.Y(n_213)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_131),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_179),
.A2(n_180),
.B1(n_136),
.B2(n_145),
.Y(n_184)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_131),
.Y(n_180)
);

OAI32xp33_ASAP7_75t_L g181 ( 
.A1(n_149),
.A2(n_119),
.A3(n_143),
.B1(n_125),
.B2(n_117),
.Y(n_181)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_183),
.B(n_203),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_184),
.A2(n_5),
.B(n_6),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_117),
.C(n_131),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_188),
.B(n_197),
.C(n_209),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_134),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_194),
.C(n_205),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_138),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_167),
.A2(n_136),
.B1(n_121),
.B2(n_139),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_195),
.A2(n_202),
.B1(n_165),
.B2(n_179),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_144),
.C(n_139),
.Y(n_197)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_152),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_200),
.A2(n_201),
.B1(n_169),
.B2(n_172),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_176),
.A2(n_146),
.B1(n_132),
.B2(n_121),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_156),
.A2(n_129),
.B1(n_3),
.B2(n_4),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_204),
.A2(n_207),
.B1(n_213),
.B2(n_191),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_147),
.B(n_13),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_2),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_177),
.C(n_178),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_150),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_208),
.B(n_153),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_164),
.B(n_5),
.C(n_6),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_162),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_211),
.B(n_212),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_161),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_190),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_214),
.B(n_230),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_216),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_163),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_218),
.B(n_222),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_219),
.A2(n_237),
.B1(n_11),
.B2(n_8),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_198),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_175),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_223),
.Y(n_245)
);

XOR2x2_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_180),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_227),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_171),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_226),
.C(n_228),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_186),
.B(n_166),
.Y(n_226)
);

XNOR2x1_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_170),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_200),
.A2(n_148),
.B1(n_157),
.B2(n_151),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_229),
.A2(n_235),
.B1(n_204),
.B2(n_209),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_185),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_188),
.B(n_148),
.C(n_158),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_240),
.C(n_208),
.Y(n_246)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_192),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_233),
.Y(n_255)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_191),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_189),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_201),
.A2(n_158),
.B1(n_6),
.B2(n_7),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_202),
.B1(n_181),
.B2(n_207),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_199),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_239),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_186),
.B(n_7),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_238),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_259),
.Y(n_268)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_243),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_246),
.B(n_254),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_247),
.A2(n_253),
.B1(n_248),
.B2(n_251),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_224),
.A2(n_197),
.B(n_182),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_248),
.A2(n_227),
.B1(n_231),
.B2(n_245),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_194),
.C(n_189),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_252),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_253),
.A2(n_262),
.B1(n_215),
.B2(n_237),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_221),
.B(n_198),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_217),
.B(n_205),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_260),
.Y(n_281)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_217),
.B(n_203),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_210),
.Y(n_261)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_261),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_220),
.A2(n_182),
.B1(n_8),
.B2(n_9),
.Y(n_262)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_264),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_251),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_249),
.B(n_236),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_267),
.B(n_283),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_269),
.A2(n_272),
.B1(n_275),
.B2(n_254),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_229),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_270),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_259),
.A2(n_219),
.B1(n_215),
.B2(n_241),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_243),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_274),
.Y(n_291)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_255),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_247),
.A2(n_228),
.B1(n_226),
.B2(n_239),
.Y(n_275)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_256),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_282),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_279),
.A2(n_257),
.B1(n_8),
.B2(n_9),
.Y(n_298)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_258),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_261),
.B(n_240),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_250),
.C(n_244),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_289),
.C(n_293),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_268),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_286),
.A2(n_273),
.B(n_276),
.Y(n_306)
);

OA21x2_ASAP7_75t_SL g287 ( 
.A1(n_281),
.A2(n_260),
.B(n_246),
.Y(n_287)
);

NOR2xp67_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_280),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_288),
.B(n_281),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_244),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_299),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_252),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_268),
.Y(n_294)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_294),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_262),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_295),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_269),
.A2(n_258),
.B(n_263),
.Y(n_296)
);

AO21x1_ASAP7_75t_L g308 ( 
.A1(n_296),
.A2(n_298),
.B(n_274),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_277),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_301),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_282),
.Y(n_305)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_305),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_308),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_271),
.C(n_279),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_310),
.C(n_311),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_297),
.A2(n_271),
.B1(n_9),
.B2(n_10),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_299),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_7),
.C(n_11),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_292),
.C(n_294),
.Y(n_311)
);

AND2x2_ASAP7_75t_SL g313 ( 
.A(n_303),
.B(n_291),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_313),
.B(n_314),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_311),
.A2(n_286),
.B1(n_291),
.B2(n_288),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_285),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_318),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_302),
.B(n_293),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_310),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_304),
.C(n_307),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_325),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_304),
.C(n_302),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_328),
.Y(n_330)
);

MAJx2_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_300),
.C(n_308),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_327),
.A2(n_315),
.B(n_320),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_11),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_323),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_329),
.A2(n_324),
.B1(n_331),
.B2(n_313),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_324),
.Y(n_333)
);

AO21x1_ASAP7_75t_L g335 ( 
.A1(n_333),
.A2(n_334),
.B(n_314),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_318),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_336),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_330),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_319),
.Y(n_339)
);


endmodule