module real_jpeg_28269_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_337, n_11, n_14, n_336, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_337;
input n_11;
input n_14;
input n_336;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_324;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_0),
.A2(n_45),
.B1(n_48),
.B2(n_49),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_0),
.A2(n_45),
.B1(n_55),
.B2(n_56),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_0),
.A2(n_32),
.B1(n_33),
.B2(n_45),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_1),
.B(n_48),
.Y(n_90)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_1),
.Y(n_95)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_1),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_2),
.A2(n_55),
.B1(n_56),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_2),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_100),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_100),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_2),
.A2(n_48),
.B1(n_49),
.B2(n_100),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_3),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_L g182 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_105),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_3),
.A2(n_55),
.B1(n_56),
.B2(n_105),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_3),
.A2(n_48),
.B1(n_49),
.B2(n_105),
.Y(n_238)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_5),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_116),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_5),
.A2(n_55),
.B1(n_56),
.B2(n_116),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_5),
.A2(n_48),
.B1(n_49),
.B2(n_116),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_23)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_6),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_6),
.A2(n_27),
.B1(n_48),
.B2(n_49),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_6),
.A2(n_27),
.B1(n_55),
.B2(n_56),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_8),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_110),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_8),
.A2(n_55),
.B1(n_56),
.B2(n_110),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_8),
.A2(n_48),
.B1(n_49),
.B2(n_110),
.Y(n_233)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_10),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_107),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_10),
.A2(n_48),
.B1(n_49),
.B2(n_107),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_10),
.A2(n_55),
.B1(n_56),
.B2(n_107),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_11),
.A2(n_43),
.B1(n_55),
.B2(n_56),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_11),
.A2(n_43),
.B1(n_48),
.B2(n_49),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_43),
.Y(n_149)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_13),
.A2(n_48),
.B1(n_49),
.B2(n_52),
.Y(n_47)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_14),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_14),
.A2(n_36),
.B1(n_55),
.B2(n_56),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_14),
.A2(n_36),
.B1(n_48),
.B2(n_49),
.Y(n_129)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_16),
.Y(n_120)
);

AOI21xp33_ASAP7_75t_SL g121 ( 
.A1(n_16),
.A2(n_29),
.B(n_33),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_16),
.A2(n_24),
.B1(n_25),
.B2(n_120),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_16),
.B(n_31),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_16),
.A2(n_55),
.B(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_16),
.B(n_55),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_16),
.B(n_70),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_16),
.A2(n_89),
.B1(n_95),
.B2(n_244),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_16),
.A2(n_32),
.B(n_260),
.Y(n_259)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_17),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_80),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_78),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_37),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_21),
.B(n_37),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_28),
.B1(n_31),
.B2(n_35),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_23),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_74)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_29),
.Y(n_30)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_25),
.A2(n_34),
.B(n_120),
.C(n_121),
.Y(n_119)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_31),
.B1(n_41),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_28),
.A2(n_31),
.B1(n_104),
.B2(n_106),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_28),
.A2(n_31),
.B1(n_106),
.B2(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_28),
.A2(n_31),
.B1(n_115),
.B2(n_188),
.Y(n_187)
);

AO22x1_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_31),
.Y(n_77)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_32),
.A2(n_62),
.B(n_64),
.C(n_65),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_32),
.B(n_62),
.Y(n_64)
);

OAI32xp33_ASAP7_75t_L g268 ( 
.A1(n_32),
.A2(n_56),
.A3(n_66),
.B1(n_261),
.B2(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_33),
.B(n_120),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_71),
.C(n_73),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_38),
.A2(n_39),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.C(n_59),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_40),
.B(n_317),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_42),
.A2(n_75),
.B1(n_77),
.B2(n_168),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_44),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_46),
.A2(n_308),
.B1(n_310),
.B2(n_311),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_46),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_46),
.A2(n_59),
.B1(n_311),
.B2(n_318),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_53),
.B(n_58),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_47),
.A2(n_53),
.B1(n_98),
.B2(n_101),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_47),
.A2(n_53),
.B1(n_101),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_47),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_47),
.A2(n_53),
.B1(n_58),
.B2(n_140),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_47),
.A2(n_53),
.B1(n_217),
.B2(n_219),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_47),
.A2(n_53),
.B1(n_219),
.B2(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_47),
.B(n_120),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_47),
.A2(n_53),
.B1(n_186),
.B2(n_286),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_48),
.B(n_52),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_48),
.B(n_249),
.Y(n_248)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI32xp33_ASAP7_75t_L g221 ( 
.A1(n_49),
.A2(n_55),
.A3(n_57),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_54)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_53),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_55),
.A2(n_56),
.B1(n_63),
.B2(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_55),
.B(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_59),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_60),
.A2(n_70),
.B1(n_109),
.B2(n_111),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_60),
.A2(n_70),
.B1(n_111),
.B2(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_60),
.A2(n_70),
.B1(n_182),
.B2(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_60),
.A2(n_68),
.B1(n_70),
.B2(n_309),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_65),
.B(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_61),
.A2(n_65),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_61),
.A2(n_65),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_61),
.A2(n_65),
.B1(n_125),
.B2(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_61),
.A2(n_65),
.B1(n_194),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_66),
.Y(n_270)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_69),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_71),
.A2(n_73),
.B1(n_74),
.B2(n_331),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_71),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_75),
.A2(n_77),
.B1(n_114),
.B2(n_117),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_75),
.A2(n_77),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_326),
.B(n_332),
.Y(n_80)
);

OAI321xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_302),
.A3(n_321),
.B1(n_324),
.B2(n_325),
.C(n_336),
.Y(n_81)
);

AOI321xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_152),
.A3(n_174),
.B1(n_296),
.B2(n_301),
.C(n_337),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_84),
.A2(n_297),
.B(n_300),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_132),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_85),
.B(n_132),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_112),
.C(n_127),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_86),
.B(n_127),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_102),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_87),
.B(n_103),
.C(n_108),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_97),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_88),
.B(n_97),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_91),
.B1(n_93),
.B2(n_96),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_89),
.A2(n_93),
.B1(n_96),
.B2(n_129),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_89),
.A2(n_129),
.B(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_89),
.A2(n_144),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_89),
.A2(n_95),
.B1(n_238),
.B2(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_89),
.A2(n_144),
.B1(n_233),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_90),
.A2(n_92),
.B1(n_94),
.B2(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_90),
.A2(n_94),
.B1(n_123),
.B2(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_90),
.A2(n_94),
.B1(n_237),
.B2(n_239),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx5_ASAP7_75t_SL g144 ( 
.A(n_94),
.Y(n_144)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_99),
.A2(n_138),
.B1(n_141),
.B2(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_104),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_109),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_112),
.B(n_208),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_118),
.C(n_124),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_113),
.B(n_124),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_118),
.B(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_119),
.B(n_122),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_120),
.B(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_130),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_131),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_151),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_145),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_145),
.C(n_151),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_142),
.B2(n_143),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_135),
.B(n_143),
.Y(n_170)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_141),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_138),
.A2(n_141),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_143),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_142),
.A2(n_166),
.B(n_169),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_145),
.Y(n_335)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_148),
.CI(n_150),
.CON(n_145),
.SN(n_145)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_148),
.C(n_150),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_147),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_149),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_153),
.B(n_154),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_172),
.B2(n_173),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_163),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_157),
.B(n_163),
.C(n_173),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_161),
.B(n_162),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_161),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_160),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_162),
.B(n_304),
.C(n_313),
.Y(n_303)
);

FAx1_ASAP7_75t_SL g323 ( 
.A(n_162),
.B(n_304),
.CI(n_313),
.CON(n_323),
.SN(n_323)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_163)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_172),
.Y(n_173)
);

NOR3xp33_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_204),
.C(n_209),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_198),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_176),
.B(n_198),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_189),
.C(n_190),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_177),
.B(n_293),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_187),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_183),
.B2(n_184),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_184),
.C(n_187),
.Y(n_201)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_294),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_189),
.Y(n_294)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.C(n_197),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_192),
.B(n_281),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_195),
.B(n_197),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_196),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_201),
.C(n_202),
.Y(n_206)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

AOI21xp33_ASAP7_75t_L g297 ( 
.A1(n_205),
.A2(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_206),
.B(n_207),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_290),
.B(n_295),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_276),
.B(n_289),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_254),
.B(n_275),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_234),
.B(n_253),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_224),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_214),
.B(n_224),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_220),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_215),
.A2(n_216),
.B1(n_220),
.B2(n_221),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_218),
.Y(n_222)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_231),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_229),
.C(n_231),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_230),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_232),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_241),
.B(n_252),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_240),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_236),
.B(n_240),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_246),
.B(n_251),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_243),
.B(n_245),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_255),
.B(n_256),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_267),
.B1(n_273),
.B2(n_274),
.Y(n_256)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_262),
.B1(n_265),
.B2(n_266),
.Y(n_257)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_258),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_262),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_266),
.C(n_274),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_264),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_267),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_271),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_271),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_277),
.B(n_278),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_282),
.B2(n_283),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_285),
.C(n_287),
.Y(n_291)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_287),
.B2(n_288),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_284),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_285),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_291),
.B(n_292),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_314),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_303),
.B(n_314),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_312),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_305),
.A2(n_306),
.B1(n_316),
.B2(n_319),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_308),
.C(n_311),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_306),
.B(n_319),
.C(n_320),
.Y(n_327)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_307),
.Y(n_312)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_308),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_320),
.Y(n_314)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_316),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_322),
.B(n_323),
.Y(n_324)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_323),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_328),
.Y(n_332)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);


endmodule