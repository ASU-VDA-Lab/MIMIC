module fake_jpeg_30163_n_72 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_72);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_72;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_71;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_32;
wire n_70;
wire n_66;

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_22),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_19),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_11),
.B(n_21),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_32),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_28),
.B1(n_24),
.B2(n_23),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_48),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_47),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_37),
.Y(n_59)
);

OR2x2_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_4),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_50),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_5),
.B(n_6),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_52),
.C(n_44),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_6),
.B(n_7),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_56),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_48),
.A2(n_37),
.B1(n_9),
.B2(n_10),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_59),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_53),
.A2(n_8),
.B1(n_12),
.B2(n_14),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_15),
.Y(n_64)
);

BUFx24_ASAP7_75t_SL g62 ( 
.A(n_54),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_64),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_57),
.C(n_61),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_65),
.Y(n_68)
);

MAJx2_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_66),
.C(n_61),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_58),
.C(n_18),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_17),
.C(n_20),
.Y(n_72)
);


endmodule