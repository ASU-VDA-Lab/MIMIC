module real_jpeg_1453_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_17;
wire n_37;
wire n_21;
wire n_35;
wire n_33;
wire n_29;
wire n_31;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_14;
wire n_25;
wire n_22;
wire n_18;
wire n_36;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_0),
.B(n_7),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_1),
.B(n_5),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_1),
.B(n_5),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_2),
.B(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_2),
.B(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_4),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_3),
.B(n_4),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_4),
.B(n_17),
.C(n_19),
.Y(n_16)
);

AOI322xp5_ASAP7_75t_SL g11 ( 
.A1(n_6),
.A2(n_12),
.A3(n_31),
.B1(n_32),
.B2(n_34),
.C1(n_35),
.C2(n_37),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_7),
.B(n_14),
.Y(n_13)
);

INVx5_ASAP7_75t_SL g34 ( 
.A(n_7),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_8),
.B(n_16),
.C(n_20),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_15),
.B1(n_21),
.B2(n_22),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_13),
.A2(n_21),
.B1(n_23),
.B2(n_36),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_25),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_26),
.B(n_30),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B(n_29),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_31),
.B(n_32),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);


endmodule