module fake_jpeg_2370_n_68 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_68);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_68;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_29),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_21),
.A2(n_18),
.B1(n_17),
.B2(n_16),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_20),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_25),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_24),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_33),
.B(n_35),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_42),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_35),
.A2(n_19),
.B(n_20),
.Y(n_40)
);

INVxp67_ASAP7_75t_SL g48 ( 
.A(n_40),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_29),
.B1(n_26),
.B2(n_21),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_34),
.Y(n_42)
);

O2A1O1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_15),
.B(n_14),
.C(n_12),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_44),
.Y(n_52)
);

NOR2x1_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_39),
.C(n_40),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_51),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_2),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_SL g55 ( 
.A(n_53),
.B(n_54),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_3),
.Y(n_54)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_58),
.Y(n_60)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_52),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_4),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_56),
.A2(n_47),
.B1(n_44),
.B2(n_8),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_55),
.Y(n_63)
);

OAI21x1_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_4),
.B(n_7),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_SL g65 ( 
.A1(n_63),
.A2(n_64),
.B(n_55),
.C(n_60),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_66),
.A2(n_7),
.B(n_8),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_9),
.Y(n_68)
);


endmodule