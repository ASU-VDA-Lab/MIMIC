module fake_jpeg_9861_n_109 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_109);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_109;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx10_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_32),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_50),
.B(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_0),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_4),
.Y(n_68)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_1),
.Y(n_65)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_55),
.Y(n_61)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_53),
.A2(n_43),
.B1(n_38),
.B2(n_44),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_63),
.A2(n_66),
.B1(n_72),
.B2(n_78),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_67),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_48),
.B1(n_37),
.B2(n_2),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_2),
.Y(n_67)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_73),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_42),
.B1(n_40),
.B2(n_8),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_5),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_74),
.B(n_76),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_6),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_9),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_81),
.C(n_16),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_13),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

OAI32xp33_ASAP7_75t_L g95 ( 
.A1(n_88),
.A2(n_89),
.A3(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_61),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

NAND2xp33_ASAP7_75t_SL g92 ( 
.A(n_71),
.B(n_17),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_96),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_97),
.A2(n_87),
.B1(n_64),
.B2(n_65),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_98),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_99),
.A2(n_93),
.B1(n_95),
.B2(n_94),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_94),
.B1(n_75),
.B2(n_83),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_102),
.A2(n_84),
.B(n_67),
.Y(n_103)
);

XOR2x2_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_69),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_85),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_18),
.B(n_21),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_23),
.B(n_24),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_25),
.Y(n_109)
);


endmodule