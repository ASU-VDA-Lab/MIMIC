module fake_jpeg_27944_n_310 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_310);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_310;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_9),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx2_ASAP7_75t_SL g43 ( 
.A(n_37),
.Y(n_43)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_41),
.Y(n_47)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_0),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_28),
.B1(n_27),
.B2(n_31),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_46),
.A2(n_50),
.B1(n_42),
.B2(n_40),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_18),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_53),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_28),
.B1(n_18),
.B2(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_55),
.Y(n_81)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_33),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_61),
.Y(n_63)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_29),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_32),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_66),
.B(n_71),
.Y(n_112)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_68),
.B(n_70),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_54),
.A2(n_28),
.B1(n_35),
.B2(n_34),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_69),
.A2(n_83),
.B1(n_85),
.B2(n_42),
.Y(n_100)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_16),
.B1(n_17),
.B2(n_20),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_80),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_37),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_37),
.Y(n_95)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_53),
.A2(n_35),
.B1(n_34),
.B2(n_16),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_35),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_84),
.A2(n_57),
.B1(n_58),
.B2(n_62),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_55),
.A2(n_35),
.B1(n_34),
.B2(n_36),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_35),
.C(n_36),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_36),
.C(n_59),
.Y(n_98)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_42),
.B1(n_40),
.B2(n_52),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_92),
.A2(n_97),
.B1(n_106),
.B2(n_107),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_95),
.B(n_81),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_72),
.A2(n_42),
.B1(n_40),
.B2(n_48),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_108),
.C(n_63),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_100),
.A2(n_109),
.B(n_115),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_76),
.A2(n_42),
.B1(n_38),
.B2(n_36),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_101),
.A2(n_102),
.B1(n_87),
.B2(n_71),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_48),
.B1(n_38),
.B2(n_36),
.Y(n_102)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_84),
.A2(n_49),
.B1(n_57),
.B2(n_44),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_84),
.A2(n_57),
.B1(n_44),
.B2(n_58),
.Y(n_107)
);

AOI21xp33_ASAP7_75t_L g108 ( 
.A1(n_63),
.A2(n_22),
.B(n_33),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_70),
.A2(n_62),
.B1(n_45),
.B2(n_22),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_73),
.B1(n_74),
.B2(n_66),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_82),
.A2(n_17),
.B1(n_20),
.B2(n_45),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_116),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_118),
.B1(n_128),
.B2(n_136),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_81),
.B1(n_86),
.B2(n_78),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_123),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_103),
.B1(n_96),
.B2(n_105),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_122),
.B(n_25),
.Y(n_175)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_124),
.A2(n_99),
.B1(n_113),
.B2(n_75),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_93),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_139),
.Y(n_154)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_132),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_94),
.A2(n_78),
.B1(n_89),
.B2(n_77),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_91),
.A2(n_77),
.B1(n_67),
.B2(n_65),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_130),
.A2(n_131),
.B1(n_133),
.B2(n_138),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_91),
.A2(n_67),
.B1(n_37),
.B2(n_31),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_91),
.A2(n_37),
.B1(n_30),
.B2(n_19),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_110),
.B(n_105),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_142),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_94),
.A2(n_37),
.B1(n_30),
.B2(n_19),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_95),
.A2(n_109),
.B1(n_92),
.B2(n_106),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_137),
.A2(n_114),
.B1(n_103),
.B2(n_96),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_102),
.A2(n_21),
.B1(n_31),
.B2(n_30),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_116),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_141),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_90),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_98),
.B(n_59),
.C(n_75),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_137),
.C(n_130),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_90),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_26),
.Y(n_173)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_59),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_135),
.A2(n_115),
.B1(n_114),
.B2(n_104),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_166),
.B1(n_176),
.B2(n_136),
.Y(n_178)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_151),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_149),
.A2(n_150),
.B1(n_152),
.B2(n_159),
.Y(n_189)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_121),
.C(n_129),
.Y(n_184)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_164),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_25),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_158),
.B(n_175),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_124),
.A2(n_99),
.B1(n_29),
.B2(n_2),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_161),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_123),
.A2(n_29),
.B1(n_1),
.B2(n_2),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_119),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_135),
.A2(n_0),
.B(n_1),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_165),
.A2(n_168),
.B(n_172),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_145),
.A2(n_59),
.B1(n_31),
.B2(n_30),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_171),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_131),
.A2(n_1),
.B(n_2),
.Y(n_172)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_121),
.A2(n_26),
.B1(n_23),
.B2(n_21),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_174),
.A2(n_138),
.B1(n_132),
.B2(n_127),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_142),
.A2(n_26),
.B1(n_23),
.B2(n_21),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_178),
.A2(n_177),
.B1(n_154),
.B2(n_166),
.Y(n_218)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_179),
.Y(n_211)
);

XNOR2x1_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_118),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_180),
.B(n_162),
.Y(n_215)
);

XOR2x1_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_133),
.Y(n_183)
);

XOR2x1_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_146),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_186),
.C(n_174),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_165),
.A2(n_125),
.B(n_139),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_185),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_129),
.C(n_140),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_171),
.B(n_25),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_187),
.B(n_13),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_169),
.A2(n_150),
.B(n_167),
.Y(n_190)
);

NAND2xp33_ASAP7_75t_SL g225 ( 
.A(n_190),
.B(n_3),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_144),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_170),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_157),
.A2(n_141),
.B1(n_26),
.B2(n_23),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_195),
.A2(n_199),
.B1(n_203),
.B2(n_172),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_146),
.A2(n_23),
.B1(n_21),
.B2(n_5),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_156),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_202),
.Y(n_207)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_148),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_155),
.A2(n_3),
.B(n_4),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_205),
.Y(n_209)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

OAI32xp33_ASAP7_75t_L g206 ( 
.A1(n_183),
.A2(n_164),
.A3(n_155),
.B1(n_168),
.B2(n_153),
.Y(n_206)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_206),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_208),
.A2(n_225),
.B(n_181),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_210),
.A2(n_218),
.B1(n_227),
.B2(n_229),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_162),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_217),
.Y(n_235)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_214),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_197),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_215),
.B(n_184),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_15),
.Y(n_219)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_226),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_193),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_223),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_186),
.Y(n_222)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_222),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_193),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_170),
.C(n_15),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_185),
.C(n_180),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_14),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_190),
.B(n_12),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_228),
.A2(n_204),
.B1(n_194),
.B2(n_182),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_208),
.A2(n_189),
.B1(n_199),
.B2(n_194),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_231),
.A2(n_246),
.B1(n_216),
.B2(n_214),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_209),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_234),
.A2(n_240),
.B1(n_229),
.B2(n_13),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_248),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_192),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_243),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_215),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_211),
.A2(n_178),
.B1(n_192),
.B2(n_195),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_210),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_211),
.A2(n_179),
.B1(n_181),
.B2(n_188),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_198),
.C(n_200),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_226),
.C(n_213),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_198),
.Y(n_248)
);

XOR2x1_ASAP7_75t_SL g249 ( 
.A(n_240),
.B(n_225),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_257),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_244),
.A2(n_207),
.B(n_241),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_251),
.A2(n_248),
.B(n_239),
.Y(n_266)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_252),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_260),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_231),
.A2(n_232),
.B1(n_246),
.B2(n_238),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_258),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_263),
.C(n_262),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_206),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_223),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_261),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_12),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_234),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_12),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_3),
.Y(n_274)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_266),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_253),
.A2(n_243),
.B(n_242),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_269),
.A2(n_275),
.B(n_249),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_235),
.C(n_237),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_273),
.C(n_262),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_239),
.C(n_11),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_274),
.B(n_276),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_254),
.A2(n_4),
.B(n_5),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_269),
.C(n_271),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_6),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_255),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_280),
.B(n_283),
.Y(n_288)
);

FAx1_ASAP7_75t_SL g281 ( 
.A(n_272),
.B(n_273),
.CI(n_264),
.CON(n_281),
.SN(n_281)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_282),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_267),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_255),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_4),
.C(n_6),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_275),
.C(n_7),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_276),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_286),
.A2(n_6),
.B(n_7),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_4),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_274),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_292),
.Y(n_298)
);

INVxp33_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_294),
.Y(n_301)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_291),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_295),
.A2(n_7),
.B(n_8),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_293),
.A2(n_284),
.B1(n_279),
.B2(n_286),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_297),
.B(n_299),
.Y(n_302)
);

OAI21x1_ASAP7_75t_L g300 ( 
.A1(n_290),
.A2(n_281),
.B(n_285),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_277),
.Y(n_303)
);

O2A1O1Ixp33_ASAP7_75t_SL g305 ( 
.A1(n_303),
.A2(n_304),
.B(n_301),
.C(n_296),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_298),
.A2(n_288),
.B(n_281),
.Y(n_304)
);

AOI21x1_ASAP7_75t_SL g306 ( 
.A1(n_305),
.A2(n_302),
.B(n_294),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_292),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_7),
.B(n_9),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_308),
.B(n_10),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_10),
.Y(n_310)
);


endmodule