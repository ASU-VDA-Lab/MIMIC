module fake_jpeg_3290_n_181 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_181);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_181;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx14_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_5),
.B(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

BUFx12f_ASAP7_75t_SL g32 ( 
.A(n_16),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_32),
.B(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_17),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_48),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_0),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_15),
.B(n_28),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_53),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

AOI21xp33_ASAP7_75t_L g51 ( 
.A1(n_14),
.A2(n_0),
.B(n_1),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_51),
.B(n_2),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_10),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_54),
.A2(n_28),
.B1(n_15),
.B2(n_25),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_29),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_56),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_14),
.B(n_1),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_29),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_SL g104 ( 
.A1(n_61),
.A2(n_69),
.B(n_72),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_73),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_42),
.A2(n_18),
.B1(n_25),
.B2(n_23),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_86),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_37),
.A2(n_23),
.B1(n_22),
.B2(n_19),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_45),
.B(n_22),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_19),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_76),
.B(n_87),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_31),
.A2(n_18),
.B1(n_3),
.B2(n_8),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_81),
.A2(n_50),
.B1(n_53),
.B2(n_57),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_41),
.B(n_2),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_88),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_35),
.B(n_3),
.C(n_8),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_38),
.B(n_9),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_9),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_10),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_75),
.A2(n_54),
.B(n_11),
.C(n_10),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_92),
.B(n_98),
.Y(n_123)
);

NAND2xp33_ASAP7_75t_SL g93 ( 
.A(n_83),
.B(n_34),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_106),
.Y(n_129)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_85),
.B(n_50),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_95),
.B(n_103),
.Y(n_117)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_107),
.B1(n_79),
.B2(n_60),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_40),
.B1(n_53),
.B2(n_57),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_64),
.B1(n_79),
.B2(n_63),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_34),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_105),
.B(n_110),
.Y(n_128)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_69),
.A2(n_72),
.B1(n_61),
.B2(n_63),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_109),
.B(n_62),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_77),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_66),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_93),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_113),
.B(n_127),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_83),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_116),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_70),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_90),
.C(n_65),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_111),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_122),
.B1(n_131),
.B2(n_97),
.Y(n_140)
);

AOI32xp33_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_60),
.A3(n_65),
.B1(n_64),
.B2(n_62),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_130),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_107),
.A2(n_58),
.B1(n_62),
.B2(n_104),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_126),
.A2(n_92),
.B(n_101),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_110),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_94),
.A2(n_96),
.B1(n_109),
.B2(n_100),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

AOI21x1_ASAP7_75t_L g150 ( 
.A1(n_134),
.A2(n_113),
.B(n_129),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_118),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_126),
.A2(n_102),
.B1(n_99),
.B2(n_103),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_136),
.A2(n_140),
.B1(n_116),
.B2(n_115),
.Y(n_149)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_142),
.B(n_144),
.Y(n_148)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_114),
.Y(n_146)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_146),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_150),
.B1(n_129),
.B2(n_117),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_128),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_151),
.B(n_152),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_133),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_135),
.C(n_95),
.Y(n_157)
);

AOI322xp5_ASAP7_75t_L g156 ( 
.A1(n_151),
.A2(n_138),
.A3(n_137),
.B1(n_139),
.B2(n_123),
.C1(n_134),
.C2(n_136),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_156),
.A2(n_149),
.B1(n_145),
.B2(n_150),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_160),
.C(n_145),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_128),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_158),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_144),
.C(n_129),
.Y(n_160)
);

XNOR2x1_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_160),
.Y(n_166)
);

OAI322xp33_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_117),
.A3(n_108),
.B1(n_91),
.B2(n_98),
.C1(n_141),
.C2(n_143),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_162),
.A2(n_91),
.B(n_108),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_163),
.B(n_165),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_166),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_167),
.B(n_155),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_171),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_164),
.B(n_157),
.Y(n_171)
);

MAJx2_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_166),
.C(n_159),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_172),
.A2(n_174),
.B(n_159),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_169),
.C(n_147),
.Y(n_174)
);

MAJx2_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_122),
.C(n_125),
.Y(n_178)
);

NAND2xp67_ASAP7_75t_SL g176 ( 
.A(n_173),
.B(n_147),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_146),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_178),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_106),
.Y(n_180)
);

FAx1_ASAP7_75t_SL g181 ( 
.A(n_180),
.B(n_178),
.CI(n_176),
.CON(n_181),
.SN(n_181)
);


endmodule