module fake_jpeg_9258_n_268 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_268);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_268;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_175;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx5p33_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_6),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_20),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_37),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx2_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_28),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_20),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_43),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_0),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_31),
.B1(n_26),
.B2(n_33),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_46),
.A2(n_66),
.B1(n_23),
.B2(n_24),
.Y(n_85)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_51),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_61),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_29),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_55),
.B(n_63),
.Y(n_76)
);

OR2x4_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_68),
.Y(n_80)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_60),
.B1(n_31),
.B2(n_25),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_23),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_25),
.B1(n_22),
.B2(n_42),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_31),
.B1(n_25),
.B2(n_26),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_24),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_36),
.A2(n_31),
.B1(n_26),
.B2(n_33),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_L g68 ( 
.A1(n_37),
.A2(n_17),
.B(n_18),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_35),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_83),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_70),
.A2(n_78),
.B1(n_84),
.B2(n_67),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_35),
.B1(n_33),
.B2(n_39),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_74),
.A2(n_79),
.B1(n_85),
.B2(n_87),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_88),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_77),
.B(n_90),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_53),
.A2(n_22),
.B1(n_33),
.B2(n_30),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_46),
.A2(n_39),
.B1(n_45),
.B2(n_22),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_38),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_64),
.A2(n_22),
.B1(n_23),
.B2(n_29),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_45),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_52),
.B(n_27),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_73),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_93),
.Y(n_117)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_70),
.B(n_69),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_80),
.B(n_38),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_77),
.C(n_29),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_73),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_97),
.Y(n_121)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_99),
.Y(n_123)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_101),
.Y(n_125)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_105),
.Y(n_132)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_104),
.Y(n_130)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

OAI32xp33_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_47),
.A3(n_24),
.B1(n_30),
.B2(n_28),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_76),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_50),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_108),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_50),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_111),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_19),
.Y(n_112)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_78),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_74),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_115),
.A2(n_118),
.B(n_16),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_80),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_122),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_85),
.B1(n_81),
.B2(n_76),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_126),
.A2(n_109),
.B1(n_101),
.B2(n_92),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_88),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_136),
.Y(n_153)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_134),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_135),
.C(n_119),
.Y(n_146)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_39),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_28),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_136),
.A2(n_98),
.B(n_93),
.Y(n_152)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_97),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_109),
.A2(n_49),
.B1(n_57),
.B2(n_48),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_138),
.A2(n_105),
.B1(n_100),
.B2(n_111),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_139),
.A2(n_143),
.B1(n_162),
.B2(n_155),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_117),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_140),
.B(n_145),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_113),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_144),
.B(n_156),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_128),
.B(n_102),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_124),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_115),
.A2(n_113),
.B(n_92),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_147),
.A2(n_148),
.B(n_152),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_121),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_133),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_149),
.B(n_163),
.C(n_164),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_150),
.Y(n_166)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_153),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_131),
.B1(n_82),
.B2(n_124),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_54),
.B(n_82),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_155),
.A2(n_158),
.B(n_152),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_127),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_132),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_159),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_134),
.A2(n_30),
.B(n_27),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_16),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_138),
.A2(n_100),
.B1(n_99),
.B2(n_82),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_160),
.A2(n_130),
.B1(n_131),
.B2(n_126),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_161),
.A2(n_130),
.B(n_129),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_136),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_129),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_62),
.C(n_54),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_120),
.B(n_65),
.C(n_99),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_165),
.A2(n_172),
.B1(n_0),
.B2(n_1),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_176),
.B1(n_180),
.B2(n_157),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_177),
.C(n_148),
.Y(n_193)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_171),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_161),
.A2(n_147),
.B(n_156),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_116),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_181),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_19),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_179),
.A2(n_182),
.B1(n_158),
.B2(n_142),
.Y(n_190)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_140),
.B(n_27),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_163),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_186),
.Y(n_200)
);

XOR2x2_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_19),
.Y(n_185)
);

XOR2x2_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_160),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_16),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_184),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_199),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_190),
.A2(n_204),
.B1(n_166),
.B2(n_183),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_159),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_193),
.C(n_198),
.Y(n_208)
);

MAJx2_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_144),
.C(n_139),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_195),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_178),
.B(n_154),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_196),
.A2(n_168),
.B(n_173),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_167),
.A2(n_151),
.B1(n_21),
.B2(n_15),
.Y(n_197)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_177),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_21),
.C(n_19),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_202),
.C(n_186),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_169),
.B(n_21),
.C(n_19),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_168),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_205),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_174),
.A2(n_13),
.B1(n_14),
.B2(n_2),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_174),
.B(n_14),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_207),
.A2(n_182),
.B(n_178),
.Y(n_210)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_165),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_214),
.C(n_215),
.Y(n_226)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_166),
.Y(n_213)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_179),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_221),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_170),
.C(n_180),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_223),
.C(n_208),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_170),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_175),
.C(n_13),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_209),
.B(n_189),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_225),
.B(n_228),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_196),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_192),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_229),
.B(n_235),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_216),
.B(n_175),
.Y(n_232)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_232),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_200),
.Y(n_233)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_233),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_234),
.B(n_220),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_206),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_238),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_219),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_224),
.A2(n_199),
.B(n_208),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_239),
.B(n_3),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_223),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_12),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_228),
.A2(n_227),
.B1(n_229),
.B2(n_226),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_242),
.A2(n_244),
.B1(n_3),
.B2(n_4),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_214),
.B1(n_202),
.B2(n_2),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_240),
.A2(n_234),
.B1(n_1),
.B2(n_2),
.Y(n_246)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_246),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_0),
.Y(n_248)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_1),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_6),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_253),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_252),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_4),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_245),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_256),
.A2(n_246),
.B(n_7),
.Y(n_262)
);

INVxp67_ASAP7_75t_SL g260 ( 
.A(n_258),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_242),
.C(n_237),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_261),
.B(n_262),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_6),
.Y(n_263)
);

AOI322xp5_ASAP7_75t_L g265 ( 
.A1(n_263),
.A2(n_259),
.A3(n_254),
.B1(n_257),
.B2(n_11),
.C1(n_8),
.C2(n_10),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_265),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_266),
.A2(n_264),
.B1(n_260),
.B2(n_7),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_267),
.B(n_7),
.Y(n_268)
);


endmodule