module fake_jpeg_14511_n_444 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_444);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_444;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_SL g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_11),
.B(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_21),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_61),
.Y(n_96)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_16),
.B(n_15),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_54),
.B(n_59),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_56),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_16),
.B(n_15),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_21),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_42),
.B(n_15),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_64),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_63),
.Y(n_136)
);

BUFx16f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx4f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_67),
.Y(n_120)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_70),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_42),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_72),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_19),
.B(n_14),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_17),
.B(n_14),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_75),
.Y(n_109)
);

BUFx24_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g141 ( 
.A(n_74),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_17),
.B(n_0),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_19),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_80),
.Y(n_126)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_22),
.B(n_12),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_84),
.Y(n_115)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_26),
.B(n_1),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_90),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_22),
.B(n_12),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_1),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_49),
.A2(n_46),
.B1(n_27),
.B2(n_18),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_93),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_74),
.A2(n_34),
.B1(n_38),
.B2(n_18),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_103),
.A2(n_124),
.B1(n_144),
.B2(n_91),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_111),
.B(n_129),
.Y(n_154)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

BUFx24_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_55),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_64),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_50),
.A2(n_46),
.B1(n_36),
.B2(n_31),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_39),
.Y(n_129)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_130),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_57),
.A2(n_46),
.B1(n_27),
.B2(n_37),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_132),
.A2(n_37),
.B1(n_51),
.B2(n_56),
.Y(n_165)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_69),
.Y(n_139)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_87),
.A2(n_36),
.B1(n_31),
.B2(n_24),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_140),
.A2(n_33),
.B1(n_45),
.B2(n_43),
.Y(n_185)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_47),
.A2(n_34),
.B1(n_38),
.B2(n_37),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_58),
.C(n_76),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_145),
.B(n_120),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_127),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_146),
.B(n_153),
.Y(n_209)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_124),
.A2(n_66),
.B1(n_36),
.B2(n_31),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_148),
.A2(n_165),
.B1(n_174),
.B2(n_190),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_114),
.Y(n_152)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_152),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_102),
.Y(n_155)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_155),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_111),
.B(n_32),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_180),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_112),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_157),
.B(n_163),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_141),
.A2(n_34),
.B1(n_38),
.B2(n_37),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_159),
.Y(n_203)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

INVx4_ASAP7_75t_SL g161 ( 
.A(n_108),
.Y(n_161)
);

INVx4_ASAP7_75t_SL g218 ( 
.A(n_161),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_109),
.B(n_78),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_162),
.B(n_164),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_96),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_126),
.B(n_43),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_141),
.A2(n_37),
.B1(n_44),
.B2(n_94),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_166),
.Y(n_216)
);

AND2x2_ASAP7_75t_SL g167 ( 
.A(n_98),
.B(n_79),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_167),
.B(n_178),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_99),
.B(n_64),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_168),
.B(n_191),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_94),
.A2(n_44),
.B1(n_117),
.B2(n_118),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_169),
.A2(n_184),
.B1(n_185),
.B2(n_120),
.Y(n_198)
);

INVx6_ASAP7_75t_SL g172 ( 
.A(n_108),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_172),
.Y(n_207)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_95),
.Y(n_173)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_110),
.Y(n_175)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

OAI32xp33_ASAP7_75t_L g176 ( 
.A1(n_115),
.A2(n_55),
.A3(n_65),
.B1(n_47),
.B2(n_88),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_176),
.B(n_179),
.Y(n_224)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_114),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_100),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_101),
.B(n_35),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_125),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_181),
.B(n_40),
.Y(n_229)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_95),
.Y(n_182)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_105),
.B(n_35),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_39),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_117),
.A2(n_44),
.B1(n_45),
.B2(n_33),
.Y(n_184)
);

BUFx2_ASAP7_75t_SL g186 ( 
.A(n_135),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_186),
.Y(n_230)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_97),
.Y(n_187)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_138),
.Y(n_188)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_188),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_144),
.A2(n_103),
.B1(n_142),
.B2(n_130),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_97),
.B(n_89),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_106),
.B(n_89),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_192),
.B(n_121),
.Y(n_226)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_128),
.Y(n_193)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_110),
.Y(n_194)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_198),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_200),
.B(n_212),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_208),
.B(n_223),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_149),
.A2(n_123),
.B1(n_122),
.B2(n_136),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_210),
.A2(n_150),
.B1(n_194),
.B2(n_175),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_116),
.Y(n_212)
);

OAI32xp33_ASAP7_75t_L g214 ( 
.A1(n_156),
.A2(n_116),
.A3(n_104),
.B1(n_121),
.B2(n_137),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_226),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_148),
.A2(n_123),
.B1(n_122),
.B2(n_136),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_219),
.A2(n_222),
.B1(n_233),
.B2(n_155),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_167),
.A2(n_145),
.B1(n_162),
.B2(n_185),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_176),
.A2(n_40),
.B(n_104),
.Y(n_223)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_147),
.Y(n_227)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_227),
.Y(n_238)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_160),
.Y(n_228)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_228),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_232),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_181),
.B(n_107),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_155),
.A2(n_193),
.B1(n_189),
.B2(n_171),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_172),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_178),
.Y(n_252)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_158),
.Y(n_236)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

O2A1O1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_167),
.A2(n_65),
.B(n_107),
.C(n_137),
.Y(n_237)
);

OA21x2_ASAP7_75t_L g250 ( 
.A1(n_237),
.A2(n_150),
.B(n_188),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_241),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_195),
.B(n_158),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_242),
.B(n_260),
.Y(n_278)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_199),
.Y(n_243)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_243),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_209),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_244),
.B(n_252),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_197),
.A2(n_163),
.B1(n_189),
.B2(n_154),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_245),
.A2(n_271),
.B1(n_237),
.B2(n_225),
.Y(n_283)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_201),
.Y(n_247)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_247),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_230),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_248),
.B(n_249),
.Y(n_291)
);

NOR2x1_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_195),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_250),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_211),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_251),
.B(n_258),
.Y(n_305)
);

INVxp33_ASAP7_75t_L g302 ( 
.A(n_253),
.Y(n_302)
);

OAI32xp33_ASAP7_75t_L g254 ( 
.A1(n_224),
.A2(n_196),
.A3(n_223),
.B1(n_200),
.B2(n_214),
.Y(n_254)
);

AOI32xp33_ASAP7_75t_L g306 ( 
.A1(n_254),
.A2(n_5),
.A3(n_8),
.B1(n_9),
.B2(n_12),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_208),
.B(n_177),
.C(n_171),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_255),
.B(n_257),
.C(n_261),
.Y(n_303)
);

AO21x2_ASAP7_75t_L g256 ( 
.A1(n_197),
.A2(n_150),
.B(n_161),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_256),
.A2(n_266),
.B1(n_269),
.B2(n_204),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_217),
.B(n_206),
.C(n_212),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_183),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_199),
.B(n_170),
.Y(n_260)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_217),
.B(n_170),
.C(n_182),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_217),
.B(n_187),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_264),
.B(n_213),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_227),
.B(n_173),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_274),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_210),
.A2(n_151),
.B1(n_88),
.B2(n_81),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_207),
.B(n_152),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_267),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_203),
.A2(n_151),
.B1(n_81),
.B2(n_44),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_215),
.Y(n_270)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_203),
.A2(n_44),
.B1(n_2),
.B2(n_4),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_205),
.Y(n_272)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_205),
.Y(n_273)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_273),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_207),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_235),
.B(n_152),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_234),
.Y(n_293)
);

BUFx24_ASAP7_75t_L g276 ( 
.A(n_218),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_276),
.A2(n_218),
.B1(n_216),
.B2(n_215),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_268),
.A2(n_216),
.B1(n_228),
.B2(n_204),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_277),
.A2(n_281),
.B1(n_292),
.B2(n_250),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_280),
.A2(n_283),
.B1(n_285),
.B2(n_297),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_239),
.A2(n_220),
.B(n_236),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_284),
.B(n_288),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_268),
.A2(n_225),
.B1(n_220),
.B2(n_201),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_262),
.A2(n_218),
.B(n_234),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_264),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_249),
.A2(n_231),
.B(n_221),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_256),
.A2(n_202),
.B1(n_213),
.B2(n_221),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_293),
.B(n_299),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_295),
.B(n_250),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_245),
.A2(n_202),
.B1(n_231),
.B2(n_4),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_257),
.A2(n_1),
.B(n_2),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_242),
.B(n_1),
.Y(n_301)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_301),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_276),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_SL g316 ( 
.A(n_304),
.B(n_306),
.C(n_308),
.Y(n_316)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_238),
.Y(n_307)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_307),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_262),
.A2(n_5),
.B(n_8),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_254),
.B(n_5),
.Y(n_310)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_310),
.Y(n_326)
);

AO21x1_ASAP7_75t_L g356 ( 
.A1(n_311),
.A2(n_299),
.B(n_301),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_293),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_313),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_305),
.B(n_246),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_314),
.B(n_315),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_282),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_289),
.A2(n_256),
.B1(n_238),
.B2(n_263),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_317),
.A2(n_322),
.B1(n_336),
.B2(n_296),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_300),
.B(n_255),
.Y(n_320)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_320),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_265),
.Y(n_321)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_321),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_303),
.B(n_261),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_324),
.B(n_330),
.C(n_334),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_309),
.Y(n_325)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_325),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_310),
.A2(n_256),
.B1(n_253),
.B2(n_266),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_327),
.A2(n_281),
.B1(n_296),
.B2(n_292),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_294),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_328),
.B(n_339),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_282),
.Y(n_329)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_329),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_270),
.C(n_260),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_332),
.B(n_278),
.Y(n_340)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_294),
.Y(n_333)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_333),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_295),
.B(n_291),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_298),
.Y(n_335)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_335),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_289),
.A2(n_256),
.B1(n_240),
.B2(n_273),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_286),
.B(n_240),
.C(n_272),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_337),
.B(n_290),
.C(n_279),
.Y(n_359)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_298),
.Y(n_338)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_338),
.Y(n_354)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_307),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_340),
.B(n_351),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_322),
.A2(n_283),
.B1(n_296),
.B2(n_284),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_342),
.A2(n_357),
.B1(n_348),
.B2(n_349),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_346),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_348),
.A2(n_356),
.B1(n_336),
.B2(n_327),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_319),
.A2(n_288),
.B(n_277),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_349),
.B(n_361),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_324),
.B(n_308),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_334),
.B(n_300),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_353),
.B(n_355),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_330),
.B(n_278),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_326),
.A2(n_297),
.B1(n_285),
.B2(n_306),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_359),
.B(n_337),
.C(n_319),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_332),
.B(n_290),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_360),
.B(n_339),
.Y(n_381)
);

NOR3xp33_ASAP7_75t_SL g361 ( 
.A(n_326),
.B(n_279),
.C(n_276),
.Y(n_361)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_347),
.Y(n_364)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_364),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_365),
.B(n_366),
.C(n_371),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_350),
.B(n_313),
.C(n_323),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_350),
.B(n_323),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_369),
.B(n_374),
.Y(n_392)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_347),
.Y(n_370)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_370),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_355),
.B(n_325),
.C(n_318),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_343),
.B(n_287),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_373),
.B(n_376),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_353),
.B(n_331),
.Y(n_374)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_375),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_359),
.B(n_312),
.C(n_328),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_377),
.B(n_383),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_360),
.B(n_328),
.C(n_335),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_379),
.B(n_381),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_358),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_380),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_345),
.B(n_333),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g389 ( 
.A(n_382),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_341),
.A2(n_316),
.B1(n_302),
.B2(n_287),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_368),
.A2(n_374),
.B(n_379),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_384),
.B(n_390),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_365),
.A2(n_342),
.B(n_352),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_378),
.A2(n_352),
.B1(n_356),
.B2(n_357),
.Y(n_393)
);

OR2x2_ASAP7_75t_L g401 ( 
.A(n_393),
.B(n_396),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_376),
.B(n_344),
.Y(n_394)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_394),
.Y(n_402)
);

FAx1_ASAP7_75t_SL g396 ( 
.A(n_366),
.B(n_340),
.CI(n_351),
.CON(n_396),
.SN(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_371),
.B(n_363),
.Y(n_397)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_397),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_392),
.B(n_369),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_403),
.B(n_404),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_392),
.B(n_372),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_395),
.A2(n_362),
.B1(n_316),
.B2(n_354),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_406),
.A2(n_393),
.B1(n_390),
.B2(n_388),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_399),
.B(n_372),
.C(n_381),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_407),
.B(n_409),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_394),
.Y(n_408)
);

CKINVDCx14_ASAP7_75t_R g422 ( 
.A(n_408),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_399),
.B(n_367),
.C(n_354),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_391),
.B(n_386),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_410),
.A2(n_412),
.B1(n_389),
.B2(n_361),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_398),
.B(n_367),
.C(n_259),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_411),
.B(n_398),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_391),
.B(n_259),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_401),
.A2(n_395),
.B1(n_387),
.B2(n_385),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_413),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_414),
.B(n_400),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_416),
.B(n_404),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_401),
.A2(n_387),
.B1(n_388),
.B2(n_385),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_417),
.B(n_418),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_405),
.A2(n_389),
.B1(n_397),
.B2(n_384),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_419),
.B(n_422),
.Y(n_426)
);

NAND2xp33_ASAP7_75t_SL g421 ( 
.A(n_402),
.B(n_396),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_421),
.A2(n_411),
.B(n_409),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_423),
.B(n_425),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_426),
.B(n_427),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_418),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_415),
.B(n_400),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_429),
.B(n_430),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_423),
.B(n_413),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_432),
.B(n_414),
.Y(n_438)
);

A2O1A1Ixp33_ASAP7_75t_L g434 ( 
.A1(n_424),
.A2(n_420),
.B(n_407),
.C(n_417),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_434),
.A2(n_428),
.B(n_415),
.Y(n_436)
);

BUFx24_ASAP7_75t_SL g440 ( 
.A(n_436),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_433),
.B(n_431),
.C(n_435),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_437),
.A2(n_438),
.B(n_428),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_439),
.A2(n_416),
.B1(n_396),
.B2(n_403),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_441),
.A2(n_440),
.B(n_269),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_442),
.B(n_247),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_443),
.A2(n_8),
.B(n_439),
.Y(n_444)
);


endmodule