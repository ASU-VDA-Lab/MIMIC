module fake_jpeg_24401_n_255 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_255);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_255;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_42),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_0),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_31),
.Y(n_52)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_17),
.B(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_43),
.B(n_26),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_49),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_17),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_50),
.B(n_52),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_30),
.B1(n_22),
.B2(n_28),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_41),
.B1(n_47),
.B2(n_25),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_30),
.B1(n_22),
.B2(n_35),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_54),
.A2(n_61),
.B1(n_41),
.B2(n_18),
.Y(n_73)
);

CKINVDCx12_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_56),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_36),
.B(n_25),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_58),
.B(n_34),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_25),
.Y(n_60)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_22),
.B1(n_35),
.B2(n_24),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_43),
.B1(n_39),
.B2(n_18),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_62),
.A2(n_63),
.B1(n_67),
.B2(n_34),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_17),
.B1(n_29),
.B2(n_18),
.Y(n_63)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_32),
.Y(n_75)
);

AO22x1_ASAP7_75t_SL g67 ( 
.A1(n_41),
.A2(n_26),
.B1(n_32),
.B2(n_29),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_26),
.Y(n_86)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_70),
.Y(n_110)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_71),
.B(n_76),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_73),
.A2(n_64),
.B1(n_47),
.B2(n_24),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_50),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_99),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_75),
.Y(n_107)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_78),
.Y(n_120)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_67),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_41),
.B(n_29),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_95),
.C(n_74),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_32),
.Y(n_80)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_81),
.B(n_92),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_32),
.Y(n_82)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_84),
.A2(n_85),
.B1(n_87),
.B2(n_98),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_86),
.Y(n_121)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_33),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_88),
.B(n_96),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_89),
.A2(n_64),
.B1(n_20),
.B2(n_27),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_93),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_58),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_57),
.B(n_34),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_47),
.A2(n_23),
.B1(n_19),
.B2(n_21),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_62),
.B(n_21),
.Y(n_99)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_109),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_52),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_119),
.Y(n_144)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_95),
.B1(n_89),
.B2(n_77),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_112),
.A2(n_124),
.B1(n_20),
.B2(n_23),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_78),
.A2(n_55),
.B1(n_49),
.B2(n_68),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_113),
.A2(n_87),
.B1(n_91),
.B2(n_79),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_116),
.A2(n_71),
.B(n_90),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_26),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_83),
.A2(n_45),
.B1(n_44),
.B2(n_27),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_26),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_127),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_45),
.Y(n_127)
);

AND2x4_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_100),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_128),
.A2(n_102),
.B(n_108),
.Y(n_171)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_129),
.B(n_132),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_110),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_130),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_133),
.B1(n_134),
.B2(n_136),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_114),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_100),
.B1(n_91),
.B2(n_72),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_138),
.C(n_141),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_37),
.C(n_94),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_140),
.B(n_142),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_37),
.C(n_94),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_69),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_148),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_76),
.Y(n_145)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_70),
.Y(n_146)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_45),
.B1(n_44),
.B2(n_93),
.Y(n_147)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_105),
.A2(n_44),
.B(n_1),
.C(n_2),
.Y(n_149)
);

A2O1A1O1Ixp25_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_115),
.B(n_116),
.C(n_105),
.D(n_118),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_150)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_123),
.B(n_16),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_151),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_104),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_152),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_15),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_154),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_123),
.B(n_14),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_158),
.A2(n_13),
.B(n_7),
.C(n_8),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_117),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_161),
.A2(n_162),
.B(n_171),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_139),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_107),
.C(n_122),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_167),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_115),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_122),
.Y(n_170)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_170),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_128),
.A2(n_102),
.B(n_126),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_172),
.A2(n_175),
.B(n_6),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_135),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_173),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_129),
.A2(n_126),
.B(n_108),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_5),
.Y(n_178)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_178),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_176),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_179),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_168),
.B(n_152),
.Y(n_181)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_181),
.Y(n_211)
);

NOR3xp33_ASAP7_75t_SL g182 ( 
.A(n_168),
.B(n_130),
.C(n_148),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_171),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_177),
.A2(n_140),
.B1(n_143),
.B2(n_136),
.Y(n_183)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_183),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_141),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_197),
.Y(n_201)
);

A2O1A1O1Ixp25_ASAP7_75t_L g187 ( 
.A1(n_162),
.A2(n_137),
.B(n_133),
.C(n_149),
.D(n_154),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_158),
.C(n_167),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_150),
.Y(n_188)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

AO221x1_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_147),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_190),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_134),
.Y(n_192)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_192),
.Y(n_203)
);

OA21x2_ASAP7_75t_L g194 ( 
.A1(n_161),
.A2(n_6),
.B(n_7),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_194),
.A2(n_195),
.B(n_172),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_196),
.A2(n_169),
.B1(n_177),
.B2(n_163),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_6),
.Y(n_197)
);

MAJx2_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_11),
.C(n_9),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_178),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_205),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_200),
.A2(n_194),
.B(n_196),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_204),
.Y(n_224)
);

INVx13_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

BUFx24_ASAP7_75t_SL g218 ( 
.A(n_208),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_213),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_212),
.A2(n_189),
.B1(n_180),
.B2(n_164),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_214),
.A2(n_216),
.B1(n_217),
.B2(n_219),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_166),
.B1(n_191),
.B2(n_182),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_215),
.A2(n_225),
.B1(n_203),
.B2(n_210),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_206),
.A2(n_166),
.B1(n_170),
.B2(n_174),
.Y(n_217)
);

AOI21x1_ASAP7_75t_L g219 ( 
.A1(n_208),
.A2(n_198),
.B(n_194),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_213),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_205),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_212),
.A2(n_157),
.B(n_165),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_202),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_210),
.A2(n_174),
.B1(n_186),
.B2(n_160),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_201),
.C(n_204),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_229),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_203),
.Y(n_227)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_227),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_201),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_230),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_207),
.C(n_211),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_231),
.B(n_233),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_223),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_232),
.A2(n_235),
.B(n_209),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_199),
.C(n_187),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_227),
.A2(n_214),
.B(n_200),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_236),
.A2(n_239),
.B(n_184),
.Y(n_244)
);

AOI322xp5_ASAP7_75t_L g239 ( 
.A1(n_234),
.A2(n_185),
.A3(n_225),
.B1(n_184),
.B2(n_209),
.C1(n_156),
.C2(n_159),
.Y(n_239)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_241),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_239),
.C(n_242),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_228),
.C(n_232),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_9),
.C(n_10),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_156),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_246),
.A2(n_247),
.B(n_163),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_169),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_248),
.A2(n_250),
.B(n_243),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_249),
.B(n_251),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_245),
.A2(n_197),
.B(n_10),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_11),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_252),
.Y(n_255)
);


endmodule