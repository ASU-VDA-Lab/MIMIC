module fake_ariane_1946_n_1667 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1667);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1667;

wire n_913;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_146;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_149;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_150;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_145;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_888;
wire n_845;
wire n_1649;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_148;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_147;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_45),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_9),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_104),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_17),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_79),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_44),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_60),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_27),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_87),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_138),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_1),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_107),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_35),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_13),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_61),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_110),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_96),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_84),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_116),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_76),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_14),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_73),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_49),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_62),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_68),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_102),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_71),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_136),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_133),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_77),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_58),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_122),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_127),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_16),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_129),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_90),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_83),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_75),
.Y(n_187)
);

INVxp33_ASAP7_75t_R g188 ( 
.A(n_30),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_65),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_91),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_10),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_25),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_135),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_23),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_3),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_98),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_26),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_10),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_28),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_50),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_19),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_53),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_45),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_48),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_27),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_123),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_86),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_39),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_21),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_137),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_70),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_100),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_121),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_97),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g215 ( 
.A(n_113),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_19),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_63),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_52),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_143),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_67),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_33),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_89),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_126),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_4),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_106),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_33),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_57),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_94),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_34),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_29),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_43),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_95),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_35),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_120),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_31),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_41),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_43),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_78),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_93),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_39),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_41),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_54),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_34),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_24),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_66),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_49),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_44),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_56),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_85),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_117),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_72),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_112),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_11),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_18),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_36),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_32),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_59),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_82),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_114),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_9),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_69),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_125),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_15),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_141),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_14),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_132),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_111),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_52),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_37),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_99),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_48),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_6),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_55),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_37),
.Y(n_274)
);

BUFx8_ASAP7_75t_SL g275 ( 
.A(n_134),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_47),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_101),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_32),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_144),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_0),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_31),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_81),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_105),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_46),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_92),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_8),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_140),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_103),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_17),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_25),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_2),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_24),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_7),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_131),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_51),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_80),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_275),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_146),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_146),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_146),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_146),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_146),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_278),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_166),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_193),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_217),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_175),
.B(n_0),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_227),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_229),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_229),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_239),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_229),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_229),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_248),
.Y(n_314)
);

BUFx6f_ASAP7_75t_SL g315 ( 
.A(n_258),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_229),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_183),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_230),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_230),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_242),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_145),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_191),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_242),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_268),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_268),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_148),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_262),
.B(n_184),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_149),
.B(n_1),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_154),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_293),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_153),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_154),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_147),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_147),
.Y(n_334)
);

INVxp33_ASAP7_75t_SL g335 ( 
.A(n_192),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_194),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_195),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_167),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_167),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_236),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_259),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_291),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_150),
.B(n_155),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_259),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_158),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_197),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_171),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_260),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_198),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_199),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_201),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_200),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_179),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_204),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_159),
.B(n_2),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_202),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_208),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_209),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_203),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_157),
.B(n_3),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_216),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_205),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_218),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_221),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_224),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_233),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_212),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_235),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_219),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_240),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_253),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_310),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_329),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_303),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_329),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_310),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_367),
.B(n_163),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_304),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_305),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_310),
.Y(n_380)
);

NAND2x1_ASAP7_75t_L g381 ( 
.A(n_355),
.B(n_159),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_298),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_329),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_329),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_298),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_329),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_325),
.B(n_258),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_306),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_343),
.B(n_172),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_332),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_348),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_353),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_311),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_332),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_299),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_333),
.B(n_180),
.Y(n_396)
);

NAND2xp33_ASAP7_75t_SL g397 ( 
.A(n_330),
.B(n_226),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_332),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_332),
.Y(n_399)
);

OR2x6_ASAP7_75t_L g400 ( 
.A(n_330),
.B(n_256),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_332),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_297),
.Y(n_402)
);

AND2x4_ASAP7_75t_L g403 ( 
.A(n_333),
.B(n_185),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_321),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_299),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_308),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_300),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_334),
.B(n_185),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_340),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_300),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_342),
.B(n_188),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_301),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_314),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_334),
.B(n_159),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_317),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_369),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_301),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_302),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_302),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_309),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_315),
.B(n_258),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_R g422 ( 
.A(n_322),
.B(n_336),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_309),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_312),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_312),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_337),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_313),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_313),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_316),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_346),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_316),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_338),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_338),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_350),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_339),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_339),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_341),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_341),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_351),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_344),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_344),
.B(n_190),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_318),
.Y(n_442)
);

BUFx4f_ASAP7_75t_L g443 ( 
.A(n_442),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_400),
.B(n_315),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_400),
.B(n_315),
.Y(n_445)
);

INVx4_ASAP7_75t_L g446 ( 
.A(n_414),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_433),
.Y(n_447)
);

NAND2x1p5_ASAP7_75t_L g448 ( 
.A(n_387),
.B(n_325),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g449 ( 
.A(n_404),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_378),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_421),
.B(n_335),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_400),
.B(n_356),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_433),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_437),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_407),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_442),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_387),
.B(n_389),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_440),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_407),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_440),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_400),
.B(n_357),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_422),
.B(n_358),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_387),
.B(n_389),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_400),
.B(n_327),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_372),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_432),
.B(n_354),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_400),
.B(n_361),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_415),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_442),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_403),
.A2(n_307),
.B1(n_348),
.B2(n_359),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_372),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_391),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_377),
.Y(n_473)
);

INVx5_ASAP7_75t_L g474 ( 
.A(n_373),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g475 ( 
.A(n_391),
.B(n_363),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_422),
.B(n_364),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_442),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_430),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_428),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_403),
.B(n_408),
.Y(n_480)
);

NAND2xp33_ASAP7_75t_L g481 ( 
.A(n_434),
.B(n_215),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_409),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_376),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_374),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_428),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_428),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_376),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_432),
.B(n_362),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_432),
.B(n_370),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_421),
.A2(n_365),
.B1(n_360),
.B2(n_328),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_432),
.B(n_345),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_380),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_407),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g494 ( 
.A(n_374),
.B(n_326),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_381),
.B(n_331),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_426),
.Y(n_496)
);

INVx5_ASAP7_75t_L g497 ( 
.A(n_373),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_439),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_410),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_410),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g501 ( 
.A(n_416),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_380),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_403),
.A2(n_286),
.B1(n_284),
.B2(n_274),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_379),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_403),
.B(n_345),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_403),
.B(n_408),
.Y(n_506)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_392),
.B(n_388),
.Y(n_507)
);

OR2x6_ASAP7_75t_L g508 ( 
.A(n_392),
.B(n_347),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_410),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g510 ( 
.A(n_408),
.Y(n_510)
);

AOI22xp33_ASAP7_75t_L g511 ( 
.A1(n_408),
.A2(n_276),
.B1(n_280),
.B2(n_290),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_414),
.B(n_206),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_408),
.B(n_347),
.Y(n_513)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_393),
.B(n_352),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_381),
.B(n_438),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_414),
.B(n_349),
.Y(n_516)
);

INVx1_ASAP7_75t_SL g517 ( 
.A(n_406),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_397),
.B(n_349),
.Y(n_518)
);

NOR3xp33_ASAP7_75t_L g519 ( 
.A(n_402),
.B(n_244),
.C(n_160),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_414),
.B(n_210),
.Y(n_520)
);

AND2x6_ASAP7_75t_L g521 ( 
.A(n_414),
.B(n_212),
.Y(n_521)
);

BUFx10_ASAP7_75t_L g522 ( 
.A(n_413),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_418),
.Y(n_523)
);

NAND2xp33_ASAP7_75t_SL g524 ( 
.A(n_396),
.B(n_151),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_418),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_438),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_377),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_438),
.B(n_366),
.Y(n_528)
);

NOR3xp33_ASAP7_75t_L g529 ( 
.A(n_438),
.B(n_160),
.C(n_151),
.Y(n_529)
);

INVx5_ASAP7_75t_L g530 ( 
.A(n_373),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_411),
.Y(n_531)
);

NOR2x1p5_ASAP7_75t_L g532 ( 
.A(n_396),
.B(n_161),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_382),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_418),
.Y(n_534)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_411),
.B(n_366),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_382),
.Y(n_536)
);

BUFx8_ASAP7_75t_SL g537 ( 
.A(n_442),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_442),
.Y(n_538)
);

INVx4_ASAP7_75t_SL g539 ( 
.A(n_373),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_442),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_441),
.B(n_368),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_441),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_385),
.Y(n_543)
);

HB1xp67_ASAP7_75t_SL g544 ( 
.A(n_385),
.Y(n_544)
);

NAND2xp33_ASAP7_75t_L g545 ( 
.A(n_412),
.B(n_215),
.Y(n_545)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_373),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_395),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_435),
.B(n_214),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_395),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_435),
.B(n_368),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_435),
.B(n_371),
.Y(n_551)
);

INVx4_ASAP7_75t_SL g552 ( 
.A(n_373),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_436),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_436),
.B(n_371),
.Y(n_554)
);

AOI22x1_ASAP7_75t_L g555 ( 
.A1(n_436),
.A2(n_169),
.B1(n_161),
.B2(n_263),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_405),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_425),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_412),
.B(n_225),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_405),
.B(n_325),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_425),
.Y(n_560)
);

OR2x2_ASAP7_75t_L g561 ( 
.A(n_417),
.B(n_169),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_417),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_419),
.B(n_186),
.Y(n_563)
);

NOR3xp33_ASAP7_75t_L g564 ( 
.A(n_419),
.B(n_265),
.C(n_281),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_384),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_420),
.B(n_234),
.Y(n_566)
);

AND2x6_ASAP7_75t_L g567 ( 
.A(n_420),
.B(n_154),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_423),
.B(n_318),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_373),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_423),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_412),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_L g572 ( 
.A(n_412),
.B(n_215),
.Y(n_572)
);

INVxp67_ASAP7_75t_SL g573 ( 
.A(n_384),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_425),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_429),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_424),
.B(n_245),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_424),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_429),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_384),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_412),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_427),
.Y(n_581)
);

INVx4_ASAP7_75t_L g582 ( 
.A(n_375),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_429),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g584 ( 
.A(n_427),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_384),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_431),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_431),
.B(n_319),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_431),
.B(n_319),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_412),
.B(n_251),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_412),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_581),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_542),
.B(n_252),
.Y(n_592)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_475),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_553),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_542),
.B(n_261),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_452),
.B(n_263),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_446),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_473),
.B(n_285),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_461),
.B(n_265),
.Y(n_599)
);

BUFx5_ASAP7_75t_L g600 ( 
.A(n_521),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_527),
.B(n_386),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_581),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_507),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_467),
.B(n_269),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_560),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_560),
.Y(n_606)
);

OR2x6_ASAP7_75t_L g607 ( 
.A(n_508),
.B(n_320),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_527),
.B(n_386),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_444),
.B(n_445),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_510),
.A2(n_464),
.B1(n_457),
.B2(n_463),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_451),
.B(n_269),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_541),
.B(n_386),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_484),
.B(n_293),
.Y(n_613)
);

O2A1O1Ixp5_ASAP7_75t_L g614 ( 
.A1(n_495),
.A2(n_386),
.B(n_390),
.C(n_401),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_510),
.A2(n_272),
.B1(n_273),
.B2(n_295),
.Y(n_615)
);

BUFx5_ASAP7_75t_L g616 ( 
.A(n_521),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_466),
.B(n_152),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_562),
.A2(n_178),
.B1(n_181),
.B2(n_177),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_466),
.B(n_152),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_488),
.B(n_156),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_488),
.B(n_156),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_514),
.B(n_162),
.Y(n_622)
);

NOR2x1p5_ASAP7_75t_L g623 ( 
.A(n_468),
.B(n_271),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_494),
.B(n_271),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_489),
.B(n_162),
.Y(n_625)
);

OR2x2_ASAP7_75t_L g626 ( 
.A(n_472),
.B(n_272),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_498),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_449),
.B(n_273),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_489),
.B(n_390),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_468),
.B(n_293),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_462),
.B(n_281),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_515),
.B(n_491),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_462),
.B(n_476),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_562),
.A2(n_177),
.B1(n_176),
.B2(n_174),
.Y(n_634)
);

O2A1O1Ixp5_ASAP7_75t_L g635 ( 
.A1(n_443),
.A2(n_520),
.B(n_512),
.C(n_479),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_450),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_521),
.A2(n_270),
.B1(n_292),
.B2(n_289),
.Y(n_637)
);

O2A1O1Ixp33_ASAP7_75t_L g638 ( 
.A1(n_528),
.A2(n_324),
.B(n_323),
.C(n_320),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_508),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_490),
.B(n_164),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_550),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_446),
.B(n_164),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_551),
.Y(n_643)
);

OR2x6_ASAP7_75t_L g644 ( 
.A(n_508),
.B(n_323),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_446),
.B(n_165),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_584),
.B(n_165),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_465),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_471),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_456),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_476),
.B(n_289),
.Y(n_650)
);

OR2x6_ASAP7_75t_L g651 ( 
.A(n_508),
.B(n_478),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_544),
.B(n_292),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_448),
.B(n_168),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_518),
.B(n_295),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_481),
.A2(n_176),
.B1(n_173),
.B2(n_174),
.Y(n_655)
);

O2A1O1Ixp5_ASAP7_75t_L g656 ( 
.A1(n_443),
.A2(n_401),
.B(n_390),
.C(n_394),
.Y(n_656)
);

INVx8_ASAP7_75t_L g657 ( 
.A(n_521),
.Y(n_657)
);

NAND2xp33_ASAP7_75t_L g658 ( 
.A(n_456),
.B(n_469),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_478),
.B(n_324),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_491),
.B(n_390),
.Y(n_660)
);

INVxp33_ASAP7_75t_L g661 ( 
.A(n_535),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_516),
.B(n_401),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_516),
.B(n_401),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_481),
.A2(n_170),
.B1(n_173),
.B2(n_178),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_516),
.B(n_170),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_526),
.B(n_394),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_485),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_578),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_561),
.B(n_231),
.Y(n_669)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_482),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_483),
.Y(n_671)
);

O2A1O1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_480),
.A2(n_398),
.B(n_394),
.C(n_237),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_578),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_450),
.B(n_181),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_487),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_517),
.B(n_241),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_492),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_583),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_529),
.B(n_220),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_502),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_587),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_587),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_583),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_485),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_588),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_521),
.A2(n_270),
.B1(n_255),
.B2(n_247),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_486),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_506),
.B(n_220),
.Y(n_688)
);

INVx8_ASAP7_75t_L g689 ( 
.A(n_521),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_504),
.B(n_243),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_522),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_588),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_526),
.B(n_398),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_447),
.B(n_398),
.Y(n_694)
);

HB1xp67_ASAP7_75t_L g695 ( 
.A(n_498),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_532),
.B(n_246),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_453),
.B(n_215),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_512),
.A2(n_264),
.B1(n_266),
.B2(n_267),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_454),
.B(n_215),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_458),
.A2(n_254),
.B1(n_294),
.B2(n_264),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_486),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_460),
.B(n_215),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_559),
.B(n_266),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_505),
.B(n_267),
.Y(n_704)
);

OAI22xp5_ASAP7_75t_L g705 ( 
.A1(n_470),
.A2(n_294),
.B1(n_288),
.B2(n_287),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_455),
.Y(n_706)
);

OR2x6_ASAP7_75t_L g707 ( 
.A(n_513),
.B(n_154),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_522),
.B(n_496),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_554),
.B(n_277),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_SL g710 ( 
.A(n_522),
.B(n_270),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_455),
.Y(n_711)
);

OAI221xp5_ASAP7_75t_L g712 ( 
.A1(n_503),
.A2(n_277),
.B1(n_279),
.B2(n_282),
.C(n_283),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_533),
.B(n_215),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_519),
.B(n_279),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_554),
.B(n_282),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_559),
.B(n_283),
.Y(n_716)
);

NAND2xp33_ASAP7_75t_L g717 ( 
.A(n_456),
.B(n_287),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_501),
.B(n_288),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_568),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_554),
.B(n_182),
.Y(n_720)
);

O2A1O1Ixp33_ASAP7_75t_L g721 ( 
.A1(n_536),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_520),
.B(n_187),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_524),
.B(n_564),
.Y(n_723)
);

BUFx5_ASAP7_75t_L g724 ( 
.A(n_590),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_559),
.B(n_5),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_563),
.B(n_189),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_479),
.B(n_196),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_568),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_459),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_511),
.B(n_7),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_524),
.B(n_238),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_479),
.B(n_249),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_543),
.B(n_232),
.Y(n_733)
);

NAND2x1_ASAP7_75t_L g734 ( 
.A(n_538),
.B(n_399),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_547),
.B(n_549),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_555),
.B(n_228),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_556),
.Y(n_737)
);

A2O1A1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_566),
.A2(n_250),
.B(n_207),
.C(n_211),
.Y(n_738)
);

OR2x6_ASAP7_75t_L g739 ( 
.A(n_548),
.B(n_154),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_570),
.B(n_257),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_469),
.B(n_296),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_577),
.B(n_223),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_565),
.B(n_222),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_586),
.Y(n_744)
);

BUFx6f_ASAP7_75t_SL g745 ( 
.A(n_567),
.Y(n_745)
);

BUFx2_ASAP7_75t_R g746 ( 
.A(n_537),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_469),
.B(n_213),
.Y(n_747)
);

OAI221xp5_ASAP7_75t_L g748 ( 
.A1(n_576),
.A2(n_399),
.B1(n_383),
.B2(n_375),
.C(n_13),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_493),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_493),
.B(n_399),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_548),
.B(n_8),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_499),
.B(n_399),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_469),
.B(n_477),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_499),
.A2(n_399),
.B1(n_383),
.B2(n_375),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_573),
.A2(n_399),
.B(n_383),
.Y(n_755)
);

BUFx2_ASAP7_75t_L g756 ( 
.A(n_670),
.Y(n_756)
);

OAI21xp5_ASAP7_75t_L g757 ( 
.A1(n_614),
.A2(n_540),
.B(n_538),
.Y(n_757)
);

INVx4_ASAP7_75t_L g758 ( 
.A(n_657),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_627),
.Y(n_759)
);

AO32x1_ASAP7_75t_L g760 ( 
.A1(n_751),
.A2(n_557),
.A3(n_500),
.B1(n_534),
.B2(n_509),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_610),
.A2(n_565),
.B1(n_579),
.B2(n_540),
.Y(n_761)
);

O2A1O1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_596),
.A2(n_599),
.B(n_604),
.C(n_654),
.Y(n_762)
);

AO21x1_ASAP7_75t_L g763 ( 
.A1(n_609),
.A2(n_633),
.B(n_697),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_593),
.B(n_579),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_607),
.Y(n_765)
);

AOI21x1_ASAP7_75t_L g766 ( 
.A1(n_753),
.A2(n_589),
.B(n_558),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_737),
.Y(n_767)
);

AOI21xp33_ASAP7_75t_L g768 ( 
.A1(n_652),
.A2(n_589),
.B(n_558),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_632),
.A2(n_540),
.B(n_538),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_624),
.B(n_531),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_607),
.B(n_644),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_632),
.A2(n_582),
.B(n_546),
.Y(n_772)
);

BUFx2_ASAP7_75t_L g773 ( 
.A(n_607),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_706),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_666),
.A2(n_693),
.B(n_612),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_600),
.B(n_477),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_617),
.B(n_523),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_693),
.A2(n_582),
.B(n_546),
.Y(n_778)
);

A2O1A1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_631),
.A2(n_557),
.B(n_534),
.C(n_575),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_735),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_612),
.A2(n_569),
.B(n_585),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_711),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_603),
.B(n_531),
.Y(n_783)
);

NOR2x1p5_ASAP7_75t_SL g784 ( 
.A(n_724),
.B(n_525),
.Y(n_784)
);

A2O1A1Ixp33_ASAP7_75t_L g785 ( 
.A1(n_650),
.A2(n_575),
.B(n_574),
.C(n_525),
.Y(n_785)
);

NAND3xp33_ASAP7_75t_SL g786 ( 
.A(n_669),
.B(n_574),
.C(n_569),
.Y(n_786)
);

NOR3xp33_ASAP7_75t_L g787 ( 
.A(n_723),
.B(n_545),
.C(n_572),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_619),
.B(n_477),
.Y(n_788)
);

NAND2x1p5_ASAP7_75t_L g789 ( 
.A(n_597),
.B(n_477),
.Y(n_789)
);

A2O1A1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_611),
.A2(n_572),
.B(n_545),
.C(n_571),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_651),
.B(n_539),
.Y(n_791)
);

OAI22xp5_ASAP7_75t_L g792 ( 
.A1(n_735),
.A2(n_580),
.B1(n_571),
.B2(n_497),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_620),
.B(n_621),
.Y(n_793)
);

CKINVDCx10_ASAP7_75t_R g794 ( 
.A(n_651),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_629),
.A2(n_580),
.B(n_571),
.Y(n_795)
);

O2A1O1Ixp33_ASAP7_75t_L g796 ( 
.A1(n_625),
.A2(n_615),
.B(n_719),
.C(n_685),
.Y(n_796)
);

O2A1O1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_681),
.A2(n_11),
.B(n_12),
.C(n_15),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_647),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_729),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_592),
.B(n_537),
.Y(n_800)
);

NAND3xp33_ASAP7_75t_L g801 ( 
.A(n_676),
.B(n_580),
.C(n_571),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_601),
.A2(n_608),
.B(n_727),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_644),
.B(n_12),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_644),
.B(n_16),
.Y(n_804)
);

AOI21x1_ASAP7_75t_L g805 ( 
.A1(n_750),
.A2(n_552),
.B(n_539),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_592),
.B(n_552),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_600),
.B(n_616),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_597),
.B(n_552),
.Y(n_808)
);

OAI21x1_ASAP7_75t_L g809 ( 
.A1(n_750),
.A2(n_552),
.B(n_539),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_728),
.A2(n_474),
.B1(n_497),
.B2(n_530),
.Y(n_810)
);

O2A1O1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_682),
.A2(n_692),
.B(n_688),
.C(n_733),
.Y(n_811)
);

O2A1O1Ixp33_ASAP7_75t_SL g812 ( 
.A1(n_738),
.A2(n_736),
.B(n_642),
.C(n_645),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_648),
.Y(n_813)
);

OAI22xp5_ASAP7_75t_L g814 ( 
.A1(n_598),
.A2(n_474),
.B1(n_497),
.B2(n_530),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_657),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_732),
.A2(n_694),
.B(n_755),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_595),
.B(n_539),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_595),
.B(n_641),
.Y(n_818)
);

AO22x1_ASAP7_75t_L g819 ( 
.A1(n_636),
.A2(n_567),
.B1(n_530),
.B2(n_474),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_600),
.B(n_530),
.Y(n_820)
);

A2O1A1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_722),
.A2(n_375),
.B(n_383),
.C(n_399),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_643),
.B(n_567),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_730),
.A2(n_680),
.B1(n_677),
.B2(n_675),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_598),
.A2(n_375),
.B1(n_383),
.B2(n_21),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_749),
.Y(n_825)
);

O2A1O1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_733),
.A2(n_18),
.B(n_20),
.C(n_22),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_646),
.B(n_567),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_734),
.A2(n_383),
.B(n_375),
.Y(n_828)
);

INVx1_ASAP7_75t_SL g829 ( 
.A(n_708),
.Y(n_829)
);

AOI21x1_ASAP7_75t_L g830 ( 
.A1(n_752),
.A2(n_567),
.B(n_64),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_704),
.B(n_567),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_600),
.B(n_20),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_662),
.A2(n_139),
.B(n_130),
.Y(n_833)
);

NAND3xp33_ASAP7_75t_L g834 ( 
.A(n_618),
.B(n_22),
.C(n_23),
.Y(n_834)
);

AOI21x1_ASAP7_75t_L g835 ( 
.A1(n_752),
.A2(n_124),
.B(n_119),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_657),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_663),
.A2(n_658),
.B(n_702),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_663),
.A2(n_115),
.B(n_109),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_651),
.B(n_26),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_594),
.B(n_28),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_671),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_591),
.B(n_29),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_602),
.B(n_36),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_659),
.B(n_38),
.Y(n_844)
);

INVx11_ASAP7_75t_L g845 ( 
.A(n_746),
.Y(n_845)
);

A2O1A1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_635),
.A2(n_38),
.B(n_40),
.C(n_42),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_659),
.B(n_40),
.Y(n_847)
);

CKINVDCx10_ASAP7_75t_R g848 ( 
.A(n_695),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_699),
.A2(n_713),
.B(n_702),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_639),
.B(n_42),
.Y(n_850)
);

INVxp67_ASAP7_75t_L g851 ( 
.A(n_628),
.Y(n_851)
);

AO21x1_ASAP7_75t_L g852 ( 
.A1(n_713),
.A2(n_74),
.B(n_47),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_744),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_743),
.A2(n_46),
.B(n_50),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_605),
.Y(n_855)
);

A2O1A1Ixp33_ASAP7_75t_L g856 ( 
.A1(n_606),
.A2(n_54),
.B(n_55),
.C(n_668),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_673),
.Y(n_857)
);

OAI22xp5_ASAP7_75t_L g858 ( 
.A1(n_678),
.A2(n_683),
.B1(n_655),
.B2(n_664),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_726),
.B(n_630),
.Y(n_859)
);

BUFx2_ASAP7_75t_L g860 ( 
.A(n_718),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_689),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_740),
.A2(n_742),
.B(n_653),
.Y(n_862)
);

O2A1O1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_622),
.A2(n_674),
.B(n_712),
.C(n_665),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_703),
.A2(n_716),
.B1(n_637),
.B2(n_689),
.Y(n_864)
);

BUFx12f_ASAP7_75t_L g865 ( 
.A(n_691),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_613),
.B(n_661),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_690),
.B(n_725),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_600),
.B(n_616),
.Y(n_868)
);

OAI22xp5_ASAP7_75t_L g869 ( 
.A1(n_667),
.A2(n_684),
.B1(n_687),
.B2(n_701),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_667),
.A2(n_684),
.B(n_701),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_741),
.A2(n_747),
.B(n_672),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_L g872 ( 
.A1(n_715),
.A2(n_720),
.B(n_638),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_709),
.A2(n_689),
.B(n_649),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_634),
.B(n_716),
.Y(n_874)
);

BUFx12f_ASAP7_75t_L g875 ( 
.A(n_623),
.Y(n_875)
);

BUFx12f_ASAP7_75t_L g876 ( 
.A(n_696),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_703),
.B(n_710),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_714),
.B(n_698),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_640),
.B(n_679),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_724),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_686),
.B(n_700),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_705),
.B(n_626),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_649),
.A2(n_731),
.B(n_717),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_696),
.B(n_724),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_649),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_724),
.B(n_600),
.Y(n_886)
);

O2A1O1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_721),
.A2(n_748),
.B(n_739),
.C(n_707),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_745),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_739),
.B(n_707),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_616),
.A2(n_724),
.B1(n_754),
.B2(n_745),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_616),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_616),
.B(n_610),
.Y(n_892)
);

AOI22x1_ASAP7_75t_L g893 ( 
.A1(n_641),
.A2(n_643),
.B1(n_737),
.B2(n_453),
.Y(n_893)
);

CKINVDCx20_ASAP7_75t_R g894 ( 
.A(n_636),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_654),
.A2(n_599),
.B(n_604),
.C(n_596),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_654),
.B(n_596),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_610),
.B(n_600),
.Y(n_897)
);

NOR2xp67_ASAP7_75t_L g898 ( 
.A(n_636),
.B(n_504),
.Y(n_898)
);

AO21x1_ASAP7_75t_L g899 ( 
.A1(n_596),
.A2(n_604),
.B(n_599),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_654),
.B(n_542),
.Y(n_900)
);

OAI21xp33_ASAP7_75t_SL g901 ( 
.A1(n_610),
.A2(n_463),
.B(n_457),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_656),
.A2(n_614),
.B(n_750),
.Y(n_902)
);

O2A1O1Ixp5_ASAP7_75t_L g903 ( 
.A1(n_614),
.A2(n_381),
.B(n_635),
.C(n_736),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_654),
.B(n_542),
.Y(n_904)
);

A2O1A1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_654),
.A2(n_599),
.B(n_604),
.C(n_596),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_651),
.Y(n_906)
);

AO22x1_ASAP7_75t_L g907 ( 
.A1(n_636),
.A2(n_450),
.B1(n_305),
.B2(n_306),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_610),
.B(n_600),
.Y(n_908)
);

AOI21x1_ASAP7_75t_L g909 ( 
.A1(n_753),
.A2(n_752),
.B(n_750),
.Y(n_909)
);

O2A1O1Ixp33_ASAP7_75t_SL g910 ( 
.A1(n_632),
.A2(n_515),
.B(n_738),
.C(n_660),
.Y(n_910)
);

NAND3xp33_ASAP7_75t_SL g911 ( 
.A(n_596),
.B(n_604),
.C(n_599),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_737),
.Y(n_912)
);

BUFx8_ASAP7_75t_L g913 ( 
.A(n_708),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_737),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_737),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_596),
.A2(n_599),
.B1(n_604),
.B2(n_654),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_654),
.B(n_542),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_607),
.Y(n_918)
);

OAI21xp33_ASAP7_75t_L g919 ( 
.A1(n_596),
.A2(n_604),
.B(n_599),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_706),
.Y(n_920)
);

A2O1A1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_896),
.A2(n_762),
.B(n_916),
.C(n_905),
.Y(n_921)
);

AOI21xp33_ASAP7_75t_L g922 ( 
.A1(n_896),
.A2(n_919),
.B(n_895),
.Y(n_922)
);

AOI21x1_ASAP7_75t_L g923 ( 
.A1(n_802),
.A2(n_775),
.B(n_816),
.Y(n_923)
);

NOR2x1_ASAP7_75t_L g924 ( 
.A(n_894),
.B(n_898),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_911),
.B(n_900),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_770),
.B(n_866),
.Y(n_926)
);

AOI21x1_ASAP7_75t_L g927 ( 
.A1(n_892),
.A2(n_908),
.B(n_897),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_911),
.A2(n_917),
.B(n_904),
.Y(n_928)
);

AO31x2_ASAP7_75t_L g929 ( 
.A1(n_763),
.A2(n_899),
.A3(n_849),
.B(n_821),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_780),
.B(n_818),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_767),
.Y(n_931)
);

OAI21x1_ASAP7_75t_L g932 ( 
.A1(n_886),
.A2(n_909),
.B(n_868),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_862),
.A2(n_837),
.B(n_910),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_901),
.B(n_793),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_823),
.B(n_798),
.Y(n_935)
);

AO31x2_ASAP7_75t_L g936 ( 
.A1(n_852),
.A2(n_785),
.A3(n_779),
.B(n_871),
.Y(n_936)
);

A2O1A1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_881),
.A2(n_863),
.B(n_879),
.C(n_878),
.Y(n_937)
);

BUFx2_ASAP7_75t_L g938 ( 
.A(n_756),
.Y(n_938)
);

CKINVDCx20_ASAP7_75t_R g939 ( 
.A(n_913),
.Y(n_939)
);

OAI21x1_ASAP7_75t_L g940 ( 
.A1(n_807),
.A2(n_868),
.B(n_757),
.Y(n_940)
);

A2O1A1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_879),
.A2(n_811),
.B(n_887),
.C(n_867),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_813),
.Y(n_942)
);

OAI21xp33_ASAP7_75t_L g943 ( 
.A1(n_882),
.A2(n_840),
.B(n_874),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_874),
.A2(n_823),
.B1(n_912),
.B2(n_915),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_774),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_851),
.B(n_783),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_903),
.A2(n_769),
.B(n_772),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_791),
.Y(n_948)
);

AO31x2_ASAP7_75t_L g949 ( 
.A1(n_846),
.A2(n_806),
.A3(n_817),
.B(n_788),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_859),
.B(n_764),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_851),
.B(n_860),
.Y(n_951)
);

AOI21xp33_ASAP7_75t_L g952 ( 
.A1(n_826),
.A2(n_796),
.B(n_800),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_778),
.A2(n_786),
.B(n_908),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_829),
.B(n_773),
.Y(n_954)
);

AO31x2_ASAP7_75t_L g955 ( 
.A1(n_824),
.A2(n_777),
.A3(n_792),
.B(n_880),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_791),
.B(n_906),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_786),
.A2(n_892),
.B(n_897),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_907),
.B(n_759),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_841),
.B(n_914),
.Y(n_959)
);

AOI21x1_ASAP7_75t_L g960 ( 
.A1(n_831),
.A2(n_776),
.B(n_781),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_839),
.B(n_771),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_853),
.B(n_893),
.Y(n_962)
);

AO31x2_ASAP7_75t_L g963 ( 
.A1(n_790),
.A2(n_760),
.A3(n_795),
.B(n_858),
.Y(n_963)
);

AO31x2_ASAP7_75t_L g964 ( 
.A1(n_760),
.A2(n_761),
.A3(n_822),
.B(n_827),
.Y(n_964)
);

OAI21x1_ASAP7_75t_L g965 ( 
.A1(n_776),
.A2(n_903),
.B(n_766),
.Y(n_965)
);

NAND3xp33_ASAP7_75t_SL g966 ( 
.A(n_803),
.B(n_804),
.C(n_877),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_812),
.A2(n_870),
.B(n_820),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_787),
.A2(n_832),
.B(n_872),
.Y(n_968)
);

O2A1O1Ixp5_ASAP7_75t_L g969 ( 
.A1(n_883),
.A2(n_832),
.B(n_854),
.C(n_808),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_771),
.B(n_839),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_765),
.B(n_918),
.Y(n_971)
);

OAI21x1_ASAP7_75t_L g972 ( 
.A1(n_820),
.A2(n_891),
.B(n_835),
.Y(n_972)
);

OAI21xp5_ASAP7_75t_L g973 ( 
.A1(n_787),
.A2(n_838),
.B(n_833),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_782),
.Y(n_974)
);

AO31x2_ASAP7_75t_L g975 ( 
.A1(n_760),
.A2(n_843),
.A3(n_842),
.B(n_825),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_799),
.B(n_920),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_834),
.A2(n_850),
.B(n_840),
.C(n_884),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_836),
.Y(n_978)
);

OAI21x1_ASAP7_75t_L g979 ( 
.A1(n_830),
.A2(n_828),
.B(n_873),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_850),
.A2(n_768),
.B(n_764),
.C(n_803),
.Y(n_980)
);

INVx6_ASAP7_75t_L g981 ( 
.A(n_913),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_836),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_765),
.B(n_918),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_804),
.B(n_876),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_869),
.A2(n_847),
.B(n_844),
.Y(n_985)
);

AND2x2_ASAP7_75t_SL g986 ( 
.A(n_864),
.B(n_889),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_836),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_864),
.A2(n_856),
.B1(n_890),
.B2(n_789),
.Y(n_988)
);

NOR2x1_ASAP7_75t_L g989 ( 
.A(n_888),
.B(n_885),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_814),
.A2(n_801),
.B(n_810),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_789),
.A2(n_797),
.B1(n_855),
.B2(n_857),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_758),
.A2(n_815),
.B(n_819),
.Y(n_992)
);

AND3x4_ASAP7_75t_L g993 ( 
.A(n_848),
.B(n_845),
.C(n_794),
.Y(n_993)
);

BUFx6f_ASAP7_75t_SL g994 ( 
.A(n_836),
.Y(n_994)
);

O2A1O1Ixp5_ASAP7_75t_L g995 ( 
.A1(n_888),
.A2(n_784),
.B(n_758),
.C(n_865),
.Y(n_995)
);

OAI21x1_ASAP7_75t_L g996 ( 
.A1(n_861),
.A2(n_809),
.B(n_902),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_861),
.A2(n_875),
.B(n_895),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_861),
.B(n_896),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_895),
.A2(n_905),
.B(n_896),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_916),
.A2(n_896),
.B1(n_905),
.B2(n_895),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_770),
.B(n_593),
.Y(n_1001)
);

OAI21x1_ASAP7_75t_L g1002 ( 
.A1(n_809),
.A2(n_902),
.B(n_805),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_896),
.B(n_780),
.Y(n_1003)
);

AO31x2_ASAP7_75t_L g1004 ( 
.A1(n_763),
.A2(n_899),
.A3(n_849),
.B(n_821),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_774),
.Y(n_1005)
);

OAI21x1_ASAP7_75t_L g1006 ( 
.A1(n_809),
.A2(n_902),
.B(n_805),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_896),
.A2(n_762),
.B(n_916),
.C(n_905),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_896),
.B(n_780),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_791),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_895),
.A2(n_905),
.B(n_896),
.Y(n_1010)
);

OAI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_895),
.A2(n_905),
.B(n_896),
.Y(n_1011)
);

NAND2x1p5_ASAP7_75t_L g1012 ( 
.A(n_791),
.B(n_758),
.Y(n_1012)
);

OAI21x1_ASAP7_75t_L g1013 ( 
.A1(n_809),
.A2(n_902),
.B(n_805),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_767),
.Y(n_1014)
);

BUFx3_ASAP7_75t_L g1015 ( 
.A(n_894),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_895),
.A2(n_905),
.B(n_896),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_894),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_767),
.Y(n_1018)
);

BUFx3_ASAP7_75t_L g1019 ( 
.A(n_894),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_895),
.A2(n_905),
.B(n_896),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_896),
.B(n_780),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_895),
.A2(n_905),
.B(n_896),
.Y(n_1022)
);

BUFx4f_ASAP7_75t_L g1023 ( 
.A(n_876),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_770),
.B(n_593),
.Y(n_1024)
);

NAND2x1p5_ASAP7_75t_L g1025 ( 
.A(n_791),
.B(n_758),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_896),
.B(n_780),
.Y(n_1026)
);

AOI21x1_ASAP7_75t_SL g1027 ( 
.A1(n_867),
.A2(n_735),
.B(n_900),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_896),
.B(n_916),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_895),
.A2(n_905),
.B(n_896),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_895),
.A2(n_905),
.B(n_896),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_809),
.A2(n_902),
.B(n_805),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_916),
.B(n_896),
.Y(n_1032)
);

AO31x2_ASAP7_75t_L g1033 ( 
.A1(n_763),
.A2(n_899),
.A3(n_849),
.B(n_821),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_767),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_895),
.A2(n_905),
.B(n_896),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_896),
.B(n_780),
.Y(n_1036)
);

INVxp67_ASAP7_75t_SL g1037 ( 
.A(n_756),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_895),
.A2(n_905),
.B(n_896),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_896),
.B(n_780),
.Y(n_1039)
);

INVx2_ASAP7_75t_SL g1040 ( 
.A(n_848),
.Y(n_1040)
);

AND2x6_ASAP7_75t_L g1041 ( 
.A(n_836),
.B(n_861),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_895),
.A2(n_905),
.B(n_896),
.Y(n_1042)
);

NAND2x1_ASAP7_75t_L g1043 ( 
.A(n_758),
.B(n_815),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_770),
.B(n_593),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_896),
.B(n_780),
.Y(n_1045)
);

INVx4_ASAP7_75t_L g1046 ( 
.A(n_791),
.Y(n_1046)
);

AOI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_896),
.A2(n_916),
.B1(n_911),
.B2(n_919),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_896),
.A2(n_762),
.B(n_916),
.C(n_905),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_896),
.B(n_780),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_896),
.B(n_780),
.Y(n_1050)
);

AND2x2_ASAP7_75t_SL g1051 ( 
.A(n_896),
.B(n_451),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_895),
.A2(n_905),
.B(n_896),
.Y(n_1052)
);

AOI21xp33_ASAP7_75t_L g1053 ( 
.A1(n_896),
.A2(n_762),
.B(n_916),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_774),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_896),
.B(n_780),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_767),
.Y(n_1056)
);

AOI21x1_ASAP7_75t_L g1057 ( 
.A1(n_802),
.A2(n_775),
.B(n_816),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_896),
.B(n_780),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_926),
.B(n_1001),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_1023),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1028),
.B(n_1003),
.Y(n_1061)
);

OR2x6_ASAP7_75t_SL g1062 ( 
.A(n_1000),
.B(n_958),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_959),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_1051),
.B(n_1047),
.Y(n_1064)
);

INVx5_ASAP7_75t_L g1065 ( 
.A(n_1041),
.Y(n_1065)
);

AOI21xp33_ASAP7_75t_SL g1066 ( 
.A1(n_1032),
.A2(n_1053),
.B(n_1000),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1003),
.B(n_1036),
.Y(n_1067)
);

OAI321xp33_ASAP7_75t_L g1068 ( 
.A1(n_999),
.A2(n_1010),
.A3(n_1011),
.B1(n_1035),
.B2(n_1042),
.C(n_943),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1024),
.B(n_1044),
.Y(n_1069)
);

AOI22xp33_ASAP7_75t_L g1070 ( 
.A1(n_1053),
.A2(n_944),
.B1(n_1042),
.B2(n_1035),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_1016),
.A2(n_1022),
.B(n_1020),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1036),
.B(n_1039),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_939),
.Y(n_1073)
);

AOI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_966),
.A2(n_944),
.B1(n_925),
.B2(n_1026),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_948),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_946),
.B(n_951),
.Y(n_1076)
);

INVx1_ASAP7_75t_SL g1077 ( 
.A(n_1015),
.Y(n_1077)
);

OR2x6_ASAP7_75t_SL g1078 ( 
.A(n_1008),
.B(n_1021),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_1029),
.A2(n_1030),
.B(n_1038),
.Y(n_1079)
);

INVx2_ASAP7_75t_SL g1080 ( 
.A(n_981),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_961),
.B(n_954),
.Y(n_1081)
);

NAND2x1p5_ASAP7_75t_L g1082 ( 
.A(n_1046),
.B(n_948),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_1039),
.B(n_1055),
.Y(n_1083)
);

AOI21xp33_ASAP7_75t_L g1084 ( 
.A1(n_999),
.A2(n_1011),
.B(n_1010),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_931),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1055),
.B(n_1058),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_1037),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_1041),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_984),
.B(n_1045),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_1049),
.B(n_1050),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_942),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1052),
.A2(n_921),
.B(n_1007),
.Y(n_1092)
);

OR2x6_ASAP7_75t_L g1093 ( 
.A(n_981),
.B(n_1046),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1005),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1058),
.B(n_1048),
.Y(n_1095)
);

CKINVDCx11_ASAP7_75t_R g1096 ( 
.A(n_1017),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_998),
.B(n_922),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_930),
.B(n_934),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1054),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_922),
.A2(n_973),
.B(n_933),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_SL g1101 ( 
.A(n_993),
.B(n_1019),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_998),
.B(n_950),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_974),
.Y(n_1103)
);

INVx1_ASAP7_75t_SL g1104 ( 
.A(n_956),
.Y(n_1104)
);

BUFx4f_ASAP7_75t_SL g1105 ( 
.A(n_1040),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_1009),
.Y(n_1106)
);

AOI21xp33_ASAP7_75t_L g1107 ( 
.A1(n_934),
.A2(n_937),
.B(n_980),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_970),
.B(n_971),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_994),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_986),
.A2(n_935),
.B1(n_1034),
.B2(n_1056),
.Y(n_1110)
);

OR2x2_ASAP7_75t_L g1111 ( 
.A(n_983),
.B(n_1014),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_928),
.B(n_941),
.Y(n_1112)
);

OAI21xp33_ASAP7_75t_L g1113 ( 
.A1(n_977),
.A2(n_952),
.B(n_968),
.Y(n_1113)
);

AOI22xp33_ASAP7_75t_L g1114 ( 
.A1(n_935),
.A2(n_1018),
.B1(n_988),
.B2(n_968),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_997),
.B(n_924),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_989),
.B(n_982),
.Y(n_1116)
);

INVx2_ASAP7_75t_SL g1117 ( 
.A(n_1012),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_978),
.B(n_987),
.Y(n_1118)
);

INVx1_ASAP7_75t_SL g1119 ( 
.A(n_976),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_978),
.Y(n_1120)
);

CKINVDCx11_ASAP7_75t_R g1121 ( 
.A(n_978),
.Y(n_1121)
);

AOI222xp33_ASAP7_75t_L g1122 ( 
.A1(n_988),
.A2(n_985),
.B1(n_991),
.B2(n_962),
.C1(n_994),
.C2(n_1041),
.Y(n_1122)
);

NAND2xp33_ASAP7_75t_L g1123 ( 
.A(n_1041),
.B(n_987),
.Y(n_1123)
);

NAND2x1p5_ASAP7_75t_L g1124 ( 
.A(n_982),
.B(n_987),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_985),
.A2(n_952),
.B(n_957),
.C(n_962),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_1025),
.B(n_991),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_969),
.A2(n_953),
.B(n_967),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_990),
.A2(n_1043),
.B1(n_947),
.B2(n_927),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_992),
.B(n_940),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_995),
.B(n_929),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_965),
.A2(n_932),
.B1(n_972),
.B2(n_1027),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_996),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_929),
.B(n_1033),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1004),
.B(n_1033),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_1004),
.B(n_1033),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_949),
.B(n_955),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_979),
.A2(n_1013),
.B(n_1006),
.C(n_1002),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_SL g1138 ( 
.A1(n_963),
.A2(n_936),
.B1(n_955),
.B2(n_949),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_963),
.B(n_975),
.Y(n_1139)
);

NOR2xp67_ASAP7_75t_L g1140 ( 
.A(n_960),
.B(n_923),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_955),
.B(n_936),
.Y(n_1141)
);

INVxp67_ASAP7_75t_SL g1142 ( 
.A(n_1057),
.Y(n_1142)
);

NOR2xp67_ASAP7_75t_R g1143 ( 
.A(n_936),
.B(n_964),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_964),
.B(n_1031),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1028),
.A2(n_896),
.B1(n_916),
.B2(n_905),
.Y(n_1145)
);

INVx5_ASAP7_75t_L g1146 ( 
.A(n_1041),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_1028),
.B(n_1032),
.Y(n_1147)
);

OAI321xp33_ASAP7_75t_L g1148 ( 
.A1(n_999),
.A2(n_896),
.A3(n_916),
.B1(n_911),
.B2(n_919),
.C(n_905),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1028),
.B(n_1003),
.Y(n_1149)
);

AOI22xp33_ASAP7_75t_L g1150 ( 
.A1(n_1028),
.A2(n_943),
.B1(n_896),
.B2(n_1051),
.Y(n_1150)
);

INVx8_ASAP7_75t_L g1151 ( 
.A(n_994),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_1023),
.Y(n_1152)
);

BUFx3_ASAP7_75t_L g1153 ( 
.A(n_1023),
.Y(n_1153)
);

CKINVDCx8_ASAP7_75t_R g1154 ( 
.A(n_938),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_959),
.Y(n_1155)
);

AND2x2_ASAP7_75t_SL g1156 ( 
.A(n_1051),
.B(n_896),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1028),
.A2(n_896),
.B1(n_916),
.B2(n_1051),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1016),
.A2(n_1022),
.B(n_1020),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1028),
.B(n_1003),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_945),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_927),
.Y(n_1161)
);

NAND2xp33_ASAP7_75t_L g1162 ( 
.A(n_921),
.B(n_919),
.Y(n_1162)
);

INVx1_ASAP7_75t_SL g1163 ( 
.A(n_938),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1028),
.B(n_1003),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_945),
.Y(n_1165)
);

BUFx12f_ASAP7_75t_L g1166 ( 
.A(n_1040),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1028),
.B(n_916),
.Y(n_1167)
);

OAI21xp33_ASAP7_75t_SL g1168 ( 
.A1(n_1028),
.A2(n_916),
.B(n_896),
.Y(n_1168)
);

INVx1_ASAP7_75t_SL g1169 ( 
.A(n_938),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_959),
.Y(n_1170)
);

INVx3_ASAP7_75t_L g1171 ( 
.A(n_1041),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_945),
.Y(n_1172)
);

AOI21xp33_ASAP7_75t_SL g1173 ( 
.A1(n_1028),
.A2(n_450),
.B(n_636),
.Y(n_1173)
);

AOI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1028),
.A2(n_896),
.B1(n_916),
.B2(n_1051),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_959),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1028),
.B(n_1003),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_945),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1028),
.B(n_1003),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_927),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_1065),
.B(n_1146),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_1136),
.Y(n_1181)
);

INVx2_ASAP7_75t_SL g1182 ( 
.A(n_1065),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_1065),
.Y(n_1183)
);

CKINVDCx11_ASAP7_75t_R g1184 ( 
.A(n_1073),
.Y(n_1184)
);

AOI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1156),
.A2(n_1157),
.B1(n_1174),
.B2(n_1064),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1161),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1161),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1179),
.Y(n_1188)
);

NAND2x1p5_ASAP7_75t_L g1189 ( 
.A(n_1065),
.B(n_1146),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1168),
.A2(n_1145),
.B(n_1167),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_1136),
.Y(n_1191)
);

OR2x2_ASAP7_75t_L g1192 ( 
.A(n_1061),
.B(n_1149),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_1129),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1085),
.Y(n_1194)
);

OAI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1074),
.A2(n_1062),
.B1(n_1149),
.B2(n_1159),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1090),
.B(n_1061),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1156),
.A2(n_1150),
.B1(n_1110),
.B2(n_1070),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1091),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1179),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1133),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_1087),
.Y(n_1201)
);

AO21x1_ASAP7_75t_SL g1202 ( 
.A1(n_1070),
.A2(n_1084),
.B(n_1107),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1150),
.A2(n_1110),
.B1(n_1162),
.B2(n_1147),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1133),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1129),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1089),
.A2(n_1122),
.B1(n_1084),
.B2(n_1176),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1135),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1134),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1139),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1134),
.Y(n_1210)
);

OAI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1159),
.A2(n_1164),
.B1(n_1178),
.B2(n_1176),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1141),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1164),
.B(n_1178),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1103),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_1151),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_1151),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1111),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_1121),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_SL g1219 ( 
.A1(n_1092),
.A2(n_1066),
.B(n_1095),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_1088),
.Y(n_1220)
);

BUFx10_ASAP7_75t_L g1221 ( 
.A(n_1152),
.Y(n_1221)
);

BUFx2_ASAP7_75t_L g1222 ( 
.A(n_1130),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1098),
.A2(n_1059),
.B1(n_1069),
.B2(n_1095),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_1171),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1171),
.Y(n_1225)
);

NAND2x1p5_ASAP7_75t_L g1226 ( 
.A(n_1126),
.B(n_1097),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_SL g1227 ( 
.A1(n_1067),
.A2(n_1086),
.B1(n_1072),
.B2(n_1078),
.Y(n_1227)
);

OA21x2_ASAP7_75t_L g1228 ( 
.A1(n_1100),
.A2(n_1127),
.B(n_1079),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_SL g1229 ( 
.A1(n_1067),
.A2(n_1086),
.B1(n_1072),
.B2(n_1102),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1098),
.A2(n_1177),
.B1(n_1172),
.B2(n_1165),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1163),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1138),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1094),
.A2(n_1099),
.B1(n_1160),
.B2(n_1107),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_SL g1234 ( 
.A1(n_1092),
.A2(n_1112),
.B(n_1079),
.Y(n_1234)
);

OA21x2_ASAP7_75t_L g1235 ( 
.A1(n_1071),
.A2(n_1158),
.B(n_1125),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1142),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1142),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1114),
.B(n_1175),
.Y(n_1238)
);

OR2x2_ASAP7_75t_L g1239 ( 
.A(n_1063),
.B(n_1155),
.Y(n_1239)
);

INVx3_ASAP7_75t_L g1240 ( 
.A(n_1132),
.Y(n_1240)
);

OAI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1148),
.A2(n_1068),
.B1(n_1101),
.B2(n_1170),
.Y(n_1241)
);

AO21x2_ASAP7_75t_L g1242 ( 
.A1(n_1140),
.A2(n_1144),
.B(n_1137),
.Y(n_1242)
);

BUFx3_ASAP7_75t_L g1243 ( 
.A(n_1151),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1169),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1119),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_1132),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1076),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1083),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_SL g1249 ( 
.A1(n_1112),
.A2(n_1108),
.B1(n_1115),
.B2(n_1104),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1113),
.A2(n_1114),
.B1(n_1081),
.B2(n_1080),
.Y(n_1250)
);

OAI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1077),
.A2(n_1093),
.B1(n_1173),
.B2(n_1154),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1120),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_SL g1253 ( 
.A1(n_1123),
.A2(n_1117),
.B1(n_1128),
.B2(n_1106),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1060),
.A2(n_1153),
.B1(n_1082),
.B2(n_1109),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1132),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1144),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1143),
.Y(n_1257)
);

HB1xp67_ASAP7_75t_L g1258 ( 
.A(n_1075),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1131),
.A2(n_1124),
.B(n_1116),
.Y(n_1259)
);

BUFx12f_ASAP7_75t_L g1260 ( 
.A(n_1096),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1118),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1124),
.Y(n_1262)
);

BUFx2_ASAP7_75t_R g1263 ( 
.A(n_1105),
.Y(n_1263)
);

BUFx2_ASAP7_75t_R g1264 ( 
.A(n_1105),
.Y(n_1264)
);

CKINVDCx11_ASAP7_75t_R g1265 ( 
.A(n_1166),
.Y(n_1265)
);

AOI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1156),
.A2(n_896),
.B1(n_1028),
.B2(n_1051),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1161),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1070),
.B(n_1147),
.Y(n_1268)
);

BUFx6f_ASAP7_75t_SL g1269 ( 
.A(n_1060),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1090),
.B(n_1061),
.Y(n_1270)
);

CKINVDCx6p67_ASAP7_75t_R g1271 ( 
.A(n_1060),
.Y(n_1271)
);

BUFx2_ASAP7_75t_R g1272 ( 
.A(n_1152),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1161),
.Y(n_1273)
);

INVxp67_ASAP7_75t_SL g1274 ( 
.A(n_1098),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1161),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1085),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1085),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1085),
.Y(n_1278)
);

INVx3_ASAP7_75t_L g1279 ( 
.A(n_1129),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1161),
.Y(n_1280)
);

OAI22xp33_ASAP7_75t_SL g1281 ( 
.A1(n_1062),
.A2(n_1064),
.B1(n_1078),
.B2(n_451),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1193),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_1184),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1257),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1190),
.A2(n_1266),
.B(n_1203),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_1201),
.Y(n_1286)
);

NAND3xp33_ASAP7_75t_L g1287 ( 
.A(n_1185),
.B(n_1268),
.C(n_1197),
.Y(n_1287)
);

AO21x1_ASAP7_75t_SL g1288 ( 
.A1(n_1257),
.A2(n_1256),
.B(n_1187),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1222),
.B(n_1209),
.Y(n_1289)
);

BUFx2_ASAP7_75t_L g1290 ( 
.A(n_1193),
.Y(n_1290)
);

INVxp67_ASAP7_75t_L g1291 ( 
.A(n_1231),
.Y(n_1291)
);

OA21x2_ASAP7_75t_L g1292 ( 
.A1(n_1234),
.A2(n_1237),
.B(n_1236),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1222),
.B(n_1209),
.Y(n_1293)
);

CKINVDCx14_ASAP7_75t_R g1294 ( 
.A(n_1184),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1268),
.B(n_1232),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1193),
.B(n_1205),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1232),
.B(n_1207),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1195),
.A2(n_1227),
.B1(n_1281),
.B2(n_1202),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1238),
.B(n_1181),
.Y(n_1299)
);

OA21x2_ASAP7_75t_L g1300 ( 
.A1(n_1237),
.A2(n_1256),
.B(n_1219),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1235),
.A2(n_1228),
.B(n_1259),
.Y(n_1301)
);

OR2x6_ASAP7_75t_L g1302 ( 
.A(n_1181),
.B(n_1191),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1238),
.B(n_1191),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1200),
.Y(n_1304)
);

OR2x2_ASAP7_75t_L g1305 ( 
.A(n_1204),
.B(n_1208),
.Y(n_1305)
);

AOI21xp33_ASAP7_75t_SL g1306 ( 
.A1(n_1211),
.A2(n_1241),
.B(n_1251),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1204),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1208),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1210),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1210),
.Y(n_1310)
);

BUFx3_ASAP7_75t_L g1311 ( 
.A(n_1180),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1248),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_1244),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1186),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1186),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1280),
.Y(n_1316)
);

OR2x2_ASAP7_75t_L g1317 ( 
.A(n_1187),
.B(n_1188),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1188),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1199),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1235),
.A2(n_1228),
.B(n_1255),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1202),
.B(n_1279),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1280),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1267),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1252),
.Y(n_1324)
);

OR2x2_ASAP7_75t_L g1325 ( 
.A(n_1273),
.B(n_1275),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1273),
.Y(n_1326)
);

INVx4_ASAP7_75t_SL g1327 ( 
.A(n_1183),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1275),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_1239),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1235),
.A2(n_1228),
.B(n_1246),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1239),
.Y(n_1331)
);

CKINVDCx16_ASAP7_75t_R g1332 ( 
.A(n_1218),
.Y(n_1332)
);

AO21x1_ASAP7_75t_SL g1333 ( 
.A1(n_1206),
.A2(n_1212),
.B(n_1250),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1235),
.A2(n_1240),
.B(n_1246),
.Y(n_1334)
);

INVxp67_ASAP7_75t_L g1335 ( 
.A(n_1217),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1274),
.B(n_1229),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1212),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1194),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1278),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1198),
.B(n_1277),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1242),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1276),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1242),
.Y(n_1343)
);

AO21x2_ASAP7_75t_L g1344 ( 
.A1(n_1242),
.A2(n_1214),
.B(n_1213),
.Y(n_1344)
);

INVx3_ASAP7_75t_L g1345 ( 
.A(n_1220),
.Y(n_1345)
);

AO21x2_ASAP7_75t_L g1346 ( 
.A1(n_1196),
.A2(n_1270),
.B(n_1245),
.Y(n_1346)
);

OA21x2_ASAP7_75t_L g1347 ( 
.A1(n_1233),
.A2(n_1230),
.B(n_1223),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1300),
.B(n_1247),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1300),
.B(n_1226),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1329),
.B(n_1192),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1289),
.B(n_1192),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1293),
.B(n_1249),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1292),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1299),
.B(n_1224),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1299),
.B(n_1224),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1292),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1292),
.Y(n_1357)
);

INVxp67_ASAP7_75t_SL g1358 ( 
.A(n_1292),
.Y(n_1358)
);

AOI31xp33_ASAP7_75t_L g1359 ( 
.A1(n_1298),
.A2(n_1253),
.A3(n_1189),
.B(n_1182),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1286),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1346),
.B(n_1258),
.Y(n_1361)
);

NOR2x1p5_ASAP7_75t_L g1362 ( 
.A(n_1311),
.B(n_1260),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1346),
.B(n_1262),
.Y(n_1363)
);

AOI21xp33_ASAP7_75t_SL g1364 ( 
.A1(n_1332),
.A2(n_1254),
.B(n_1260),
.Y(n_1364)
);

INVx3_ASAP7_75t_L g1365 ( 
.A(n_1334),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1303),
.B(n_1225),
.Y(n_1366)
);

BUFx3_ASAP7_75t_L g1367 ( 
.A(n_1302),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1284),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1317),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1346),
.B(n_1262),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1331),
.B(n_1303),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1301),
.B(n_1320),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1346),
.B(n_1261),
.Y(n_1373)
);

INVx4_ASAP7_75t_L g1374 ( 
.A(n_1327),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1314),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1314),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1320),
.B(n_1330),
.Y(n_1377)
);

AND2x2_ASAP7_75t_SL g1378 ( 
.A(n_1290),
.B(n_1183),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1302),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1317),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1315),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1315),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1316),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1325),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1325),
.B(n_1218),
.Y(n_1385)
);

AOI221xp5_ASAP7_75t_L g1386 ( 
.A1(n_1348),
.A2(n_1306),
.B1(n_1287),
.B2(n_1285),
.C(n_1295),
.Y(n_1386)
);

OAI221xp5_ASAP7_75t_L g1387 ( 
.A1(n_1359),
.A2(n_1285),
.B1(n_1287),
.B2(n_1336),
.C(n_1295),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1351),
.B(n_1313),
.Y(n_1388)
);

NAND3xp33_ASAP7_75t_L g1389 ( 
.A(n_1361),
.B(n_1312),
.C(n_1336),
.Y(n_1389)
);

OAI221xp5_ASAP7_75t_L g1390 ( 
.A1(n_1359),
.A2(n_1361),
.B1(n_1373),
.B2(n_1370),
.C(n_1363),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1360),
.B(n_1369),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1360),
.B(n_1291),
.Y(n_1392)
);

NAND3xp33_ASAP7_75t_L g1393 ( 
.A(n_1353),
.B(n_1324),
.C(n_1319),
.Y(n_1393)
);

NAND3xp33_ASAP7_75t_L g1394 ( 
.A(n_1353),
.B(n_1328),
.C(n_1318),
.Y(n_1394)
);

NAND4xp25_ASAP7_75t_L g1395 ( 
.A(n_1368),
.B(n_1321),
.C(n_1323),
.D(n_1318),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1369),
.B(n_1340),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_SL g1397 ( 
.A(n_1364),
.B(n_1332),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1380),
.B(n_1340),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1385),
.A2(n_1294),
.B1(n_1302),
.B2(n_1218),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_SL g1400 ( 
.A(n_1364),
.B(n_1283),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1354),
.B(n_1288),
.Y(n_1401)
);

AND2x2_ASAP7_75t_SL g1402 ( 
.A(n_1378),
.B(n_1296),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1350),
.B(n_1218),
.Y(n_1403)
);

OAI21xp5_ASAP7_75t_SL g1404 ( 
.A1(n_1356),
.A2(n_1357),
.B(n_1368),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1380),
.B(n_1335),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1352),
.A2(n_1333),
.B1(n_1347),
.B2(n_1297),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_1350),
.B(n_1271),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1355),
.B(n_1288),
.Y(n_1408)
);

OAI221xp5_ASAP7_75t_SL g1409 ( 
.A1(n_1358),
.A2(n_1342),
.B1(n_1339),
.B2(n_1338),
.C(n_1310),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1384),
.B(n_1344),
.Y(n_1410)
);

OAI21xp5_ASAP7_75t_SL g1411 ( 
.A1(n_1356),
.A2(n_1297),
.B(n_1319),
.Y(n_1411)
);

OAI221xp5_ASAP7_75t_L g1412 ( 
.A1(n_1373),
.A2(n_1338),
.B1(n_1339),
.B2(n_1342),
.C(n_1322),
.Y(n_1412)
);

NAND3xp33_ASAP7_75t_L g1413 ( 
.A(n_1357),
.B(n_1358),
.C(n_1348),
.Y(n_1413)
);

AOI221xp5_ASAP7_75t_L g1414 ( 
.A1(n_1348),
.A2(n_1304),
.B1(n_1310),
.B2(n_1308),
.C(n_1307),
.Y(n_1414)
);

OAI21xp5_ASAP7_75t_SL g1415 ( 
.A1(n_1368),
.A2(n_1322),
.B(n_1323),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1355),
.B(n_1282),
.Y(n_1416)
);

OAI221xp5_ASAP7_75t_SL g1417 ( 
.A1(n_1349),
.A2(n_1307),
.B1(n_1308),
.B2(n_1305),
.C(n_1328),
.Y(n_1417)
);

OAI221xp5_ASAP7_75t_L g1418 ( 
.A1(n_1363),
.A2(n_1326),
.B1(n_1337),
.B2(n_1343),
.C(n_1341),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1366),
.B(n_1282),
.Y(n_1419)
);

NAND3xp33_ASAP7_75t_L g1420 ( 
.A(n_1372),
.B(n_1326),
.C(n_1305),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1350),
.B(n_1309),
.Y(n_1421)
);

NAND3xp33_ASAP7_75t_L g1422 ( 
.A(n_1372),
.B(n_1341),
.C(n_1337),
.Y(n_1422)
);

OAI221xp5_ASAP7_75t_SL g1423 ( 
.A1(n_1349),
.A2(n_1341),
.B1(n_1343),
.B2(n_1271),
.C(n_1333),
.Y(n_1423)
);

NOR3xp33_ASAP7_75t_L g1424 ( 
.A(n_1365),
.B(n_1341),
.C(n_1345),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1422),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1391),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1414),
.B(n_1375),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1401),
.B(n_1367),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1421),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1412),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1394),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1420),
.B(n_1375),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1394),
.Y(n_1433)
);

INVxp33_ASAP7_75t_L g1434 ( 
.A(n_1403),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_SL g1435 ( 
.A(n_1387),
.B(n_1374),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1400),
.B(n_1265),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1396),
.B(n_1371),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1398),
.B(n_1371),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1388),
.B(n_1371),
.Y(n_1439)
);

AOI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1386),
.A2(n_1406),
.B1(n_1390),
.B2(n_1352),
.Y(n_1440)
);

BUFx3_ASAP7_75t_L g1441 ( 
.A(n_1402),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1410),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1420),
.B(n_1376),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1401),
.B(n_1377),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1408),
.B(n_1377),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1415),
.B(n_1376),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1408),
.B(n_1377),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1402),
.B(n_1379),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1402),
.B(n_1379),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1411),
.B(n_1381),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1405),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1393),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1393),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1413),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1422),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1413),
.B(n_1381),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1418),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1404),
.B(n_1382),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1444),
.B(n_1416),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1430),
.B(n_1431),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1431),
.B(n_1382),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1441),
.B(n_1424),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1432),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1425),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1425),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1432),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1444),
.B(n_1419),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1445),
.B(n_1419),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1433),
.B(n_1383),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1441),
.B(n_1362),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1443),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1443),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1445),
.B(n_1447),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1425),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1456),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1455),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1456),
.Y(n_1477)
);

NOR3xp33_ASAP7_75t_L g1478 ( 
.A(n_1454),
.B(n_1409),
.C(n_1417),
.Y(n_1478)
);

AOI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1440),
.A2(n_1352),
.B1(n_1389),
.B2(n_1407),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1429),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1429),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1427),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1430),
.B(n_1433),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1427),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1437),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1455),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1437),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1452),
.B(n_1383),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1438),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1438),
.Y(n_1490)
);

INVx2_ASAP7_75t_SL g1491 ( 
.A(n_1441),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1461),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1461),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1460),
.B(n_1452),
.Y(n_1494)
);

A2O1A1Ixp33_ASAP7_75t_L g1495 ( 
.A1(n_1478),
.A2(n_1440),
.B(n_1457),
.C(n_1435),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1473),
.B(n_1454),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1478),
.B(n_1457),
.Y(n_1497)
);

INVxp67_ASAP7_75t_L g1498 ( 
.A(n_1460),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1482),
.B(n_1453),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1469),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1473),
.B(n_1428),
.Y(n_1501)
);

INVxp33_ASAP7_75t_L g1502 ( 
.A(n_1483),
.Y(n_1502)
);

OR3x2_ASAP7_75t_L g1503 ( 
.A(n_1483),
.B(n_1484),
.C(n_1482),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1469),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1488),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1459),
.B(n_1428),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1459),
.B(n_1428),
.Y(n_1507)
);

NOR2x1_ASAP7_75t_L g1508 ( 
.A(n_1464),
.B(n_1436),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1488),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1464),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1485),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1485),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1487),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1487),
.B(n_1439),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1464),
.Y(n_1515)
);

INVxp33_ASAP7_75t_L g1516 ( 
.A(n_1470),
.Y(n_1516)
);

AOI21x1_ASAP7_75t_SL g1517 ( 
.A1(n_1462),
.A2(n_1470),
.B(n_1458),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1489),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1489),
.Y(n_1519)
);

OAI21xp33_ASAP7_75t_L g1520 ( 
.A1(n_1484),
.A2(n_1455),
.B(n_1453),
.Y(n_1520)
);

INVx3_ASAP7_75t_L g1521 ( 
.A(n_1470),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1490),
.B(n_1450),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1490),
.B(n_1450),
.Y(n_1523)
);

NOR2x1_ASAP7_75t_SL g1524 ( 
.A(n_1491),
.B(n_1448),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1463),
.B(n_1446),
.Y(n_1525)
);

OAI32xp33_ASAP7_75t_L g1526 ( 
.A1(n_1465),
.A2(n_1458),
.A3(n_1446),
.B1(n_1395),
.B2(n_1434),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1465),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1480),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1480),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1481),
.Y(n_1530)
);

AO22x1_ASAP7_75t_L g1531 ( 
.A1(n_1470),
.A2(n_1448),
.B1(n_1449),
.B2(n_1428),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1463),
.B(n_1451),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1466),
.B(n_1451),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1465),
.B(n_1426),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1528),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1494),
.B(n_1466),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1503),
.Y(n_1537)
);

INVxp67_ASAP7_75t_L g1538 ( 
.A(n_1508),
.Y(n_1538)
);

CKINVDCx16_ASAP7_75t_R g1539 ( 
.A(n_1497),
.Y(n_1539)
);

INVx1_ASAP7_75t_SL g1540 ( 
.A(n_1494),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1524),
.B(n_1491),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1521),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1529),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1530),
.Y(n_1544)
);

INVx1_ASAP7_75t_SL g1545 ( 
.A(n_1521),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1499),
.B(n_1471),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1514),
.B(n_1471),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1521),
.B(n_1491),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1503),
.A2(n_1495),
.B1(n_1479),
.B2(n_1516),
.Y(n_1549)
);

CKINVDCx16_ASAP7_75t_R g1550 ( 
.A(n_1496),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1511),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1506),
.B(n_1507),
.Y(n_1552)
);

INVx1_ASAP7_75t_SL g1553 ( 
.A(n_1502),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1498),
.B(n_1472),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1502),
.B(n_1520),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1512),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1506),
.B(n_1459),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1513),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1495),
.B(n_1472),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1516),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1496),
.B(n_1475),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1507),
.B(n_1467),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1510),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1518),
.Y(n_1564)
);

INVx2_ASAP7_75t_SL g1565 ( 
.A(n_1531),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1510),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1519),
.Y(n_1567)
);

INVx2_ASAP7_75t_SL g1568 ( 
.A(n_1534),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1515),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1532),
.Y(n_1570)
);

A2O1A1Ixp33_ASAP7_75t_L g1571 ( 
.A1(n_1537),
.A2(n_1526),
.B(n_1479),
.C(n_1486),
.Y(n_1571)
);

NOR3xp33_ASAP7_75t_L g1572 ( 
.A(n_1539),
.B(n_1476),
.C(n_1474),
.Y(n_1572)
);

AOI221xp5_ASAP7_75t_L g1573 ( 
.A1(n_1537),
.A2(n_1476),
.B1(n_1486),
.B2(n_1474),
.C(n_1525),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1535),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_SL g1575 ( 
.A(n_1549),
.B(n_1474),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1535),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1543),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1550),
.B(n_1522),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1542),
.Y(n_1579)
);

INVx2_ASAP7_75t_SL g1580 ( 
.A(n_1542),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1552),
.Y(n_1581)
);

NAND4xp25_ASAP7_75t_L g1582 ( 
.A(n_1560),
.B(n_1545),
.C(n_1555),
.D(n_1553),
.Y(n_1582)
);

OA21x2_ASAP7_75t_L g1583 ( 
.A1(n_1559),
.A2(n_1486),
.B(n_1476),
.Y(n_1583)
);

OAI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1538),
.A2(n_1477),
.B(n_1475),
.Y(n_1584)
);

AOI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1565),
.A2(n_1477),
.B(n_1533),
.Y(n_1585)
);

AOI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1565),
.A2(n_1435),
.B1(n_1527),
.B2(n_1515),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_L g1587 ( 
.A(n_1540),
.B(n_1265),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1552),
.Y(n_1588)
);

OAI21x1_ASAP7_75t_SL g1589 ( 
.A1(n_1567),
.A2(n_1517),
.B(n_1522),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1543),
.Y(n_1590)
);

OAI221xp5_ASAP7_75t_L g1591 ( 
.A1(n_1561),
.A2(n_1523),
.B1(n_1527),
.B2(n_1500),
.C(n_1509),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1544),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1544),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1570),
.B(n_1492),
.Y(n_1594)
);

A2O1A1Ixp33_ASAP7_75t_L g1595 ( 
.A1(n_1541),
.A2(n_1523),
.B(n_1462),
.C(n_1423),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1572),
.B(n_1570),
.Y(n_1596)
);

BUFx2_ASAP7_75t_L g1597 ( 
.A(n_1579),
.Y(n_1597)
);

AOI21xp33_ASAP7_75t_SL g1598 ( 
.A1(n_1572),
.A2(n_1541),
.B(n_1567),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1578),
.B(n_1568),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1580),
.B(n_1568),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1574),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_L g1602 ( 
.A(n_1587),
.B(n_1552),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1581),
.B(n_1557),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1576),
.Y(n_1604)
);

NAND3xp33_ASAP7_75t_L g1605 ( 
.A(n_1571),
.B(n_1548),
.C(n_1556),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1588),
.B(n_1557),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1587),
.B(n_1548),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1584),
.B(n_1562),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1577),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1583),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1585),
.B(n_1562),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1590),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1592),
.B(n_1548),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1582),
.B(n_1551),
.Y(n_1614)
);

OAI221xp5_ASAP7_75t_L g1615 ( 
.A1(n_1605),
.A2(n_1571),
.B1(n_1575),
.B2(n_1610),
.C(n_1595),
.Y(n_1615)
);

NAND4xp25_ASAP7_75t_L g1616 ( 
.A(n_1602),
.B(n_1595),
.C(n_1593),
.D(n_1591),
.Y(n_1616)
);

AOI221xp5_ASAP7_75t_L g1617 ( 
.A1(n_1598),
.A2(n_1575),
.B1(n_1573),
.B2(n_1589),
.C(n_1594),
.Y(n_1617)
);

AOI31xp33_ASAP7_75t_L g1618 ( 
.A1(n_1614),
.A2(n_1263),
.A3(n_1264),
.B(n_1554),
.Y(n_1618)
);

OAI21xp33_ASAP7_75t_SL g1619 ( 
.A1(n_1611),
.A2(n_1586),
.B(n_1536),
.Y(n_1619)
);

OAI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1596),
.A2(n_1547),
.B1(n_1536),
.B2(n_1546),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1610),
.Y(n_1621)
);

AOI222xp33_ASAP7_75t_L g1622 ( 
.A1(n_1608),
.A2(n_1569),
.B1(n_1566),
.B2(n_1563),
.C1(n_1583),
.C2(n_1551),
.Y(n_1622)
);

OAI21xp5_ASAP7_75t_SL g1623 ( 
.A1(n_1608),
.A2(n_1554),
.B(n_1558),
.Y(n_1623)
);

AOI221xp5_ASAP7_75t_L g1624 ( 
.A1(n_1601),
.A2(n_1564),
.B1(n_1558),
.B2(n_1546),
.C(n_1566),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1607),
.A2(n_1583),
.B1(n_1569),
.B2(n_1563),
.Y(n_1625)
);

OAI211xp5_ASAP7_75t_SL g1626 ( 
.A1(n_1599),
.A2(n_1564),
.B(n_1547),
.C(n_1505),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1620),
.B(n_1597),
.Y(n_1627)
);

NAND4xp75_ASAP7_75t_L g1628 ( 
.A(n_1619),
.B(n_1600),
.C(n_1613),
.D(n_1603),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1623),
.B(n_1597),
.Y(n_1629)
);

NAND4xp25_ASAP7_75t_L g1630 ( 
.A(n_1617),
.B(n_1607),
.C(n_1603),
.D(n_1606),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1622),
.B(n_1613),
.Y(n_1631)
);

NOR2x1p5_ASAP7_75t_L g1632 ( 
.A(n_1616),
.B(n_1607),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1624),
.B(n_1606),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1621),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1625),
.B(n_1604),
.Y(n_1635)
);

OAI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1615),
.A2(n_1609),
.B1(n_1601),
.B2(n_1612),
.C(n_1534),
.Y(n_1636)
);

NOR2x1_ASAP7_75t_L g1637 ( 
.A(n_1628),
.B(n_1609),
.Y(n_1637)
);

NAND4xp25_ASAP7_75t_L g1638 ( 
.A(n_1630),
.B(n_1626),
.C(n_1618),
.D(n_1462),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1632),
.B(n_1493),
.Y(n_1639)
);

AND4x1_ASAP7_75t_L g1640 ( 
.A(n_1629),
.B(n_1272),
.C(n_1501),
.D(n_1221),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1627),
.B(n_1504),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1637),
.Y(n_1642)
);

NOR3xp33_ASAP7_75t_L g1643 ( 
.A(n_1638),
.B(n_1631),
.C(n_1636),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1639),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1641),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1640),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1637),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1642),
.Y(n_1648)
);

OAI211xp5_ASAP7_75t_L g1649 ( 
.A1(n_1647),
.A2(n_1635),
.B(n_1633),
.C(n_1634),
.Y(n_1649)
);

OAI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1643),
.A2(n_1462),
.B(n_1481),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1645),
.Y(n_1651)
);

INVxp67_ASAP7_75t_SL g1652 ( 
.A(n_1643),
.Y(n_1652)
);

INVx2_ASAP7_75t_SL g1653 ( 
.A(n_1648),
.Y(n_1653)
);

NAND2x1_ASAP7_75t_L g1654 ( 
.A(n_1651),
.B(n_1646),
.Y(n_1654)
);

OAI211xp5_ASAP7_75t_SL g1655 ( 
.A1(n_1649),
.A2(n_1644),
.B(n_1392),
.C(n_1397),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1654),
.Y(n_1656)
);

NOR5xp2_ASAP7_75t_L g1657 ( 
.A(n_1656),
.B(n_1652),
.C(n_1655),
.D(n_1650),
.E(n_1653),
.Y(n_1657)
);

AOI21xp5_ASAP7_75t_L g1658 ( 
.A1(n_1657),
.A2(n_1501),
.B(n_1215),
.Y(n_1658)
);

OAI21xp5_ASAP7_75t_SL g1659 ( 
.A1(n_1657),
.A2(n_1221),
.B(n_1269),
.Y(n_1659)
);

AO21x2_ASAP7_75t_L g1660 ( 
.A1(n_1658),
.A2(n_1468),
.B(n_1467),
.Y(n_1660)
);

AO21x2_ASAP7_75t_L g1661 ( 
.A1(n_1659),
.A2(n_1468),
.B(n_1467),
.Y(n_1661)
);

OAI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1660),
.A2(n_1215),
.B(n_1216),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1660),
.B(n_1661),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1663),
.B(n_1221),
.Y(n_1664)
);

NAND3xp33_ASAP7_75t_L g1665 ( 
.A(n_1664),
.B(n_1662),
.C(n_1243),
.Y(n_1665)
);

AOI221xp5_ASAP7_75t_L g1666 ( 
.A1(n_1665),
.A2(n_1269),
.B1(n_1216),
.B2(n_1243),
.C(n_1442),
.Y(n_1666)
);

AOI211xp5_ASAP7_75t_L g1667 ( 
.A1(n_1666),
.A2(n_1269),
.B(n_1399),
.C(n_1426),
.Y(n_1667)
);


endmodule