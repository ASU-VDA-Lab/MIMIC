module fake_jpeg_16550_n_99 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_99);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_99;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

INVx8_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_25),
.B(n_7),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_48),
.B(n_49),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_0),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_1),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_51),
.B(n_37),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_51),
.A2(n_42),
.B1(n_41),
.B2(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_61),
.Y(n_66)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_50),
.A2(n_42),
.B1(n_41),
.B2(n_37),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_60),
.A2(n_44),
.B1(n_36),
.B2(n_6),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_8),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_SL g64 ( 
.A(n_62),
.B(n_43),
.C(n_36),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_64),
.A2(n_69),
.B(n_72),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_1),
.C(n_3),
.Y(n_67)
);

NOR4xp25_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_73),
.C(n_75),
.D(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_71),
.Y(n_81)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_3),
.B(n_4),
.C(n_6),
.Y(n_72)
);

BUFx2_ASAP7_75t_SL g73 ( 
.A(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_74),
.B(n_9),
.Y(n_79)
);

AND2x4_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_44),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_36),
.B(n_55),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_76),
.A2(n_77),
.B(n_82),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_55),
.B1(n_20),
.B2(n_23),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_75),
.B(n_11),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_80),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_18),
.B1(n_32),
.B2(n_31),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_67),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_86),
.B(n_87),
.Y(n_92)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_82),
.C(n_84),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_89),
.Y(n_90)
);

OAI32xp33_ASAP7_75t_L g93 ( 
.A1(n_90),
.A2(n_91),
.A3(n_85),
.B1(n_88),
.B2(n_80),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_92),
.B1(n_78),
.B2(n_13),
.Y(n_94)
);

AOI31xp33_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_83),
.A3(n_24),
.B(n_14),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_95),
.A2(n_19),
.B1(n_29),
.B2(n_15),
.Y(n_96)
);

AOI21x1_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_26),
.B(n_28),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_97),
.A2(n_16),
.B(n_17),
.Y(n_98)
);

AOI221xp5_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_27),
.B1(n_33),
.B2(n_10),
.C(n_12),
.Y(n_99)
);


endmodule