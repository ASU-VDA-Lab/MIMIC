module real_jpeg_12880_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_274, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_274;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_255;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_89;

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_3),
.A2(n_29),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_3),
.A2(n_37),
.B1(n_44),
.B2(n_45),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_4),
.A2(n_66),
.B1(n_67),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_4),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_4),
.A2(n_44),
.B1(n_45),
.B2(n_70),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_4),
.A2(n_61),
.B1(n_64),
.B2(n_70),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_4),
.A2(n_29),
.B1(n_36),
.B2(n_70),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_5),
.A2(n_66),
.B1(n_67),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_5),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_5),
.A2(n_61),
.B1(n_64),
.B2(n_72),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_72),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_5),
.A2(n_29),
.B1(n_36),
.B2(n_72),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_7),
.A2(n_61),
.B1(n_64),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_7),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_7),
.A2(n_66),
.B1(n_67),
.B2(n_137),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_7),
.A2(n_44),
.B1(n_45),
.B2(n_137),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_7),
.A2(n_29),
.B1(n_36),
.B2(n_137),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_8),
.A2(n_61),
.B1(n_64),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_8),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_81),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_8),
.A2(n_66),
.B1(n_67),
.B2(n_81),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_8),
.A2(n_29),
.B1(n_36),
.B2(n_81),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_9),
.A2(n_66),
.B1(n_67),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_9),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_9),
.A2(n_61),
.B1(n_64),
.B2(n_104),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_9),
.A2(n_44),
.B1(n_45),
.B2(n_104),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_9),
.A2(n_29),
.B1(n_36),
.B2(n_104),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_11),
.A2(n_44),
.B1(n_45),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_11),
.A2(n_29),
.B1(n_36),
.B2(n_54),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_11),
.A2(n_54),
.B1(n_61),
.B2(n_64),
.Y(n_110)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_12),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_13),
.B(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_13),
.Y(n_155)
);

AOI21xp33_ASAP7_75t_L g163 ( 
.A1(n_13),
.A2(n_66),
.B(n_164),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_L g189 ( 
.A1(n_13),
.A2(n_44),
.B1(n_45),
.B2(n_155),
.Y(n_189)
);

O2A1O1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_13),
.A2(n_44),
.B(n_50),
.C(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_13),
.B(n_111),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_13),
.B(n_33),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_13),
.B(n_55),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_13),
.A2(n_64),
.B(n_75),
.C(n_226),
.Y(n_225)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_15),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_15),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_15),
.A2(n_47),
.B1(n_61),
.B2(n_64),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_15),
.A2(n_29),
.B1(n_36),
.B2(n_47),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_16),
.A2(n_29),
.B1(n_36),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_16),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_113)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

XNOR2x2_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_127),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_126),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_105),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_22),
.B(n_105),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_83),
.C(n_89),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_23),
.B(n_83),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_56),
.B2(n_57),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_24),
.B(n_58),
.C(n_73),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_40),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_26),
.A2(n_27),
.B1(n_40),
.B2(n_41),
.Y(n_259)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_28),
.A2(n_33),
.B(n_38),
.Y(n_85)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_28),
.A2(n_33),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_28),
.A2(n_33),
.B1(n_144),
.B2(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_28),
.A2(n_33),
.B1(n_95),
.B2(n_145),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_28),
.A2(n_33),
.B1(n_158),
.B2(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_28),
.A2(n_33),
.B1(n_155),
.B2(n_211),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_28),
.A2(n_33),
.B1(n_204),
.B2(n_211),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_29),
.A2(n_36),
.B1(n_50),
.B2(n_51),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_29),
.B(n_213),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_32),
.A2(n_35),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_32),
.A2(n_93),
.B1(n_203),
.B2(n_205),
.Y(n_202)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_36),
.A2(n_51),
.B(n_155),
.Y(n_192)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_48),
.B1(n_53),
.B2(n_55),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_43),
.A2(n_52),
.B1(n_97),
.B2(n_99),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_45),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_44),
.A2(n_45),
.B1(n_77),
.B2(n_78),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_44),
.B(n_78),
.Y(n_156)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI32xp33_ASAP7_75t_L g153 ( 
.A1(n_45),
.A2(n_64),
.A3(n_77),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_48),
.A2(n_53),
.B1(n_55),
.B2(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_48),
.A2(n_55),
.B1(n_87),
.B2(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_48),
.A2(n_55),
.B1(n_147),
.B2(n_149),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_48),
.A2(n_55),
.B1(n_98),
.B2(n_149),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_48),
.A2(n_55),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_48),
.A2(n_55),
.B1(n_190),
.B2(n_197),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_52),
.A2(n_99),
.B1(n_148),
.B2(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_73),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_69),
.B2(n_71),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_59),
.A2(n_60),
.B1(n_69),
.B2(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_59),
.A2(n_60),
.B1(n_71),
.B2(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_59),
.A2(n_60),
.B1(n_163),
.B2(n_166),
.Y(n_162)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_59),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_65),
.Y(n_59)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_60),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_60)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_64),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_61),
.B(n_155),
.Y(n_154)
);

OAI32xp33_ASAP7_75t_L g178 ( 
.A1(n_61),
.A2(n_63),
.A3(n_66),
.B1(n_165),
.B2(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_63),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_62),
.B(n_64),
.Y(n_179)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_67),
.B(n_155),
.Y(n_165)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_79),
.B1(n_80),
.B2(n_82),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_74),
.A2(n_79),
.B1(n_80),
.B2(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_74),
.A2(n_79),
.B1(n_139),
.B2(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_75),
.A2(n_111),
.B1(n_135),
.B2(n_138),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_75),
.A2(n_111),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_79),
.A2(n_136),
.B(n_225),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_86),
.B2(n_88),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_88),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_84),
.A2(n_85),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_89),
.B(n_271),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_100),
.C(n_102),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_90),
.A2(n_91),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_96),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_92),
.B(n_96),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_100),
.B(n_102),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_101),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_103),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_125),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_115),
.B1(n_116),
.B2(n_124),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_112),
.B(n_114),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_112),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_123),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_117),
.Y(n_123)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_268),
.B(n_272),
.Y(n_127)
);

OAI221xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_255),
.B1(n_266),
.B2(n_267),
.C(n_274),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_239),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_182),
.B(n_238),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_159),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_132),
.B(n_159),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_146),
.C(n_150),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_133),
.B(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_140),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_134),
.B(n_141),
.C(n_143),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_143),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_142),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_146),
.A2(n_150),
.B1(n_151),
.B2(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_146),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_157),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_152),
.A2(n_153),
.B1(n_157),
.B2(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_154),
.Y(n_226)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_157),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_173),
.B2(n_181),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_160),
.B(n_174),
.C(n_180),
.Y(n_240)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_167),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_162),
.B(n_168),
.C(n_172),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_166),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_167)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_168),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_169),
.Y(n_248)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_170),
.Y(n_172)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_180),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_175),
.B(n_178),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_232),
.B(n_237),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_220),
.B(n_231),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_200),
.B(n_219),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_193),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_186),
.B(n_193),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_191),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_187),
.A2(n_188),
.B1(n_191),
.B2(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_198),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_196),
.C(n_198),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_197),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_199),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_208),
.B(n_218),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_206),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_202),
.B(n_206),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_214),
.B(n_217),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_215),
.B(n_216),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_221),
.B(n_222),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_229),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_227),
.C(n_229),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_233),
.B(n_234),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_241),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_244),
.C(n_245),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_254),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_250),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_250),
.C(n_254),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_257),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_265),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_263),
.B2(n_264),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_259),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_264),
.C(n_265),
.Y(n_269)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_260),
.Y(n_264)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_270),
.Y(n_272)
);


endmodule