module real_aes_2742_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g564 ( .A(n_0), .B(n_184), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_1), .B(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g145 ( .A(n_2), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_3), .B(n_487), .Y(n_519) );
NAND2xp33_ASAP7_75t_SL g513 ( .A(n_4), .B(n_166), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_5), .B(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g506 ( .A(n_6), .Y(n_506) );
INVx1_ASAP7_75t_L g243 ( .A(n_7), .Y(n_243) );
CKINVDCx16_ASAP7_75t_R g806 ( .A(n_8), .Y(n_806) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_9), .Y(n_235) );
AND2x2_ASAP7_75t_L g517 ( .A(n_10), .B(n_135), .Y(n_517) );
INVx2_ASAP7_75t_L g136 ( .A(n_11), .Y(n_136) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_12), .Y(n_115) );
INVx1_ASAP7_75t_L g185 ( .A(n_13), .Y(n_185) );
AOI221x1_ASAP7_75t_L g509 ( .A1(n_14), .A2(n_168), .B1(n_486), .B2(n_510), .C(n_512), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_15), .B(n_487), .Y(n_495) );
INVx1_ASAP7_75t_L g119 ( .A(n_16), .Y(n_119) );
INVx1_ASAP7_75t_L g182 ( .A(n_17), .Y(n_182) );
INVx1_ASAP7_75t_SL g157 ( .A(n_18), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_19), .B(n_160), .Y(n_199) );
AOI33xp33_ASAP7_75t_L g252 ( .A1(n_20), .A2(n_51), .A3(n_142), .B1(n_153), .B2(n_253), .B3(n_254), .Y(n_252) );
AOI221xp5_ASAP7_75t_SL g485 ( .A1(n_21), .A2(n_40), .B1(n_486), .B2(n_487), .C(n_488), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_22), .A2(n_486), .B(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_23), .B(n_184), .Y(n_522) );
INVx1_ASAP7_75t_L g776 ( .A(n_24), .Y(n_776) );
INVx1_ASAP7_75t_L g228 ( .A(n_25), .Y(n_228) );
OR2x2_ASAP7_75t_L g137 ( .A(n_26), .B(n_92), .Y(n_137) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_26), .A2(n_92), .B(n_136), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_27), .B(n_187), .Y(n_499) );
INVxp67_ASAP7_75t_L g508 ( .A(n_28), .Y(n_508) );
AND2x2_ASAP7_75t_L g553 ( .A(n_29), .B(n_134), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_30), .B(n_140), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_31), .A2(n_486), .B(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_32), .B(n_187), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g765 ( .A1(n_33), .A2(n_43), .B1(n_766), .B2(n_767), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_33), .Y(n_766) );
AND2x2_ASAP7_75t_L g147 ( .A(n_34), .B(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g152 ( .A(n_34), .Y(n_152) );
AND2x2_ASAP7_75t_L g166 ( .A(n_34), .B(n_145), .Y(n_166) );
OR2x6_ASAP7_75t_L g117 ( .A(n_35), .B(n_118), .Y(n_117) );
NOR3xp33_ASAP7_75t_L g804 ( .A(n_35), .B(n_115), .C(n_805), .Y(n_804) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_36), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_37), .B(n_140), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_38), .A2(n_169), .B1(n_175), .B2(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_39), .B(n_201), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_41), .A2(n_81), .B1(n_150), .B2(n_486), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_42), .B(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g767 ( .A(n_43), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_44), .B(n_184), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g785 ( .A1(n_45), .A2(n_786), .B1(n_787), .B2(n_790), .Y(n_785) );
INVx1_ASAP7_75t_L g790 ( .A(n_45), .Y(n_790) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_46), .B(n_203), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_47), .B(n_160), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_48), .Y(n_196) );
AND2x2_ASAP7_75t_L g567 ( .A(n_49), .B(n_134), .Y(n_567) );
OAI22xp5_ASAP7_75t_SL g787 ( .A1(n_49), .A2(n_77), .B1(n_788), .B2(n_789), .Y(n_787) );
INVxp67_ASAP7_75t_L g788 ( .A(n_49), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_50), .B(n_134), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_52), .B(n_160), .Y(n_274) );
INVx1_ASAP7_75t_L g143 ( .A(n_53), .Y(n_143) );
INVx1_ASAP7_75t_L g162 ( .A(n_53), .Y(n_162) );
AND2x2_ASAP7_75t_L g275 ( .A(n_54), .B(n_134), .Y(n_275) );
AOI221xp5_ASAP7_75t_L g241 ( .A1(n_55), .A2(n_73), .B1(n_140), .B2(n_150), .C(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_56), .B(n_140), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_57), .B(n_487), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_58), .B(n_169), .Y(n_237) );
AOI21xp5_ASAP7_75t_SL g208 ( .A1(n_59), .A2(n_150), .B(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g532 ( .A(n_60), .B(n_134), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_61), .B(n_187), .Y(n_565) );
INVx1_ASAP7_75t_L g178 ( .A(n_62), .Y(n_178) );
AND2x2_ASAP7_75t_SL g500 ( .A(n_63), .B(n_135), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_64), .B(n_184), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_65), .A2(n_486), .B(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g273 ( .A(n_66), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_67), .B(n_187), .Y(n_523) );
AND2x2_ASAP7_75t_SL g538 ( .A(n_68), .B(n_203), .Y(n_538) );
OAI22xp5_ASAP7_75t_SL g796 ( .A1(n_69), .A2(n_91), .B1(n_797), .B2(n_798), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_69), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_70), .A2(n_150), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g148 ( .A(n_71), .Y(n_148) );
INVx1_ASAP7_75t_L g164 ( .A(n_71), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_72), .B(n_140), .Y(n_255) );
AND2x2_ASAP7_75t_L g167 ( .A(n_74), .B(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g179 ( .A(n_75), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_76), .A2(n_150), .B(n_156), .Y(n_149) );
INVx1_ASAP7_75t_L g789 ( .A(n_77), .Y(n_789) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_78), .A2(n_150), .B(n_198), .C(n_202), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_79), .B(n_487), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_80), .A2(n_84), .B1(n_140), .B2(n_487), .Y(n_536) );
INVx1_ASAP7_75t_L g120 ( .A(n_82), .Y(n_120) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_82), .B(n_119), .Y(n_803) );
AND2x2_ASAP7_75t_SL g206 ( .A(n_83), .B(n_168), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g249 ( .A1(n_85), .A2(n_150), .B1(n_250), .B2(n_251), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_86), .B(n_184), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_87), .B(n_184), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_88), .B(n_112), .Y(n_111) );
XNOR2x2_ASAP7_75t_SL g763 ( .A(n_89), .B(n_764), .Y(n_763) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_90), .A2(n_486), .B(n_528), .Y(n_527) );
NOR2xp33_ASAP7_75t_SL g416 ( .A(n_91), .B(n_417), .Y(n_416) );
OAI21xp5_ASAP7_75t_L g469 ( .A1(n_91), .A2(n_470), .B(n_471), .Y(n_469) );
OAI21xp5_ASAP7_75t_L g472 ( .A1(n_91), .A2(n_417), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g798 ( .A(n_91), .Y(n_798) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_93), .Y(n_808) );
INVx1_ASAP7_75t_L g210 ( .A(n_94), .Y(n_210) );
XNOR2xp5_ASAP7_75t_L g764 ( .A(n_95), .B(n_765), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_96), .B(n_187), .Y(n_529) );
AND2x2_ASAP7_75t_L g256 ( .A(n_97), .B(n_168), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_98), .A2(n_226), .B(n_227), .C(n_229), .Y(n_225) );
INVxp67_ASAP7_75t_L g511 ( .A(n_99), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_100), .B(n_487), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_101), .B(n_187), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_102), .A2(n_486), .B(n_497), .Y(n_496) );
BUFx2_ASAP7_75t_L g110 ( .A(n_103), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_104), .B(n_160), .Y(n_211) );
AOI21xp33_ASAP7_75t_SL g105 ( .A1(n_106), .A2(n_800), .B(n_807), .Y(n_105) );
OA22x2_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_110), .B1(n_121), .B2(n_780), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
OAI21xp5_ASAP7_75t_L g780 ( .A1(n_111), .A2(n_781), .B(n_783), .Y(n_780) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_R g782 ( .A(n_114), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
AND2x6_ASAP7_75t_SL g477 ( .A(n_115), .B(n_117), .Y(n_477) );
OR2x6_ASAP7_75t_SL g762 ( .A(n_115), .B(n_116), .Y(n_762) );
OR2x2_ASAP7_75t_L g779 ( .A(n_115), .B(n_117), .Y(n_779) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
OAI21xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_763), .B(n_768), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_124), .A2(n_474), .B1(n_478), .B2(n_760), .Y(n_123) );
INVx1_ASAP7_75t_L g770 ( .A(n_124), .Y(n_770) );
NAND3xp33_ASAP7_75t_L g124 ( .A(n_125), .B(n_469), .C(n_472), .Y(n_124) );
NAND4xp25_ASAP7_75t_L g125 ( .A(n_126), .B(n_356), .C(n_416), .D(n_444), .Y(n_125) );
INVx1_ASAP7_75t_L g473 ( .A(n_126), .Y(n_473) );
NAND3x1_ASAP7_75t_L g792 ( .A(n_126), .B(n_356), .C(n_793), .Y(n_792) );
AND3x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_295), .C(n_323), .Y(n_126) );
AOI221x1_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_218), .B1(n_257), .B2(n_261), .C(n_281), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_189), .B(n_213), .Y(n_129) );
AND2x4_ASAP7_75t_L g365 ( .A(n_130), .B(n_215), .Y(n_365) );
AND2x4_ASAP7_75t_SL g130 ( .A(n_131), .B(n_171), .Y(n_130) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_131), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_131), .B(n_347), .Y(n_464) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g214 ( .A(n_132), .B(n_173), .Y(n_214) );
INVx2_ASAP7_75t_L g288 ( .A(n_132), .Y(n_288) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_132), .Y(n_348) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_132), .Y(n_355) );
AND2x2_ASAP7_75t_L g360 ( .A(n_132), .B(n_172), .Y(n_360) );
INVx1_ASAP7_75t_L g390 ( .A(n_132), .Y(n_390) );
OR2x2_ASAP7_75t_L g443 ( .A(n_132), .B(n_205), .Y(n_443) );
AO21x2_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_138), .B(n_167), .Y(n_132) );
AO21x2_ASAP7_75t_L g525 ( .A1(n_133), .A2(n_526), .B(n_532), .Y(n_525) );
AO21x2_ASAP7_75t_L g546 ( .A1(n_133), .A2(n_547), .B(n_553), .Y(n_546) );
AO21x2_ASAP7_75t_L g610 ( .A1(n_133), .A2(n_547), .B(n_553), .Y(n_610) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_134), .Y(n_133) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_134), .A2(n_485), .B(n_491), .Y(n_484) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_SL g135 ( .A(n_136), .B(n_137), .Y(n_135) );
AND2x4_ASAP7_75t_L g175 ( .A(n_136), .B(n_137), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_149), .Y(n_138) );
INVx1_ASAP7_75t_L g238 ( .A(n_140), .Y(n_238) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_140), .A2(n_150), .B1(n_505), .B2(n_507), .Y(n_504) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_146), .Y(n_140) );
INVx1_ASAP7_75t_L g194 ( .A(n_141), .Y(n_194) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
OR2x6_ASAP7_75t_L g158 ( .A(n_142), .B(n_154), .Y(n_158) );
INVxp33_ASAP7_75t_L g253 ( .A(n_142), .Y(n_253) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g155 ( .A(n_143), .B(n_145), .Y(n_155) );
AND2x4_ASAP7_75t_L g187 ( .A(n_143), .B(n_163), .Y(n_187) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g195 ( .A(n_146), .Y(n_195) );
BUFx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AND2x6_ASAP7_75t_L g486 ( .A(n_147), .B(n_155), .Y(n_486) );
INVx2_ASAP7_75t_L g154 ( .A(n_148), .Y(n_154) );
AND2x6_ASAP7_75t_L g184 ( .A(n_148), .B(n_161), .Y(n_184) );
INVxp67_ASAP7_75t_L g236 ( .A(n_150), .Y(n_236) );
AND2x4_ASAP7_75t_L g150 ( .A(n_151), .B(n_155), .Y(n_150) );
NOR2x1p5_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
INVx1_ASAP7_75t_L g254 ( .A(n_153), .Y(n_254) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
O2A1O1Ixp33_ASAP7_75t_SL g156 ( .A1(n_157), .A2(n_158), .B(n_159), .C(n_165), .Y(n_156) );
OAI22xp5_ASAP7_75t_L g177 ( .A1(n_158), .A2(n_178), .B1(n_179), .B2(n_180), .Y(n_177) );
INVx2_ASAP7_75t_L g201 ( .A(n_158), .Y(n_201) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_158), .A2(n_165), .B(n_210), .C(n_211), .Y(n_209) );
INVxp67_ASAP7_75t_L g226 ( .A(n_158), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_SL g242 ( .A1(n_158), .A2(n_165), .B(n_243), .C(n_244), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g272 ( .A1(n_158), .A2(n_165), .B(n_273), .C(n_274), .Y(n_272) );
INVx1_ASAP7_75t_L g180 ( .A(n_160), .Y(n_180) );
AND2x4_ASAP7_75t_L g487 ( .A(n_160), .B(n_166), .Y(n_487) );
AND2x4_ASAP7_75t_L g160 ( .A(n_161), .B(n_163), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_165), .B(n_175), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_165), .A2(n_199), .B(n_200), .Y(n_198) );
INVx1_ASAP7_75t_L g250 ( .A(n_165), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_165), .A2(n_489), .B(n_490), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_165), .A2(n_498), .B(n_499), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_165), .A2(n_522), .B(n_523), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_165), .A2(n_529), .B(n_530), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_165), .A2(n_550), .B(n_551), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_165), .A2(n_564), .B(n_565), .Y(n_563) );
INVx5_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
HB1xp67_ASAP7_75t_L g229 ( .A(n_166), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g224 ( .A1(n_168), .A2(n_225), .B1(n_230), .B2(n_231), .Y(n_224) );
INVx3_ASAP7_75t_L g231 ( .A(n_168), .Y(n_231) );
INVx4_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_169), .B(n_234), .Y(n_233) );
AOI21x1_ASAP7_75t_L g560 ( .A1(n_169), .A2(n_561), .B(n_567), .Y(n_560) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
BUFx4f_ASAP7_75t_L g203 ( .A(n_170), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g370 ( .A(n_171), .B(n_205), .Y(n_370) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AND2x4_ASAP7_75t_L g260 ( .A(n_172), .B(n_191), .Y(n_260) );
AND2x2_ASAP7_75t_L g347 ( .A(n_172), .B(n_217), .Y(n_347) );
INVx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g318 ( .A(n_173), .Y(n_318) );
NOR2x1_ASAP7_75t_SL g379 ( .A(n_173), .B(n_205), .Y(n_379) );
AND2x2_ASAP7_75t_L g400 ( .A(n_173), .B(n_191), .Y(n_400) );
AND2x4_ASAP7_75t_L g173 ( .A(n_174), .B(n_176), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_175), .A2(n_208), .B(n_212), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_175), .B(n_506), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_175), .B(n_508), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_175), .B(n_511), .Y(n_510) );
NOR3xp33_ASAP7_75t_L g512 ( .A(n_175), .B(n_180), .C(n_513), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_175), .A2(n_519), .B(n_520), .Y(n_518) );
OAI21xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_181), .B(n_188), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_180), .B(n_228), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B1(n_185), .B2(n_186), .Y(n_181) );
INVxp67_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVxp67_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g396 ( .A(n_189), .B(n_286), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_189), .B(n_425), .Y(n_424) );
AND2x4_ASAP7_75t_SL g189 ( .A(n_190), .B(n_204), .Y(n_189) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g217 ( .A(n_191), .Y(n_217) );
INVx1_ASAP7_75t_L g285 ( .A(n_191), .Y(n_285) );
AND2x2_ASAP7_75t_L g343 ( .A(n_191), .B(n_205), .Y(n_343) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_197), .Y(n_191) );
NOR3xp33_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .C(n_196), .Y(n_193) );
AO21x2_ASAP7_75t_L g247 ( .A1(n_202), .A2(n_248), .B(n_256), .Y(n_247) );
AO21x2_ASAP7_75t_L g294 ( .A1(n_202), .A2(n_248), .B(n_256), .Y(n_294) );
AOI21x1_ASAP7_75t_L g534 ( .A1(n_202), .A2(n_535), .B(n_538), .Y(n_534) );
INVx2_ASAP7_75t_SL g202 ( .A(n_203), .Y(n_202) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_203), .A2(n_241), .B(n_245), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_203), .A2(n_495), .B(n_496), .Y(n_494) );
NOR2x1_ASAP7_75t_L g258 ( .A(n_204), .B(n_259), .Y(n_258) );
AND2x4_ASAP7_75t_L g284 ( .A(n_204), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g322 ( .A(n_204), .B(n_214), .Y(n_322) );
INVx4_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g303 ( .A(n_205), .Y(n_303) );
AND2x4_ASAP7_75t_L g332 ( .A(n_205), .B(n_285), .Y(n_332) );
BUFx6f_ASAP7_75t_L g368 ( .A(n_205), .Y(n_368) );
AND2x2_ASAP7_75t_L g467 ( .A(n_205), .B(n_318), .Y(n_467) );
OR2x6_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
OAI21xp33_ASAP7_75t_SL g465 ( .A1(n_213), .A2(n_466), .B(n_468), .Y(n_465) );
AND2x2_ASAP7_75t_SL g213 ( .A(n_214), .B(n_215), .Y(n_213) );
NOR2xp33_ASAP7_75t_SL g340 ( .A(n_214), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_SL g422 ( .A(n_215), .Y(n_422) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx3_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_220), .A2(n_290), .B1(n_331), .B2(n_347), .Y(n_386) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_239), .Y(n_220) );
INVx1_ASAP7_75t_L g441 ( .A(n_221), .Y(n_441) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g383 ( .A(n_222), .B(n_376), .Y(n_383) );
AND2x2_ASAP7_75t_L g421 ( .A(n_222), .B(n_239), .Y(n_421) );
INVx1_ASAP7_75t_L g435 ( .A(n_222), .Y(n_435) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g265 ( .A(n_223), .Y(n_265) );
AND2x4_ASAP7_75t_L g299 ( .A(n_223), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g308 ( .A(n_223), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_223), .B(n_268), .Y(n_338) );
OR2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_232), .Y(n_223) );
AO21x2_ASAP7_75t_L g268 ( .A1(n_231), .A2(n_269), .B(n_275), .Y(n_268) );
AO21x2_ASAP7_75t_L g314 ( .A1(n_231), .A2(n_269), .B(n_275), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_236), .B1(n_237), .B2(n_238), .Y(n_232) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g279 ( .A(n_239), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g319 ( .A(n_239), .B(n_320), .Y(n_319) );
AND2x4_ASAP7_75t_L g362 ( .A(n_239), .B(n_363), .Y(n_362) );
AND2x4_ASAP7_75t_L g239 ( .A(n_240), .B(n_246), .Y(n_239) );
INVx1_ASAP7_75t_L g277 ( .A(n_240), .Y(n_277) );
INVx2_ASAP7_75t_L g300 ( .A(n_240), .Y(n_300) );
INVx1_ASAP7_75t_L g315 ( .A(n_240), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_240), .B(n_294), .Y(n_339) );
INVxp67_ASAP7_75t_L g395 ( .A(n_240), .Y(n_395) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g264 ( .A(n_247), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g298 ( .A(n_247), .Y(n_298) );
AND2x4_ASAP7_75t_L g414 ( .A(n_247), .B(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_249), .B(n_255), .Y(n_248) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
BUFx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g342 ( .A(n_259), .Y(n_342) );
OAI21xp5_ASAP7_75t_L g452 ( .A1(n_259), .A2(n_453), .B(n_454), .Y(n_452) );
INVx4_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g302 ( .A(n_260), .B(n_303), .Y(n_302) );
NAND2xp33_ASAP7_75t_SL g261 ( .A(n_262), .B(n_278), .Y(n_261) );
OR2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_266), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g468 ( .A(n_264), .B(n_313), .Y(n_468) );
AND2x2_ASAP7_75t_L g291 ( .A(n_265), .B(n_277), .Y(n_291) );
AND2x2_ASAP7_75t_L g336 ( .A(n_265), .B(n_314), .Y(n_336) );
NOR2xp67_ASAP7_75t_L g363 ( .A(n_265), .B(n_314), .Y(n_363) );
NAND2x1p5_ASAP7_75t_L g266 ( .A(n_267), .B(n_276), .Y(n_266) );
INVx3_ASAP7_75t_L g280 ( .A(n_267), .Y(n_280) );
AND2x4_ASAP7_75t_L g292 ( .A(n_267), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_267), .B(n_308), .Y(n_328) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_268), .B(n_294), .Y(n_310) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_268), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_276), .B(n_327), .Y(n_326) );
INVx3_ASAP7_75t_L g372 ( .A(n_276), .Y(n_372) );
BUFx3_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_280), .B(n_291), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_280), .B(n_348), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_282), .B(n_289), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OAI21xp5_ASAP7_75t_L g432 ( .A1(n_283), .A2(n_433), .B(n_434), .Y(n_432) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
AND2x2_ASAP7_75t_L g316 ( .A(n_284), .B(n_317), .Y(n_316) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_284), .Y(n_324) );
AND2x2_ASAP7_75t_L g438 ( .A(n_284), .B(n_439), .Y(n_438) );
NOR3xp33_ASAP7_75t_L g325 ( .A(n_286), .B(n_326), .C(n_328), .Y(n_325) );
INVx1_ASAP7_75t_L g450 ( .A(n_286), .Y(n_450) );
INVx1_ASAP7_75t_L g460 ( .A(n_286), .Y(n_460) );
AND2x2_ASAP7_75t_L g466 ( .A(n_286), .B(n_467), .Y(n_466) );
INVx3_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_287), .Y(n_439) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_290), .B(n_368), .Y(n_446) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
INVx2_ASAP7_75t_L g350 ( .A(n_291), .Y(n_350) );
INVx1_ASAP7_75t_L g349 ( .A(n_292), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_292), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g327 ( .A(n_293), .Y(n_327) );
AND2x2_ASAP7_75t_L g376 ( .A(n_293), .B(n_314), .Y(n_376) );
AND2x2_ASAP7_75t_L g394 ( .A(n_293), .B(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AOI222xp33_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_302), .B1(n_304), .B2(n_316), .C1(n_319), .C2(n_322), .Y(n_295) );
NAND2xp33_ASAP7_75t_SL g296 ( .A(n_297), .B(n_301), .Y(n_296) );
INVx2_ASAP7_75t_SL g384 ( .A(n_297), .Y(n_384) );
NAND2x1_ASAP7_75t_SL g297 ( .A(n_298), .B(n_299), .Y(n_297) );
OR2x2_ASAP7_75t_L g367 ( .A(n_298), .B(n_350), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_298), .B(n_312), .Y(n_453) );
INVx3_ASAP7_75t_L g403 ( .A(n_299), .Y(n_403) );
AND2x2_ASAP7_75t_L g413 ( .A(n_299), .B(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_302), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g392 ( .A(n_303), .Y(n_392) );
NAND2xp33_ASAP7_75t_L g304 ( .A(n_305), .B(n_311), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OAI21xp33_ASAP7_75t_SL g447 ( .A1(n_306), .A2(n_448), .B(n_451), .Y(n_447) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_307), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g312 ( .A(n_308), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NOR2x1_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx2_ASAP7_75t_L g415 ( .A(n_314), .Y(n_415) );
AND2x2_ASAP7_75t_L g331 ( .A(n_317), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NOR2x1_ASAP7_75t_L g391 ( .A(n_318), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AOI211xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_325), .B(n_329), .C(n_344), .Y(n_323) );
NAND2x1p5_ASAP7_75t_L g335 ( .A(n_327), .B(n_336), .Y(n_335) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_333), .B1(n_337), .B2(n_340), .Y(n_329) );
INVxp67_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g433 ( .A(n_332), .B(n_425), .Y(n_433) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_334), .A2(n_389), .B1(n_393), .B2(n_396), .Y(n_388) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g371 ( .A(n_335), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g393 ( .A(n_336), .B(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx2_ASAP7_75t_SL g405 ( .A(n_338), .Y(n_405) );
INVx2_ASAP7_75t_L g436 ( .A(n_339), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
AND2x2_ASAP7_75t_L g352 ( .A(n_343), .B(n_353), .Y(n_352) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_343), .A2(n_378), .B1(n_402), .B2(n_406), .Y(n_401) );
AND2x2_ASAP7_75t_L g427 ( .A(n_343), .B(n_428), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_349), .B1(n_350), .B2(n_351), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
AND2x2_ASAP7_75t_SL g385 ( .A(n_347), .B(n_368), .Y(n_385) );
INVx2_ASAP7_75t_L g411 ( .A(n_347), .Y(n_411) );
BUFx2_ASAP7_75t_L g425 ( .A(n_348), .Y(n_425) );
NOR2xp33_ASAP7_75t_SL g440 ( .A(n_349), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g378 ( .A(n_353), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVxp67_ASAP7_75t_L g470 ( .A(n_356), .Y(n_470) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_380), .Y(n_356) );
AOI21xp33_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_368), .B(n_369), .Y(n_357) );
OAI21xp33_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_361), .B(n_364), .Y(n_358) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
OAI21xp33_ASAP7_75t_L g364 ( .A1(n_360), .A2(n_365), .B(n_366), .Y(n_364) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AOI22xp33_ASAP7_75t_SL g437 ( .A1(n_362), .A2(n_438), .B1(n_440), .B2(n_442), .Y(n_437) );
AOI22xp33_ASAP7_75t_SL g382 ( .A1(n_365), .A2(n_383), .B1(n_384), .B2(n_385), .Y(n_382) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g398 ( .A(n_368), .B(n_399), .Y(n_398) );
OR2x6_ASAP7_75t_L g410 ( .A(n_368), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g412 ( .A(n_368), .B(n_400), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_371), .B1(n_373), .B2(n_377), .Y(n_369) );
NOR2xp67_ASAP7_75t_SL g374 ( .A(n_372), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g457 ( .A(n_372), .Y(n_457) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g429 ( .A(n_379), .Y(n_429) );
NOR2xp67_ASAP7_75t_L g380 ( .A(n_381), .B(n_387), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_386), .Y(n_381) );
NAND4xp25_ASAP7_75t_L g387 ( .A(n_388), .B(n_397), .C(n_401), .D(n_408), .Y(n_387) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
AND2x2_ASAP7_75t_L g399 ( .A(n_390), .B(n_400), .Y(n_399) );
NAND2x1p5_ASAP7_75t_L g430 ( .A(n_394), .B(n_405), .Y(n_430) );
NAND2xp33_ASAP7_75t_SL g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g420 ( .A(n_407), .Y(n_420) );
OAI21xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_412), .B(n_413), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g459 ( .A(n_414), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g793 ( .A(n_418), .B(n_794), .Y(n_793) );
AOI211x1_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_422), .B(n_423), .C(n_431), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_422), .B(n_450), .Y(n_451) );
AOI31xp33_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_426), .A3(n_429), .B(n_430), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_437), .Y(n_431) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_436), .B(n_462), .Y(n_461) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_439), .Y(n_455) );
INVx2_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g471 ( .A(n_444), .Y(n_471) );
AOI21xp33_ASAP7_75t_SL g444 ( .A1(n_445), .A2(n_452), .B(n_456), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g794 ( .A1(n_445), .A2(n_452), .B(n_456), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVxp33_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OAI211xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_458), .B(n_461), .C(n_465), .Y(n_456) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OAI21x1_ASAP7_75t_L g769 ( .A1(n_474), .A2(n_770), .B(n_771), .Y(n_769) );
CKINVDCx6p67_ASAP7_75t_R g474 ( .A(n_475), .Y(n_474) );
INVx3_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g476 ( .A(n_477), .Y(n_476) );
NAND2x1_ASAP7_75t_SL g771 ( .A(n_478), .B(n_772), .Y(n_771) );
INVx4_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
OR2x6_ASAP7_75t_L g479 ( .A(n_480), .B(n_673), .Y(n_479) );
NAND3xp33_ASAP7_75t_SL g480 ( .A(n_481), .B(n_583), .C(n_623), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_501), .B(n_514), .C(n_539), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_482), .B(n_588), .Y(n_622) );
NOR2x1p5_ASAP7_75t_L g482 ( .A(n_483), .B(n_492), .Y(n_482) );
BUFx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g558 ( .A(n_484), .Y(n_558) );
INVx2_ASAP7_75t_L g574 ( .A(n_484), .Y(n_574) );
OR2x2_ASAP7_75t_L g586 ( .A(n_484), .B(n_493), .Y(n_586) );
AND2x2_ASAP7_75t_L g600 ( .A(n_484), .B(n_559), .Y(n_600) );
INVx1_ASAP7_75t_L g628 ( .A(n_484), .Y(n_628) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_484), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_484), .B(n_493), .Y(n_734) );
OR2x2_ASAP7_75t_L g555 ( .A(n_492), .B(n_556), .Y(n_555) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_492), .Y(n_690) );
AND2x2_ASAP7_75t_L g695 ( .A(n_492), .B(n_557), .Y(n_695) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x4_ASAP7_75t_L g501 ( .A(n_493), .B(n_502), .Y(n_501) );
OR2x2_ASAP7_75t_L g554 ( .A(n_493), .B(n_503), .Y(n_554) );
OR2x2_ASAP7_75t_L g573 ( .A(n_493), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g602 ( .A(n_493), .Y(n_602) );
AND2x4_ASAP7_75t_SL g641 ( .A(n_493), .B(n_503), .Y(n_641) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_493), .Y(n_645) );
OR2x2_ASAP7_75t_L g662 ( .A(n_493), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g672 ( .A(n_493), .B(n_579), .Y(n_672) );
INVx1_ASAP7_75t_L g701 ( .A(n_493), .Y(n_701) );
OR2x6_ASAP7_75t_L g493 ( .A(n_494), .B(n_500), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_501), .B(n_630), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_502), .B(n_559), .Y(n_576) );
AND2x2_ASAP7_75t_L g588 ( .A(n_502), .B(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g606 ( .A(n_502), .B(n_573), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_502), .B(n_627), .Y(n_626) );
INVx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x4_ASAP7_75t_L g579 ( .A(n_503), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g601 ( .A(n_503), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g636 ( .A(n_503), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_503), .B(n_559), .Y(n_660) );
AND2x4_ASAP7_75t_L g503 ( .A(n_504), .B(n_509), .Y(n_503) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_524), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_515), .B(n_592), .Y(n_591) );
AND2x4_ASAP7_75t_L g609 ( .A(n_515), .B(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_515), .B(n_525), .Y(n_614) );
NAND3xp33_ASAP7_75t_L g629 ( .A(n_515), .B(n_630), .C(n_631), .Y(n_629) );
AND2x2_ASAP7_75t_L g677 ( .A(n_515), .B(n_582), .Y(n_677) );
INVx5_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g544 ( .A(n_516), .B(n_545), .Y(n_544) );
AND2x4_ASAP7_75t_SL g581 ( .A(n_516), .B(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g597 ( .A(n_516), .Y(n_597) );
OR2x2_ASAP7_75t_L g620 ( .A(n_516), .B(n_610), .Y(n_620) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_516), .Y(n_637) );
AND2x2_ASAP7_75t_SL g655 ( .A(n_516), .B(n_543), .Y(n_655) );
AND2x4_ASAP7_75t_L g670 ( .A(n_516), .B(n_546), .Y(n_670) );
AND2x2_ASAP7_75t_L g684 ( .A(n_516), .B(n_525), .Y(n_684) );
OR2x2_ASAP7_75t_L g705 ( .A(n_516), .B(n_533), .Y(n_705) );
OR2x6_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
AND2x2_ASAP7_75t_L g759 ( .A(n_524), .B(n_637), .Y(n_759) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_533), .Y(n_524) );
AND2x4_ASAP7_75t_L g582 ( .A(n_525), .B(n_545), .Y(n_582) );
INVx2_ASAP7_75t_L g593 ( .A(n_525), .Y(n_593) );
AND2x2_ASAP7_75t_L g598 ( .A(n_525), .B(n_543), .Y(n_598) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_525), .Y(n_631) );
OR2x2_ASAP7_75t_L g654 ( .A(n_525), .B(n_546), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_525), .B(n_546), .Y(n_657) );
INVx1_ASAP7_75t_L g666 ( .A(n_525), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_531), .Y(n_526) );
AND2x2_ASAP7_75t_L g569 ( .A(n_533), .B(n_546), .Y(n_569) );
BUFx2_ASAP7_75t_L g618 ( .A(n_533), .Y(n_618) );
AND2x2_ASAP7_75t_L g713 ( .A(n_533), .B(n_593), .Y(n_713) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_534), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
OAI221xp5_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_554), .B1(n_555), .B2(n_568), .C(n_570), .Y(n_539) );
INVx1_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_544), .Y(n_541) );
NOR2x1_ASAP7_75t_L g615 ( .A(n_542), .B(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_542), .B(n_609), .Y(n_649) );
OR2x2_ASAP7_75t_L g661 ( .A(n_542), .B(n_657), .Y(n_661) );
OR2x2_ASAP7_75t_L g664 ( .A(n_542), .B(n_665), .Y(n_664) );
OR2x2_ASAP7_75t_L g753 ( .A(n_542), .B(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x4_ASAP7_75t_L g592 ( .A(n_543), .B(n_593), .Y(n_592) );
OA33x2_ASAP7_75t_L g625 ( .A1(n_543), .A2(n_586), .A3(n_626), .B1(n_629), .B2(n_632), .B3(n_635), .Y(n_625) );
OR2x2_ASAP7_75t_L g656 ( .A(n_543), .B(n_657), .Y(n_656) );
OR2x2_ASAP7_75t_L g680 ( .A(n_543), .B(n_681), .Y(n_680) );
OR2x2_ASAP7_75t_L g688 ( .A(n_543), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g708 ( .A(n_543), .B(n_582), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_543), .B(n_597), .Y(n_746) );
INVx2_ASAP7_75t_L g616 ( .A(n_544), .Y(n_616) );
AOI322xp5_ASAP7_75t_L g686 ( .A1(n_544), .A2(n_599), .A3(n_687), .B1(n_690), .B2(n_691), .C1(n_693), .C2(n_695), .Y(n_686) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_546), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_552), .Y(n_547) );
OR2x2_ASAP7_75t_L g668 ( .A(n_554), .B(n_647), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_554), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g741 ( .A(n_554), .Y(n_741) );
INVx1_ASAP7_75t_SL g607 ( .A(n_555), .Y(n_607) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g640 ( .A(n_557), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
INVx2_ASAP7_75t_L g580 ( .A(n_559), .Y(n_580) );
INVx1_ASAP7_75t_L g589 ( .A(n_559), .Y(n_589) );
INVx1_ASAP7_75t_L g630 ( .A(n_559), .Y(n_630) );
OR2x2_ASAP7_75t_L g647 ( .A(n_559), .B(n_574), .Y(n_647) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_559), .Y(n_722) );
INVx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_566), .Y(n_561) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_SL g691 ( .A(n_569), .B(n_692), .Y(n_691) );
OAI21xp5_ASAP7_75t_SL g570 ( .A1(n_571), .A2(n_577), .B(n_581), .Y(n_570) );
A2O1A1Ixp33_ASAP7_75t_L g644 ( .A1(n_571), .A2(n_645), .B(n_646), .C(n_648), .Y(n_644) );
AND2x4_ASAP7_75t_L g571 ( .A(n_572), .B(n_575), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g709 ( .A(n_573), .B(n_710), .Y(n_709) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_574), .Y(n_578) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g733 ( .A(n_576), .B(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
AND2x2_ASAP7_75t_SL g702 ( .A(n_579), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g710 ( .A(n_579), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_579), .B(n_701), .Y(n_718) );
INVx3_ASAP7_75t_SL g643 ( .A(n_582), .Y(n_643) );
AOI221xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_590), .B1(n_594), .B2(n_599), .C(n_603), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_589), .Y(n_634) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AOI21xp5_ASAP7_75t_L g697 ( .A1(n_592), .A2(n_619), .B(n_691), .Y(n_697) );
AND2x2_ASAP7_75t_L g723 ( .A(n_592), .B(n_670), .Y(n_723) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_593), .Y(n_611) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_597), .B(n_713), .Y(n_712) );
OR2x2_ASAP7_75t_L g732 ( .A(n_597), .B(n_654), .Y(n_732) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx2_ASAP7_75t_L g681 ( .A(n_600), .Y(n_681) );
OAI21xp33_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_608), .B(n_612), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .Y(n_608) );
INVx2_ASAP7_75t_L g754 ( .A(n_609), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_610), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g683 ( .A(n_610), .B(n_684), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_611), .B(n_633), .Y(n_632) );
OAI31xp33_ASAP7_75t_SL g612 ( .A1(n_613), .A2(n_615), .A3(n_617), .B(n_621), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_616), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
OR2x2_ASAP7_75t_L g694 ( .A(n_618), .B(n_620), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_618), .B(n_670), .Y(n_749) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NOR5xp2_ASAP7_75t_L g623 ( .A(n_624), .B(n_638), .C(n_650), .D(n_659), .E(n_667), .Y(n_623) );
INVxp67_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_628), .B(n_630), .Y(n_663) );
INVx1_ASAP7_75t_L g703 ( .A(n_628), .Y(n_703) );
INVxp67_ASAP7_75t_SL g740 ( .A(n_628), .Y(n_740) );
INVx1_ASAP7_75t_L g692 ( .A(n_631), .Y(n_692) );
INVxp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp33_ASAP7_75t_SL g635 ( .A(n_636), .B(n_637), .Y(n_635) );
OAI321xp33_ASAP7_75t_L g675 ( .A1(n_636), .A2(n_676), .A3(n_678), .B1(n_682), .B2(n_685), .C(n_686), .Y(n_675) );
INVx1_ASAP7_75t_L g729 ( .A(n_637), .Y(n_729) );
OAI21xp33_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_642), .B(n_644), .Y(n_638) );
INVx1_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_640), .A2(n_713), .B1(n_720), .B2(n_723), .Y(n_719) );
AND2x2_ASAP7_75t_L g748 ( .A(n_641), .B(n_722), .Y(n_748) );
INVx1_ASAP7_75t_L g658 ( .A(n_646), .Y(n_658) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AOI21xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_656), .B(n_658), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_657), .A2(n_668), .B1(n_669), .B2(n_671), .Y(n_667) );
INVx1_ASAP7_75t_L g730 ( .A(n_657), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_661), .B1(n_662), .B2(n_664), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_666), .B(n_670), .Y(n_669) );
OAI221xp5_ASAP7_75t_L g744 ( .A1(n_668), .A2(n_745), .B1(n_747), .B2(n_749), .C(n_750), .Y(n_744) );
INVx1_ASAP7_75t_L g751 ( .A(n_668), .Y(n_751) );
OAI221xp5_ASAP7_75t_L g725 ( .A1(n_669), .A2(n_726), .B1(n_733), .B2(n_735), .C(n_736), .Y(n_725) );
OAI21xp5_ASAP7_75t_L g696 ( .A1(n_671), .A2(n_697), .B(n_698), .Y(n_696) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_724), .Y(n_673) );
NOR3xp33_ASAP7_75t_L g674 ( .A(n_675), .B(n_696), .C(n_714), .Y(n_674) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_677), .Y(n_743) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx3_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g742 ( .A(n_685), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_687), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g735 ( .A(n_695), .Y(n_735) );
AOI21xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_704), .B(n_706), .Y(n_698) );
INVxp67_ASAP7_75t_L g756 ( .A(n_699), .Y(n_756) );
AND2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_702), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_SL g711 ( .A(n_702), .Y(n_711) );
INVx1_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
OAI22xp33_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_709), .B1(n_711), .B2(n_712), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OAI21xp33_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_716), .B(n_719), .Y(n_714) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g757 ( .A(n_720), .Y(n_757) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
NOR3xp33_ASAP7_75t_L g724 ( .A(n_725), .B(n_744), .C(n_755), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_727), .B(n_731), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_SL g728 ( .A(n_729), .B(n_730), .Y(n_728) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
OAI21xp5_ASAP7_75t_SL g736 ( .A1(n_737), .A2(n_742), .B(n_743), .Y(n_736) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_739), .B(n_741), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVxp67_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
OAI21xp5_ASAP7_75t_L g750 ( .A1(n_748), .A2(n_751), .B(n_752), .Y(n_750) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
AOI21xp33_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_757), .B(n_758), .Y(n_755) );
INVx1_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_761), .Y(n_774) );
CKINVDCx11_ASAP7_75t_R g761 ( .A(n_762), .Y(n_761) );
AOI21xp33_ASAP7_75t_SL g768 ( .A1(n_763), .A2(n_769), .B(n_775), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_773), .Y(n_772) );
BUFx4f_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_776), .B(n_777), .Y(n_775) );
INVx1_ASAP7_75t_SL g777 ( .A(n_778), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_SL g781 ( .A(n_782), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_785), .B1(n_791), .B2(n_799), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g799 ( .A(n_791), .Y(n_799) );
XOR2x2_ASAP7_75t_L g791 ( .A(n_792), .B(n_795), .Y(n_791) );
CKINVDCx5p33_ASAP7_75t_R g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_SL g810 ( .A(n_801), .Y(n_810) );
INVx3_ASAP7_75t_SL g801 ( .A(n_802), .Y(n_801) );
AND2x2_ASAP7_75t_SL g802 ( .A(n_803), .B(n_804), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .Y(n_807) );
HB1xp67_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
endmodule