module real_jpeg_4083_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_0),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_0),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_0),
.B(n_187),
.Y(n_186)
);

AND2x2_ASAP7_75t_SL g214 ( 
.A(n_0),
.B(n_215),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_0),
.B(n_230),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_0),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_0),
.B(n_248),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_0),
.B(n_425),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_1),
.Y(n_522)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_2),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_2),
.Y(n_257)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_2),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_2),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_2),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_3),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_3),
.Y(n_103)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_3),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_3),
.Y(n_171)
);

INVx6_ASAP7_75t_L g453 ( 
.A(n_3),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_3),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_4),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_4),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_4),
.B(n_239),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_4),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_4),
.B(n_57),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_4),
.B(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_4),
.B(n_50),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_5),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_5),
.B(n_192),
.Y(n_191)
);

AND2x2_ASAP7_75t_SL g217 ( 
.A(n_5),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_5),
.B(n_396),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_5),
.B(n_439),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_6),
.B(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_6),
.B(n_227),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_6),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_6),
.B(n_306),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_6),
.B(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_6),
.B(n_285),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_6),
.B(n_402),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_6),
.B(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_7),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_7),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_7),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_7),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_7),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_7),
.B(n_192),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_7),
.B(n_387),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_7),
.B(n_312),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_8),
.Y(n_100)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_8),
.Y(n_118)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_8),
.Y(n_143)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_9),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_10),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_10),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_10),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_10),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_10),
.B(n_159),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g383 ( 
.A(n_10),
.B(n_384),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_10),
.B(n_448),
.Y(n_447)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_11),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g312 ( 
.A(n_11),
.Y(n_312)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_13),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_13),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_13),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_14),
.B(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_14),
.Y(n_71)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_14),
.B(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_14),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_14),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_14),
.B(n_163),
.Y(n_162)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_16),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_16),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_16),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_16),
.B(n_126),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_16),
.B(n_255),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_16),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_16),
.B(n_312),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_16),
.B(n_434),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_17),
.B(n_233),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_17),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_17),
.B(n_283),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_17),
.B(n_293),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_17),
.B(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_17),
.B(n_239),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_17),
.B(n_437),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_17),
.B(n_476),
.Y(n_475)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_19),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_19),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_19),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_19),
.B(n_303),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_19),
.B(n_312),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g342 ( 
.A(n_19),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_19),
.B(n_212),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_517),
.B(n_519),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_173),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_172),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_151),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_24),
.B(n_151),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_109),
.C(n_121),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_25),
.B(n_503),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_77),
.C(n_90),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g505 ( 
.A(n_26),
.B(n_506),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_46),
.C(n_59),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_27),
.B(n_46),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_28),
.B(n_38),
.C(n_45),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_29),
.B(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_29),
.B(n_251),
.Y(n_250)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_31),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_38),
.B1(n_39),
.B2(n_45),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g248 ( 
.A(n_35),
.Y(n_248)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_37),
.Y(n_134)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_37),
.Y(n_228)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_37),
.Y(n_441)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_43),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_43),
.Y(n_344)
);

INVx6_ASAP7_75t_L g398 ( 
.A(n_43),
.Y(n_398)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g216 ( 
.A(n_44),
.Y(n_216)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_44),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_44),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_46),
.B(n_466),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_46),
.B(n_462),
.C(n_466),
.Y(n_487)
);

FAx1_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_51),
.CI(n_54),
.CON(n_46),
.SN(n_46)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_58),
.Y(n_231)
);

INVx5_ASAP7_75t_L g286 ( 
.A(n_58),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_59),
.B(n_495),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_65),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_60),
.B(n_66),
.C(n_76),
.Y(n_119)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_62),
.Y(n_196)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_64),
.Y(n_206)
);

INVx6_ASAP7_75t_L g428 ( 
.A(n_64),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_70),
.B2(n_76),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_66),
.A2(n_67),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_66),
.B(n_112),
.C(n_116),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_93),
.C(n_97),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_70),
.A2(n_76),
.B1(n_93),
.B2(n_94),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_75),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_75),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_77),
.A2(n_90),
.B1(n_91),
.B2(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_77),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_78),
.B(n_82),
.C(n_85),
.Y(n_139)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_89),
.Y(n_163)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_101),
.C(n_104),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_92),
.B(n_493),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_93),
.A2(n_94),
.B1(n_447),
.B2(n_449),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_93),
.B(n_447),
.C(n_450),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_96),
.Y(n_194)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_96),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_97),
.B(n_464),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_100),
.Y(n_199)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_100),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_101),
.A2(n_102),
.B1(n_104),
.B2(n_105),
.Y(n_493)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_104),
.A2(n_105),
.B1(n_475),
.B2(n_477),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_105),
.B(n_477),
.C(n_491),
.Y(n_490)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_108),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_109),
.B(n_121),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_119),
.C(n_120),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_110),
.B(n_509),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_116),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_112),
.A2(n_113),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_113),
.B(n_131),
.C(n_135),
.Y(n_167)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx5_ASAP7_75t_L g316 ( 
.A(n_115),
.Y(n_316)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_119),
.B(n_120),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_138),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_136),
.B2(n_137),
.Y(n_122)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_137),
.C(n_138),
.Y(n_152)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_129),
.B1(n_130),
.B2(n_135),
.Y(n_124)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_128),
.Y(n_212)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_131),
.A2(n_132),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_144),
.C(n_150),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_144),
.B1(n_145),
.B2(n_150),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_141),
.Y(n_150)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_143),
.Y(n_437)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_165),
.B2(n_166),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_162),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

AO21x1_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_498),
.B(n_514),
.Y(n_173)
);

OAI21x1_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_482),
.B(n_497),
.Y(n_174)
);

AOI21x1_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_457),
.B(n_481),
.Y(n_175)
);

OAI21x1_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_411),
.B(n_456),
.Y(n_176)
);

AOI21x1_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_373),
.B(n_410),
.Y(n_177)
);

AO21x1_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_296),
.B(n_372),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_276),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_180),
.B(n_276),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_223),
.B2(n_275),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_181),
.B(n_224),
.C(n_258),
.Y(n_409)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_200),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_183),
.B(n_201),
.C(n_222),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_195),
.C(n_197),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_184),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_190),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_185),
.A2(n_186),
.B1(n_190),
.B2(n_191),
.Y(n_281)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_195),
.B(n_197),
.Y(n_295)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_208),
.B1(n_221),
.B2(n_222),
.Y(n_200)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_201),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B(n_207),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_203),
.Y(n_207)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_207),
.B(n_389),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_207),
.B(n_378),
.C(n_389),
.Y(n_418)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_208),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_213),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_209),
.B(n_214),
.C(n_217),
.Y(n_408)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.Y(n_213)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx8_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_223),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_258),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_235),
.C(n_249),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_225),
.B(n_278),
.Y(n_277)
);

BUFx24_ASAP7_75t_SL g524 ( 
.A(n_225),
.Y(n_524)
);

FAx1_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_229),
.CI(n_232),
.CON(n_225),
.SN(n_225)
);

MAJx2_ASAP7_75t_L g274 ( 
.A(n_226),
.B(n_229),
.C(n_232),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_228),
.Y(n_261)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_234),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_235),
.A2(n_236),
.B1(n_249),
.B2(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

MAJx2_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_241),
.C(n_246),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_237),
.A2(n_238),
.B1(n_246),
.B2(n_247),
.Y(n_365)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx8_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_241),
.B(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_249),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_254),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_254),
.Y(n_273)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

BUFx8_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_253),
.Y(n_269)
);

BUFx5_ASAP7_75t_L g293 ( 
.A(n_253),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_253),
.Y(n_387)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_257),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_272),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_259),
.B(n_273),
.C(n_274),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

MAJx2_ASAP7_75t_L g389 ( 
.A(n_260),
.B(n_267),
.C(n_270),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_267),
.B1(n_270),
.B2(n_271),
.Y(n_262)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_263),
.Y(n_270)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx8_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_267),
.Y(n_271)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_280),
.C(n_294),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_277),
.B(n_370),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_280),
.B(n_294),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.C(n_287),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_281),
.B(n_282),
.Y(n_358)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_287),
.B(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_292),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_288),
.B(n_292),
.Y(n_338)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

OAI21x1_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_367),
.B(n_371),
.Y(n_296)
);

OA21x2_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_352),
.B(n_366),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_335),
.B(n_351),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_300),
.A2(n_325),
.B(n_334),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_308),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_301),
.B(n_308),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_305),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_302),
.B(n_305),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_302),
.B(n_330),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

BUFx5_ASAP7_75t_L g448 ( 
.A(n_304),
.Y(n_448)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_310),
.B1(n_317),
.B2(n_318),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_313),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_311),
.B(n_313),
.C(n_317),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_323),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_319),
.B(n_323),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_329),
.B(n_333),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_328),
.Y(n_333)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_350),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_336),
.B(n_350),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_340),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_338),
.B(n_339),
.C(n_354),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_340),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_341),
.B(n_345),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_341),
.B(n_347),
.C(n_349),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

INVx11_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_347),
.B1(n_348),
.B2(n_349),
.Y(n_345)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_346),
.Y(n_349)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_355),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_353),
.B(n_355),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_356),
.A2(n_357),
.B1(n_359),
.B2(n_360),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_356),
.B(n_362),
.C(n_363),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_362),
.B1(n_363),
.B2(n_364),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_364),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_369),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_368),
.B(n_369),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_374),
.B(n_409),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_374),
.B(n_409),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_391),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_376),
.B(n_377),
.C(n_391),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_379),
.B1(n_388),
.B2(n_390),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_381),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_380),
.B(n_383),
.C(n_385),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_382),
.A2(n_383),
.B1(n_385),
.B2(n_386),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_388),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_392),
.B(n_393),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_392),
.B(n_394),
.C(n_404),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_404),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_399),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_395),
.B(n_400),
.C(n_401),
.Y(n_443)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_401),
.Y(n_399)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_408),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_406),
.B(n_407),
.C(n_408),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_413),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_412),
.B(n_413),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_415),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_414),
.B(n_431),
.C(n_454),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_416),
.A2(n_431),
.B1(n_454),
.B2(n_455),
.Y(n_415)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_416),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_417),
.A2(n_418),
.B1(n_419),
.B2(n_430),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_417),
.B(n_420),
.C(n_421),
.Y(n_459)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_419),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_420),
.B(n_421),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_429),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_423),
.B(n_424),
.C(n_429),
.Y(n_472)
);

INVx6_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx5_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_431),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_442),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_432),
.B(n_443),
.C(n_444),
.Y(n_470)
);

BUFx24_ASAP7_75t_SL g527 ( 
.A(n_432),
.Y(n_527)
);

FAx1_ASAP7_75t_SL g432 ( 
.A(n_433),
.B(n_436),
.CI(n_438),
.CON(n_432),
.SN(n_432)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_433),
.B(n_436),
.C(n_438),
.Y(n_478)
);

INVx5_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_444),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_445),
.A2(n_446),
.B1(n_450),
.B2(n_451),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_447),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_458),
.B(n_480),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_458),
.B(n_480),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_460),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_459),
.B(n_461),
.C(n_468),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_468),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_462),
.A2(n_463),
.B1(n_465),
.B2(n_467),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_465),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_469),
.A2(n_470),
.B1(n_471),
.B2(n_479),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_469),
.B(n_472),
.C(n_473),
.Y(n_484)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_471),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_472),
.B(n_473),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_478),
.Y(n_473)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_475),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_478),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_483),
.B(n_496),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_483),
.B(n_496),
.Y(n_497)
);

BUFx24_ASAP7_75t_SL g525 ( 
.A(n_483),
.Y(n_525)
);

FAx1_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_485),
.CI(n_494),
.CON(n_483),
.SN(n_483)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_484),
.B(n_485),
.C(n_494),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_486),
.A2(n_487),
.B1(n_488),
.B2(n_489),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_486),
.B(n_490),
.C(n_492),
.Y(n_510)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_492),
.Y(n_489)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_511),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_501),
.A2(n_515),
.B(n_516),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_502),
.B(n_504),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_502),
.B(n_504),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_508),
.C(n_510),
.Y(n_504)
);

FAx1_ASAP7_75t_SL g512 ( 
.A(n_505),
.B(n_508),
.CI(n_510),
.CON(n_512),
.SN(n_512)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_513),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_512),
.B(n_513),
.Y(n_515)
);

BUFx24_ASAP7_75t_SL g523 ( 
.A(n_512),
.Y(n_523)
);

INVx8_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx13_ASAP7_75t_L g521 ( 
.A(n_518),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_522),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);


endmodule