module fake_jpeg_8593_n_29 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_29);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_29;

wire n_13;
wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_12;
wire n_15;

INVx13_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_8),
.B(n_3),
.Y(n_13)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_10),
.A2(n_0),
.B(n_5),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g15 ( 
.A(n_4),
.B(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_17),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_19),
.Y(n_24)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_1),
.C(n_2),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_21),
.C(n_22),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_1),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_21),
.A2(n_12),
.B1(n_13),
.B2(n_16),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_26),
.B(n_27),
.Y(n_28)
);

OAI321xp33_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_25),
.A3(n_7),
.B1(n_9),
.B2(n_6),
.C(n_19),
.Y(n_29)
);


endmodule