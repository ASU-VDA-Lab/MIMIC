module fake_jpeg_8267_n_275 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_275);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_275;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_42),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_17),
.B(n_7),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_33),
.B1(n_22),
.B2(n_18),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_44),
.A2(n_31),
.B1(n_21),
.B2(n_30),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_42),
.B(n_32),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_19),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_20),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_59),
.Y(n_84)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_48),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_27),
.Y(n_48)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_27),
.Y(n_58)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_20),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_60),
.Y(n_69)
);

HAxp5_ASAP7_75t_SL g61 ( 
.A(n_40),
.B(n_17),
.CON(n_61),
.SN(n_61)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_61),
.A2(n_62),
.B1(n_32),
.B2(n_19),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_35),
.A2(n_33),
.B1(n_22),
.B2(n_18),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_20),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_64),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_32),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_51),
.A2(n_35),
.B1(n_43),
.B2(n_39),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_67),
.A2(n_70),
.B1(n_72),
.B2(n_66),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_35),
.B1(n_39),
.B2(n_22),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_39),
.B1(n_33),
.B2(n_18),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_74),
.B(n_77),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_75)
);

AO21x1_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_86),
.B(n_89),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_52),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_83),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_37),
.C(n_41),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_55),
.C(n_37),
.Y(n_98)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_65),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_52),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_51),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_55),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_54),
.A2(n_19),
.B1(n_31),
.B2(n_21),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_89),
.B1(n_56),
.B2(n_45),
.Y(n_100)
);

AO22x1_ASAP7_75t_SL g89 ( 
.A1(n_63),
.A2(n_37),
.B1(n_41),
.B2(n_34),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_91),
.A2(n_107),
.B1(n_110),
.B2(n_113),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_77),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_47),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_94),
.B(n_60),
.Y(n_131)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_87),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_106),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_99),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_101),
.C(n_102),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_89),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_100),
.A2(n_109),
.B1(n_28),
.B2(n_23),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_46),
.C(n_37),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_60),
.C(n_41),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_88),
.B1(n_85),
.B2(n_83),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_72),
.A2(n_34),
.B(n_16),
.C(n_50),
.Y(n_104)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_104),
.A2(n_75),
.B(n_77),
.C(n_57),
.D(n_50),
.Y(n_124)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_107),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_49),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_66),
.B1(n_29),
.B2(n_23),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_111),
.Y(n_121)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_113),
.Y(n_134)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_118),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_116),
.A2(n_122),
.B1(n_136),
.B2(n_100),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_68),
.B1(n_71),
.B2(n_76),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_117),
.A2(n_123),
.B1(n_26),
.B2(n_24),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_68),
.B1(n_71),
.B2(n_70),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_124),
.A2(n_126),
.B1(n_137),
.B2(n_29),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_108),
.A2(n_81),
.B1(n_75),
.B2(n_69),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_130),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_69),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_98),
.C(n_102),
.Y(n_140)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_133),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_106),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_96),
.B(n_81),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_138),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_97),
.A2(n_28),
.B1(n_30),
.B2(n_24),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_93),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_126),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_142),
.Y(n_181)
);

AND2x6_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_94),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_143),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_119),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_144),
.B(n_150),
.Y(n_168)
);

AND2x6_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_94),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_146),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_101),
.Y(n_147)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_133),
.Y(n_148)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_115),
.A2(n_105),
.B1(n_91),
.B2(n_108),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_114),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_91),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_151),
.A2(n_161),
.B(n_163),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_92),
.C(n_109),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_140),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_104),
.Y(n_153)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_155),
.A2(n_159),
.B1(n_137),
.B2(n_163),
.Y(n_180)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_156),
.B(n_157),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_138),
.B(n_25),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_116),
.A2(n_24),
.B1(n_29),
.B2(n_26),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_158),
.A2(n_128),
.B1(n_26),
.B2(n_29),
.Y(n_175)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_123),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_124),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_134),
.A2(n_60),
.B(n_50),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_129),
.B(n_24),
.Y(n_162)
);

XNOR2x1_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_129),
.Y(n_179)
);

OAI21x1_ASAP7_75t_R g163 ( 
.A1(n_121),
.A2(n_16),
.B(n_50),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_176),
.C(n_152),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_163),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_170),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_179),
.B(n_139),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_125),
.Y(n_174)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_180),
.B1(n_184),
.B2(n_186),
.Y(n_193)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_188),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_130),
.Y(n_182)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_150),
.A2(n_156),
.B1(n_155),
.B2(n_151),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_151),
.A2(n_128),
.B1(n_130),
.B2(n_118),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_145),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_168),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_194),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_192),
.C(n_199),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_147),
.C(n_143),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_178),
.B(n_148),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_181),
.A2(n_146),
.B1(n_162),
.B2(n_164),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_195),
.A2(n_177),
.B1(n_166),
.B2(n_10),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_173),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_203),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_139),
.C(n_153),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_160),
.C(n_161),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_202),
.C(n_208),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_164),
.C(n_49),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_26),
.Y(n_206)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_180),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_49),
.C(n_1),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_0),
.C(n_1),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_187),
.C(n_171),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_186),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_221),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_198),
.A2(n_177),
.B1(n_183),
.B2(n_171),
.Y(n_214)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_215),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_205),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_217),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_166),
.C(n_179),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_224),
.C(n_200),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_187),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_208),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_6),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_206),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_226),
.A2(n_220),
.B1(n_197),
.B2(n_222),
.Y(n_227)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_223),
.A2(n_204),
.B1(n_191),
.B2(n_193),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_235),
.C(n_212),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_218),
.A2(n_201),
.B1(n_196),
.B2(n_195),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_236),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_234),
.Y(n_242)
);

MAJx2_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_209),
.C(n_9),
.Y(n_234)
);

XNOR2x1_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_6),
.Y(n_235)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_238),
.B(n_225),
.Y(n_241)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_241),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_238),
.B(n_210),
.Y(n_244)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_244),
.Y(n_256)
);

A2O1A1Ixp33_ASAP7_75t_L g245 ( 
.A1(n_233),
.A2(n_215),
.B(n_219),
.C(n_213),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_245),
.A2(n_236),
.B(n_231),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_248),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_212),
.C(n_228),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_242),
.C(n_240),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_237),
.B(n_9),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_250),
.A2(n_252),
.B(n_11),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_243),
.A2(n_230),
.B1(n_235),
.B2(n_234),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_245),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_243),
.A2(n_228),
.B1(n_9),
.B2(n_11),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_257),
.C(n_5),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_249),
.C(n_242),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_258),
.A2(n_252),
.B1(n_4),
.B2(n_14),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_254),
.C(n_257),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_255),
.B(n_5),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_260),
.A2(n_261),
.B(n_262),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_4),
.Y(n_262)
);

AOI322xp5_ASAP7_75t_L g263 ( 
.A1(n_256),
.A2(n_4),
.A3(n_14),
.B1(n_13),
.B2(n_12),
.C1(n_15),
.C2(n_3),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_15),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_265),
.Y(n_270)
);

AO21x1_ASAP7_75t_L g271 ( 
.A1(n_267),
.A2(n_268),
.B(n_0),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_259),
.A2(n_15),
.B(n_1),
.Y(n_268)
);

OAI21x1_ASAP7_75t_L g269 ( 
.A1(n_266),
.A2(n_0),
.B(n_2),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_269),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_272),
.A2(n_270),
.B1(n_271),
.B2(n_3),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_3),
.C(n_0),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_2),
.Y(n_275)
);


endmodule