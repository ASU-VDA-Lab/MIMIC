module fake_netlist_1_8552_n_32 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_32);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_32;
wire n_20;
wire n_23;
wire n_8;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_2), .Y(n_8) );
INVx1_ASAP7_75t_SL g9 ( .A(n_1), .Y(n_9) );
OAI22xp5_ASAP7_75t_SL g10 ( .A1(n_7), .A2(n_2), .B1(n_6), .B2(n_4), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_5), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_3), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_11), .Y(n_13) );
AOI21xp5_ASAP7_75t_L g14 ( .A1(n_11), .A2(n_0), .B(n_3), .Y(n_14) );
INVx3_ASAP7_75t_L g15 ( .A(n_8), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_12), .B(n_5), .Y(n_16) );
NAND3xp33_ASAP7_75t_SL g17 ( .A(n_9), .B(n_0), .C(n_4), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_13), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_13), .Y(n_19) );
OR2x6_ASAP7_75t_L g20 ( .A(n_14), .B(n_10), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_20), .B(n_15), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_18), .Y(n_22) );
AND2x4_ASAP7_75t_L g23 ( .A(n_20), .B(n_15), .Y(n_23) );
INVx1_ASAP7_75t_SL g24 ( .A(n_21), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_22), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
AOI322xp5_ASAP7_75t_L g27 ( .A1(n_24), .A2(n_23), .A3(n_17), .B1(n_15), .B2(n_16), .C1(n_19), .C2(n_10), .Y(n_27) );
INVx2_ASAP7_75t_SL g28 ( .A(n_26), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_26), .Y(n_29) );
NOR2xp67_ASAP7_75t_L g30 ( .A(n_27), .B(n_23), .Y(n_30) );
HB1xp67_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
AOI22xp5_ASAP7_75t_SL g32 ( .A1(n_31), .A2(n_29), .B1(n_23), .B2(n_30), .Y(n_32) );
endmodule