module fake_jpeg_9113_n_279 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_279);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_181;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_128;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_33),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_37),
.Y(n_46)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_22),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_54),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_34),
.A2(n_16),
.B1(n_18),
.B2(n_25),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_39),
.A2(n_16),
.B1(n_34),
.B2(n_36),
.Y(n_64)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_50),
.Y(n_67)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_29),
.B(n_19),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_28),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_60),
.Y(n_77)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_53),
.A2(n_16),
.B1(n_18),
.B2(n_25),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_74),
.B1(n_36),
.B2(n_52),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_SL g90 ( 
.A(n_62),
.Y(n_90)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_66),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_64),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_65),
.Y(n_92)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_28),
.C(n_35),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_38),
.C(n_47),
.Y(n_91)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_71),
.Y(n_85)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_72),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_75),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_34),
.B1(n_36),
.B2(n_31),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_54),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_78),
.A2(n_93),
.B(n_97),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_80),
.A2(n_36),
.B1(n_48),
.B2(n_31),
.Y(n_106)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_82),
.Y(n_99)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_46),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_88),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_95),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_46),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_91),
.B(n_96),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_54),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_75),
.B(n_55),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_30),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_35),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_105),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_100),
.B(n_102),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_84),
.B(n_24),
.Y(n_102)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_107),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_56),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_106),
.A2(n_52),
.B1(n_33),
.B2(n_31),
.Y(n_128)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_108),
.A2(n_82),
.B1(n_92),
.B2(n_89),
.Y(n_137)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_111),
.Y(n_136)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

AND2x4_ASAP7_75t_SL g112 ( 
.A(n_78),
.B(n_50),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_112),
.A2(n_93),
.B(n_97),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_87),
.A2(n_52),
.B1(n_31),
.B2(n_70),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_89),
.B1(n_79),
.B2(n_14),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_56),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_115),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_60),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_97),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_42),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_57),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_118),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_57),
.Y(n_119)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_122),
.B(n_124),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_99),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_106),
.A2(n_87),
.B1(n_91),
.B2(n_78),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_125),
.A2(n_127),
.B1(n_140),
.B2(n_113),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_126),
.A2(n_131),
.B(n_139),
.Y(n_145)
);

AO22x1_ASAP7_75t_SL g127 ( 
.A1(n_112),
.A2(n_93),
.B1(n_80),
.B2(n_33),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_SL g148 ( 
.A1(n_128),
.A2(n_137),
.B(n_108),
.C(n_104),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_110),
.B(n_29),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_132),
.Y(n_164)
);

NAND2xp33_ASAP7_75t_SL g131 ( 
.A(n_112),
.B(n_33),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_41),
.C(n_95),
.Y(n_132)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_111),
.Y(n_151)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_135),
.B(n_142),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_110),
.A2(n_37),
.B(n_19),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_118),
.Y(n_143)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_101),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_143),
.B(n_159),
.Y(n_176)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_153),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_117),
.Y(n_147)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_148),
.A2(n_116),
.B1(n_108),
.B2(n_104),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_112),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_150),
.A2(n_126),
.B(n_139),
.Y(n_167)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_156),
.Y(n_173)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_136),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_117),
.Y(n_154)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_117),
.Y(n_155)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

XOR2x2_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_112),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_157),
.A2(n_110),
.B(n_125),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_103),
.Y(n_158)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_121),
.B(n_102),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_140),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_165),
.Y(n_184)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_162),
.Y(n_177)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_163),
.A2(n_131),
.B1(n_115),
.B2(n_105),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_120),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_98),
.Y(n_166)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_167),
.A2(n_175),
.B(n_143),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_129),
.C(n_132),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_164),
.C(n_145),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_149),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_155),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_145),
.A2(n_122),
.B(n_123),
.Y(n_175)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_98),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_182),
.A2(n_185),
.B(n_76),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_163),
.A2(n_120),
.B1(n_116),
.B2(n_113),
.Y(n_183)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_183),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_162),
.A2(n_114),
.B1(n_101),
.B2(n_107),
.Y(n_186)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_186),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_187),
.A2(n_156),
.B1(n_161),
.B2(n_150),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_157),
.A2(n_109),
.B1(n_98),
.B2(n_20),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_188),
.A2(n_21),
.B1(n_20),
.B2(n_158),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_189),
.A2(n_198),
.B1(n_172),
.B2(n_169),
.Y(n_214)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_177),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_196),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_184),
.A2(n_153),
.B1(n_152),
.B2(n_148),
.Y(n_193)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_195),
.A2(n_207),
.B(n_175),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_197),
.B(n_200),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_148),
.B1(n_154),
.B2(n_147),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_199),
.Y(n_220)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_201),
.B(n_203),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_168),
.C(n_185),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_187),
.A2(n_150),
.B1(n_148),
.B2(n_146),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_204),
.A2(n_174),
.B1(n_172),
.B2(n_169),
.Y(n_212)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_205),
.A2(n_206),
.B1(n_181),
.B2(n_171),
.Y(n_210)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_218),
.C(n_204),
.Y(n_225)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

NAND3xp33_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_188),
.C(n_167),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_214),
.Y(n_226)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_178),
.C(n_174),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_217),
.C(n_219),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_178),
.C(n_92),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_65),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_62),
.C(n_76),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_191),
.A2(n_24),
.B1(n_21),
.B2(n_22),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_223),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_237),
.C(n_219),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_190),
.C(n_203),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_235),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_215),
.A2(n_201),
.B1(n_196),
.B2(n_14),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_232),
.A2(n_222),
.B(n_220),
.Y(n_242)
);

BUFx24_ASAP7_75t_SL g233 ( 
.A(n_210),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_236),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_208),
.A2(n_15),
.B1(n_26),
.B2(n_8),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_234),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_27),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_27),
.C(n_23),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_7),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_244),
.C(n_245),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_226),
.A2(n_216),
.B(n_224),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_241),
.B(n_249),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_248),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_209),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_228),
.A2(n_212),
.B(n_8),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_250),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_27),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_229),
.A2(n_7),
.B(n_12),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_27),
.C(n_23),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_239),
.A2(n_236),
.B1(n_232),
.B2(n_237),
.Y(n_252)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_243),
.B(n_26),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_255),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_240),
.A2(n_6),
.B1(n_10),
.B2(n_7),
.Y(n_255)
);

INVxp33_ASAP7_75t_SL g257 ( 
.A(n_244),
.Y(n_257)
);

AOI21xp33_ASAP7_75t_L g267 ( 
.A1(n_257),
.A2(n_258),
.B(n_6),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_248),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_23),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_256),
.Y(n_262)
);

OAI21xp33_ASAP7_75t_L g271 ( 
.A1(n_262),
.A2(n_0),
.B(n_1),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_251),
.A2(n_26),
.B1(n_15),
.B2(n_5),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_265),
.Y(n_268)
);

AO21x1_ASAP7_75t_L g264 ( 
.A1(n_254),
.A2(n_5),
.B(n_6),
.Y(n_264)
);

MAJx2_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_267),
.C(n_10),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_5),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_270),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_261),
.A2(n_260),
.B(n_266),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_271),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_272),
.B(n_266),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_274),
.A2(n_273),
.B(n_268),
.Y(n_275)
);

AOI21x1_ASAP7_75t_L g276 ( 
.A1(n_275),
.A2(n_1),
.B(n_2),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_1),
.C(n_2),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_2),
.B1(n_3),
.B2(n_272),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_3),
.Y(n_279)
);


endmodule