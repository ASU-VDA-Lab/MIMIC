module fake_jpeg_16054_n_86 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_86);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_86;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

BUFx2_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_17),
.B(n_20),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_22),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_10),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_16),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_13),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_8),
.B(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

OAI32xp33_ASAP7_75t_L g30 ( 
.A1(n_23),
.A2(n_17),
.A3(n_13),
.B1(n_12),
.B2(n_15),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_30),
.A2(n_34),
.B1(n_9),
.B2(n_10),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_23),
.B(n_19),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_14),
.Y(n_42)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_37),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_26),
.A2(n_11),
.B1(n_12),
.B2(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_10),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_19),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_1),
.B(n_2),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_32),
.B(n_6),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_SL g50 ( 
.A(n_46),
.B(n_47),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_25),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_22),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_9),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_SL g51 ( 
.A1(n_48),
.A2(n_30),
.B(n_25),
.C(n_33),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_51),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_36),
.B1(n_6),
.B2(n_3),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_53),
.C(n_47),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_19),
.C(n_22),
.Y(n_53)
);

NAND3xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_36),
.C(n_2),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_55),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_1),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_59),
.Y(n_64)
);

FAx1_ASAP7_75t_SL g71 ( 
.A(n_60),
.B(n_4),
.CI(n_5),
.CON(n_71),
.SN(n_71)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

OA21x2_ASAP7_75t_SL g67 ( 
.A1(n_63),
.A2(n_51),
.B(n_56),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_45),
.C(n_4),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_1),
.Y(n_69)
);

INVxp33_ASAP7_75t_SL g72 ( 
.A(n_67),
.Y(n_72)
);

FAx1_ASAP7_75t_SL g68 ( 
.A(n_61),
.B(n_56),
.CI(n_51),
.CON(n_68),
.SN(n_68)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_66),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_71),
.Y(n_75)
);

NOR2xp67_ASAP7_75t_SL g73 ( 
.A(n_67),
.B(n_62),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_68),
.Y(n_78)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_75),
.B(n_70),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_77),
.B(n_68),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_68),
.C(n_71),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_72),
.B(n_70),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_79),
.A2(n_81),
.B(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_82),
.A2(n_78),
.B1(n_71),
.B2(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_83),
.Y(n_86)
);


endmodule