module fake_jpeg_722_n_513 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_513);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_513;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_341;
wire n_151;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_SL g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_49),
.Y(n_117)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_51),
.Y(n_119)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_54),
.Y(n_132)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g162 ( 
.A(n_56),
.Y(n_162)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_59),
.B(n_77),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_61),
.B(n_68),
.Y(n_121)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_62),
.Y(n_140)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_65),
.Y(n_142)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_27),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_20),
.B(n_0),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_70),
.Y(n_147)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_73),
.Y(n_151)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_75),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_20),
.B(n_0),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_76),
.B(n_80),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_37),
.B(n_1),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_78),
.Y(n_155)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

CKINVDCx6p67_ASAP7_75t_R g144 ( 
.A(n_79),
.Y(n_144)
);

BUFx4f_ASAP7_75t_SL g80 ( 
.A(n_27),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_81),
.Y(n_156)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_15),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_83),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_84),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_15),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_85),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_87),
.Y(n_159)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_89),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_14),
.B(n_1),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_92),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

BUFx10_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_14),
.B(n_1),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_15),
.Y(n_96)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_15),
.Y(n_97)
);

BUFx10_ASAP7_75t_L g158 ( 
.A(n_97),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_100),
.Y(n_163)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_101),
.B(n_35),
.Y(n_146)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_36),
.B1(n_64),
.B2(n_70),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_29),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_35),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_61),
.A2(n_30),
.B1(n_42),
.B2(n_29),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_104),
.A2(n_33),
.B1(n_17),
.B2(n_16),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_92),
.A2(n_36),
.B1(n_42),
.B2(n_29),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_120),
.A2(n_139),
.B1(n_154),
.B2(n_161),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_146),
.Y(n_168)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_68),
.B(n_42),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_133),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_76),
.A2(n_36),
.B1(n_42),
.B2(n_35),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_83),
.A2(n_41),
.B1(n_38),
.B2(n_34),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_150),
.A2(n_44),
.B1(n_16),
.B2(n_13),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_85),
.A2(n_35),
.B1(n_32),
.B2(n_41),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_47),
.A2(n_32),
.B1(n_38),
.B2(n_18),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_49),
.A2(n_32),
.B1(n_18),
.B2(n_33),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_44),
.B1(n_33),
.B2(n_25),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_166),
.B(n_167),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_115),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_169),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_144),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_170),
.B(n_172),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_144),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_171),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_110),
.B(n_1),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_1),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_173),
.B(n_182),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_174),
.Y(n_235)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_175),
.Y(n_242)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_177),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_121),
.B(n_67),
.C(n_96),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_178),
.B(n_185),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_113),
.Y(n_179)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_111),
.Y(n_180)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_180),
.Y(n_232)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_181),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_121),
.B(n_2),
.Y(n_182)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_117),
.Y(n_183)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_183),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_161),
.A2(n_164),
.B1(n_118),
.B2(n_154),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_184),
.A2(n_190),
.B1(n_199),
.B2(n_206),
.Y(n_225)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_140),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_126),
.B(n_2),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_186),
.B(n_201),
.Y(n_247)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_137),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_127),
.Y(n_188)
);

NOR3xp33_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_194),
.C(n_196),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_126),
.B(n_2),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_192),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_105),
.B(n_2),
.Y(n_192)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_193),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_159),
.B(n_2),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_152),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_195),
.Y(n_228)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_128),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_106),
.B(n_79),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_197),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_141),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_198),
.Y(n_233)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_143),
.Y(n_200)
);

INVx11_ASAP7_75t_L g241 ( 
.A(n_200),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_107),
.B(n_80),
.Y(n_201)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_148),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_202),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_114),
.A2(n_94),
.B1(n_84),
.B2(n_98),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_203),
.A2(n_204),
.B1(n_207),
.B2(n_25),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_132),
.B(n_25),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_208),
.Y(n_231)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_141),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_135),
.A2(n_103),
.B1(n_51),
.B2(n_95),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_142),
.Y(n_208)
);

AND2x2_ASAP7_75t_SL g209 ( 
.A(n_155),
.B(n_74),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_211),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_116),
.Y(n_210)
);

OA22x2_ASAP7_75t_L g212 ( 
.A1(n_210),
.A2(n_17),
.B1(n_46),
.B2(n_44),
.Y(n_212)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_109),
.Y(n_211)
);

INVx11_ASAP7_75t_L g267 ( 
.A(n_212),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_173),
.B(n_160),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_214),
.B(n_210),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_216),
.A2(n_230),
.B1(n_236),
.B2(n_237),
.Y(n_249)
);

AOI32xp33_ASAP7_75t_L g224 ( 
.A1(n_191),
.A2(n_156),
.A3(n_147),
.B1(n_112),
.B2(n_163),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_176),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_168),
.A2(n_122),
.B1(n_136),
.B2(n_58),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_165),
.A2(n_130),
.B1(n_119),
.B2(n_125),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_168),
.A2(n_130),
.B1(n_119),
.B2(n_125),
.Y(n_237)
);

A2O1A1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_182),
.A2(n_13),
.B(n_16),
.C(n_17),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_244),
.B(n_245),
.Y(n_256)
);

A2O1A1Ixp33_ASAP7_75t_L g245 ( 
.A1(n_178),
.A2(n_46),
.B(n_13),
.C(n_109),
.Y(n_245)
);

A2O1A1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_189),
.A2(n_46),
.B(n_162),
.C(n_43),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_209),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_248),
.A2(n_250),
.B(n_254),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_234),
.A2(n_176),
.B1(n_184),
.B2(n_168),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_209),
.C(n_197),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_251),
.B(n_252),
.C(n_255),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_197),
.C(n_192),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_218),
.Y(n_253)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_253),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_223),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_218),
.Y(n_257)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

BUFx24_ASAP7_75t_SL g258 ( 
.A(n_247),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_258),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_227),
.B(n_205),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_259),
.B(n_261),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_223),
.B(n_195),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_264),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_208),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_225),
.A2(n_204),
.B1(n_145),
.B2(n_149),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_262),
.A2(n_269),
.B1(n_270),
.B2(n_237),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_263),
.B(n_265),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_167),
.C(n_166),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_214),
.B(n_245),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_244),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_266),
.B(n_274),
.Y(n_297)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_218),
.Y(n_268)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_268),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_236),
.A2(n_196),
.B1(n_183),
.B2(n_193),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_216),
.A2(n_181),
.B1(n_200),
.B2(n_149),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_219),
.B(n_198),
.C(n_177),
.Y(n_271)
);

MAJx2_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_273),
.C(n_215),
.Y(n_295)
);

INVx11_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_272),
.A2(n_243),
.B1(n_171),
.B2(n_174),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_215),
.B(n_210),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_242),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_230),
.A2(n_187),
.B1(n_145),
.B2(n_131),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_275),
.A2(n_243),
.B1(n_239),
.B2(n_228),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_175),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_212),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_248),
.B(n_238),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_277),
.Y(n_320)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_279),
.Y(n_307)
);

AND2x6_ASAP7_75t_L g280 ( 
.A(n_250),
.B(n_224),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_280),
.B(n_300),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_246),
.B(n_238),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_282),
.A2(n_288),
.B(n_306),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_267),
.A2(n_219),
.B1(n_217),
.B2(n_246),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_284),
.A2(n_301),
.B1(n_272),
.B2(n_235),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_267),
.A2(n_217),
.B1(n_233),
.B2(n_242),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_285),
.A2(n_287),
.B1(n_294),
.B2(n_262),
.Y(n_321)
);

INVxp33_ASAP7_75t_L g286 ( 
.A(n_276),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_286),
.B(n_212),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_249),
.A2(n_247),
.B1(n_233),
.B2(n_239),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_251),
.B(n_222),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_256),
.Y(n_291)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_291),
.Y(n_332)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_253),
.Y(n_292)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_292),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_295),
.B(n_264),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_254),
.A2(n_229),
.B1(n_228),
.B2(n_242),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_296),
.A2(n_275),
.B1(n_274),
.B2(n_226),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_256),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_299),
.B(n_273),
.Y(n_322)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_257),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_267),
.A2(n_229),
.B1(n_179),
.B2(n_202),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_302),
.Y(n_315)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_268),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_261),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_278),
.B(n_255),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_309),
.B(n_314),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_252),
.C(n_260),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_310),
.B(n_309),
.C(n_313),
.Y(n_343)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_311),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_252),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_313),
.B(n_316),
.Y(n_352)
);

MAJx2_ASAP7_75t_L g314 ( 
.A(n_278),
.B(n_295),
.C(n_289),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_295),
.B(n_260),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_259),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_317),
.B(n_318),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_297),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_277),
.B(n_264),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_319),
.B(n_220),
.Y(n_362)
);

OA22x2_ASAP7_75t_L g359 ( 
.A1(n_321),
.A2(n_290),
.B1(n_283),
.B2(n_281),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_322),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_323),
.B(n_290),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_293),
.B(n_265),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_324),
.B(n_327),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_287),
.A2(n_249),
.B1(n_270),
.B2(n_269),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_325),
.A2(n_328),
.B1(n_331),
.B2(n_333),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_297),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_326),
.B(n_329),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_303),
.B(n_263),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_301),
.Y(n_329)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_330),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_291),
.A2(n_271),
.B1(n_221),
.B2(n_240),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_293),
.B(n_213),
.Y(n_334)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_334),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_294),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_336),
.A2(n_283),
.B(n_305),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_315),
.A2(n_299),
.B(n_289),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_338),
.A2(n_340),
.B(n_341),
.Y(n_378)
);

AOI22x1_ASAP7_75t_L g339 ( 
.A1(n_308),
.A2(n_285),
.B1(n_282),
.B2(n_284),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_339),
.A2(n_350),
.B1(n_365),
.B2(n_366),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_312),
.A2(n_302),
.B(n_296),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_326),
.A2(n_277),
.B(n_280),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_343),
.B(n_354),
.C(n_356),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_323),
.B(n_277),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_345),
.B(n_220),
.Y(n_382)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_335),
.Y(n_348)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_348),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_336),
.A2(n_279),
.B1(n_280),
.B2(n_288),
.Y(n_350)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_351),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_310),
.B(n_288),
.C(n_300),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_335),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g393 ( 
.A1(n_355),
.A2(n_358),
.B1(n_363),
.B2(n_241),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_314),
.B(n_288),
.C(n_292),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_357),
.B(n_360),
.C(n_362),
.Y(n_387)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_311),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_359),
.B(n_328),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_319),
.B(n_281),
.C(n_226),
.Y(n_360)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_318),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_307),
.A2(n_221),
.B1(n_240),
.B2(n_306),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_307),
.A2(n_321),
.B1(n_332),
.B2(n_312),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_368),
.B(n_373),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_361),
.B(n_317),
.Y(n_369)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_369),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_342),
.A2(n_308),
.B1(n_332),
.B2(n_325),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_370),
.A2(n_374),
.B1(n_376),
.B2(n_362),
.Y(n_396)
);

OR2x4_ASAP7_75t_L g371 ( 
.A(n_340),
.B(n_320),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_371),
.Y(n_395)
);

BUFx12_ASAP7_75t_L g372 ( 
.A(n_351),
.Y(n_372)
);

CKINVDCx14_ASAP7_75t_R g405 ( 
.A(n_372),
.Y(n_405)
);

CKINVDCx14_ASAP7_75t_R g373 ( 
.A(n_344),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_342),
.A2(n_320),
.B1(n_329),
.B2(n_331),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_347),
.B(n_346),
.Y(n_375)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_375),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_366),
.A2(n_324),
.B1(n_333),
.B2(n_316),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_347),
.B(n_212),
.Y(n_377)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_377),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_359),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_379),
.B(n_391),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_359),
.B(n_212),
.Y(n_381)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_381),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_382),
.B(n_392),
.Y(n_398)
);

AOI322xp5_ASAP7_75t_L g384 ( 
.A1(n_338),
.A2(n_272),
.A3(n_221),
.B1(n_158),
.B2(n_131),
.C1(n_153),
.C2(n_148),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_384),
.B(n_385),
.Y(n_397)
);

BUFx12_ASAP7_75t_L g385 ( 
.A(n_339),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_354),
.B(n_157),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_386),
.B(n_393),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_364),
.B(n_232),
.Y(n_388)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_388),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_353),
.B(n_232),
.Y(n_389)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_389),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_349),
.B(n_235),
.Y(n_391)
);

OAI32xp33_ASAP7_75t_L g392 ( 
.A1(n_339),
.A2(n_241),
.A3(n_185),
.B1(n_235),
.B2(n_123),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_390),
.A2(n_350),
.B1(n_341),
.B2(n_359),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_394),
.A2(n_404),
.B1(n_416),
.B2(n_374),
.Y(n_419)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_396),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_367),
.A2(n_337),
.B1(n_356),
.B2(n_357),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_399),
.B(n_415),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_390),
.A2(n_365),
.B1(n_348),
.B2(n_360),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_383),
.B(n_343),
.C(n_352),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_406),
.B(n_412),
.C(n_417),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_378),
.A2(n_345),
.B(n_352),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_409),
.A2(n_369),
.B(n_375),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_383),
.B(n_337),
.C(n_157),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_392),
.B(n_102),
.Y(n_414)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_414),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_386),
.B(n_211),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_376),
.A2(n_86),
.B1(n_75),
.B2(n_69),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_387),
.B(n_180),
.C(n_124),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_419),
.B(n_397),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_405),
.A2(n_378),
.B(n_371),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_420),
.A2(n_433),
.B(n_417),
.Y(n_442)
);

MAJx2_ASAP7_75t_L g440 ( 
.A(n_421),
.B(n_394),
.C(n_398),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_SL g423 ( 
.A(n_409),
.B(n_396),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_423),
.B(n_408),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_402),
.B(n_380),
.Y(n_424)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_424),
.Y(n_454)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_401),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_425),
.B(n_427),
.Y(n_446)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_401),
.Y(n_427)
);

INVxp33_ASAP7_75t_L g428 ( 
.A(n_413),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_428),
.A2(n_430),
.B1(n_435),
.B2(n_438),
.Y(n_455)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_400),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_402),
.B(n_380),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_431),
.A2(n_437),
.B(n_377),
.Y(n_451)
);

OR2x2_ASAP7_75t_L g432 ( 
.A(n_403),
.B(n_391),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_432),
.A2(n_381),
.B1(n_414),
.B2(n_385),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_410),
.B(n_387),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_406),
.B(n_382),
.C(n_370),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_434),
.B(n_436),
.Y(n_448)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_407),
.Y(n_435)
);

BUFx24_ASAP7_75t_SL g436 ( 
.A(n_395),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_395),
.B(n_379),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_404),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_439),
.A2(n_442),
.B1(n_452),
.B2(n_437),
.Y(n_464)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_440),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_422),
.B(n_412),
.C(n_411),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_441),
.B(n_443),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_422),
.B(n_411),
.C(n_399),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_434),
.B(n_398),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_444),
.B(n_447),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_445),
.B(n_153),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_418),
.B(n_415),
.C(n_368),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_418),
.B(n_416),
.C(n_372),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_449),
.B(n_451),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_429),
.A2(n_414),
.B1(n_385),
.B2(n_372),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_450),
.A2(n_426),
.B1(n_162),
.B2(n_151),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_421),
.B(n_241),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_453),
.B(n_52),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_423),
.B(n_158),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_456),
.B(n_426),
.Y(n_467)
);

INVx6_ASAP7_75t_L g457 ( 
.A(n_428),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_457),
.B(n_432),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_454),
.A2(n_429),
.B1(n_431),
.B2(n_424),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_458),
.A2(n_464),
.B1(n_472),
.B2(n_457),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_441),
.B(n_419),
.C(n_420),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_459),
.B(n_462),
.Y(n_484)
);

BUFx24_ASAP7_75t_SL g461 ( 
.A(n_448),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_461),
.B(n_463),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_439),
.B(n_444),
.C(n_443),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_467),
.B(n_473),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_468),
.B(n_471),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_449),
.B(n_72),
.C(n_158),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_470),
.B(n_462),
.C(n_465),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_446),
.A2(n_32),
.B1(n_88),
.B2(n_62),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_475),
.A2(n_472),
.B1(n_4),
.B2(n_5),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_469),
.A2(n_447),
.B(n_445),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_476),
.A2(n_485),
.B(n_474),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_477),
.B(n_480),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_460),
.B(n_455),
.C(n_440),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_479),
.B(n_481),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_459),
.B(n_453),
.C(n_450),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_466),
.B(n_3),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_482),
.B(n_486),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_458),
.A2(n_153),
.B(n_43),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_483),
.A2(n_3),
.B(n_5),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_471),
.A2(n_43),
.B(n_23),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_470),
.B(n_43),
.C(n_23),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_484),
.B(n_473),
.Y(n_487)
);

AO21x1_ASAP7_75t_L g497 ( 
.A1(n_487),
.A2(n_496),
.B(n_474),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_490),
.Y(n_498)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_491),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_477),
.B(n_3),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_492),
.B(n_493),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_478),
.B(n_12),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_476),
.B(n_12),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_494),
.B(n_11),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_495),
.A2(n_485),
.B(n_6),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_497),
.B(n_500),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_502),
.B(n_5),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_504),
.A2(n_505),
.B(n_506),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_498),
.B(n_488),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_501),
.A2(n_487),
.B(n_489),
.Y(n_506)
);

AO221x1_ASAP7_75t_L g507 ( 
.A1(n_503),
.A2(n_499),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_507),
.B(n_5),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_509),
.B(n_7),
.Y(n_510)
);

AO21x1_ASAP7_75t_L g511 ( 
.A1(n_510),
.A2(n_508),
.B(n_10),
.Y(n_511)
);

MAJx2_ASAP7_75t_L g512 ( 
.A(n_511),
.B(n_9),
.C(n_10),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_512),
.A2(n_10),
.B(n_11),
.Y(n_513)
);


endmodule