module real_jpeg_28757_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_176;
wire n_221;
wire n_166;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_191;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_202;
wire n_244;
wire n_128;
wire n_179;
wire n_167;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

INVx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_1),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_1),
.A2(n_3),
.B(n_57),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_1),
.A2(n_60),
.B1(n_61),
.B2(n_142),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_1),
.B(n_38),
.Y(n_202)
);

A2O1A1O1Ixp25_ASAP7_75t_L g204 ( 
.A1(n_1),
.A2(n_38),
.B(n_42),
.C(n_202),
.D(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_1),
.B(n_71),
.Y(n_209)
);

OAI21xp33_ASAP7_75t_L g233 ( 
.A1(n_1),
.A2(n_24),
.B(n_215),
.Y(n_233)
);

A2O1A1O1Ixp25_ASAP7_75t_L g243 ( 
.A1(n_1),
.A2(n_58),
.B(n_70),
.C(n_154),
.D(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_1),
.B(n_58),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_2),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_2),
.A2(n_40),
.B1(n_57),
.B2(n_58),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_2),
.A2(n_25),
.B1(n_29),
.B2(n_40),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_3),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_3),
.A2(n_56),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_4),
.A2(n_60),
.B1(n_61),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_4),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_4),
.A2(n_57),
.B1(n_58),
.B2(n_67),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_4),
.A2(n_38),
.B1(n_39),
.B2(n_67),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_4),
.A2(n_25),
.B1(n_29),
.B2(n_67),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_6),
.A2(n_60),
.B1(n_61),
.B2(n_98),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_6),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_6),
.A2(n_57),
.B1(n_58),
.B2(n_98),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_6),
.A2(n_38),
.B1(n_39),
.B2(n_98),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_6),
.A2(n_25),
.B1(n_29),
.B2(n_98),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_7),
.A2(n_38),
.B1(n_39),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_7),
.A2(n_25),
.B1(n_29),
.B2(n_48),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_7),
.A2(n_48),
.B1(n_57),
.B2(n_58),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_8),
.A2(n_57),
.B1(n_58),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_8),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_8),
.A2(n_38),
.B1(n_39),
.B2(n_77),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_8),
.A2(n_60),
.B1(n_61),
.B2(n_77),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_8),
.A2(n_25),
.B1(n_29),
.B2(n_77),
.Y(n_191)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_10),
.A2(n_60),
.B1(n_61),
.B2(n_64),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_10),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_10),
.A2(n_57),
.B1(n_58),
.B2(n_64),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_10),
.A2(n_25),
.B1(n_29),
.B2(n_64),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_10),
.A2(n_38),
.B1(n_39),
.B2(n_64),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_11),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_11),
.A2(n_30),
.B1(n_38),
.B2(n_39),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_12),
.A2(n_38),
.B(n_43),
.C(n_44),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_12),
.B(n_38),
.Y(n_43)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_13),
.A2(n_25),
.B1(n_29),
.B2(n_35),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_13),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_109)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_15),
.A2(n_38),
.B1(n_39),
.B2(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_15),
.Y(n_74)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_16),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_127),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_125),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_104),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_20),
.B(n_104),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_81),
.C(n_88),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_21),
.B(n_81),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_50),
.B1(n_51),
.B2(n_80),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_22),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_23),
.B(n_36),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B1(n_31),
.B2(n_34),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_24),
.A2(n_31),
.B(n_34),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_24),
.A2(n_28),
.B1(n_91),
.B2(n_93),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_24),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_24),
.A2(n_93),
.B1(n_148),
.B2(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_24),
.A2(n_214),
.B(n_215),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_24),
.B(n_217),
.Y(n_231)
);

NAND2x1_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_27),
.Y(n_24)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_25),
.A2(n_29),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_25),
.B(n_46),
.Y(n_203)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI32xp33_ASAP7_75t_L g201 ( 
.A1(n_29),
.A2(n_39),
.A3(n_45),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_29),
.B(n_235),
.Y(n_234)
);

INVx5_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_32),
.A2(n_92),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_32),
.B(n_216),
.Y(n_215)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_33),
.B(n_142),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_47),
.B2(n_49),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_37),
.A2(n_41),
.B1(n_49),
.B2(n_95),
.Y(n_94)
);

AOI32xp33_ASAP7_75t_L g251 ( 
.A1(n_38),
.A2(n_57),
.A3(n_244),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_SL g253 ( 
.A(n_39),
.B(n_75),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_41),
.A2(n_263),
.B(n_264),
.Y(n_262)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_42),
.A2(n_44),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_42),
.A2(n_44),
.B1(n_85),
.B2(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_42),
.B(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_42),
.A2(n_44),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_47),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_49),
.A2(n_95),
.B(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_49),
.B(n_170),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_49),
.A2(n_168),
.B(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_49),
.B(n_142),
.Y(n_228)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_68),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_52),
.B(n_68),
.C(n_80),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_62),
.B(n_65),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_54),
.A2(n_55),
.B1(n_63),
.B2(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_54),
.B(n_66),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_54),
.A2(n_172),
.B(n_173),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_59),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_55),
.B(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_56),
.A2(n_60),
.B(n_142),
.C(n_143),
.Y(n_141)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_57),
.A2(n_58),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_65),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_76),
.B1(n_78),
.B2(n_79),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_69),
.A2(n_151),
.B(n_153),
.Y(n_150)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_70),
.B(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_70),
.A2(n_71),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_70),
.A2(n_71),
.B1(n_152),
.B2(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_73),
.Y(n_70)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_75),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_78),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_78),
.B(n_103),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_78),
.A2(n_101),
.B(n_176),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_79),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_86),
.B2(n_87),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_87),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_87),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_88),
.B(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_96),
.C(n_99),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_89),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_90),
.B(n_94),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_93),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_93),
.A2(n_222),
.B(n_230),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_96),
.A2(n_99),
.B1(n_100),
.B2(n_132),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_96),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_97),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_124),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_114),
.B1(n_115),
.B2(n_123),
.Y(n_105)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_110),
.B(n_113),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_110),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_122),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_120),
.B(n_121),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_121),
.B(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_119),
.B(n_142),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_157),
.B(n_273),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_155),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_129),
.B(n_155),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.C(n_134),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_130),
.B(n_133),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_134),
.A2(n_135),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.C(n_149),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_136),
.A2(n_137),
.B1(n_149),
.B2(n_150),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_140),
.A2(n_141),
.B1(n_144),
.B2(n_145),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_146),
.A2(n_221),
.B1(n_223),
.B2(n_224),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_194),
.Y(n_157)
);

INVxp33_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_180),
.B(n_193),
.Y(n_159)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_160),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_177),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_161),
.B(n_177),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.C(n_165),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_165),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_171),
.C(n_174),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_166),
.A2(n_167),
.B1(n_174),
.B2(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_171),
.B(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_174),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_178),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_181),
.B(n_183),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.C(n_188),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_184),
.B(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_187),
.B(n_188),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.C(n_192),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_189),
.B(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_190),
.B(n_192),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_191),
.Y(n_250)
);

NOR3xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_271),
.C(n_272),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_266),
.B(n_270),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_255),
.B(n_265),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_239),
.B(n_254),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_218),
.B(n_238),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_206),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_200),
.B(n_206),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_204),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_205),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_213),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_211),
.C(n_213),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_212),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_214),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_226),
.B(n_237),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_225),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_220),
.B(n_225),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_224),
.A2(n_231),
.B(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_232),
.B(n_236),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_228),
.B(n_229),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_240),
.B(n_241),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_248),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_245),
.C(n_248),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_247),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_251),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_256),
.B(n_257),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_261),
.C(n_262),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_267),
.B(n_268),
.Y(n_270)
);


endmodule