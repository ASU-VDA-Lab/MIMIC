module real_jpeg_5006_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_164;
wire n_48;
wire n_184;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_97;
wire n_75;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_1),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_2),
.A2(n_66),
.B1(n_70),
.B2(n_71),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_2),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_2),
.A2(n_70),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_4),
.Y(n_77)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_4),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_4),
.Y(n_146)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_5),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_6),
.B(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_6),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_6),
.B(n_122),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_6),
.A2(n_29),
.B1(n_119),
.B2(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_6),
.B(n_170),
.C(n_171),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_6),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_6),
.B(n_164),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_7),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_7),
.A2(n_38),
.B1(n_86),
.B2(n_90),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_7),
.A2(n_38),
.B1(n_128),
.B2(n_131),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_8),
.A2(n_139),
.B1(n_141),
.B2(n_142),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_8),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_9),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_9),
.A2(n_31),
.B1(n_187),
.B2(n_192),
.Y(n_186)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_10),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_157),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_155),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_92),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_14),
.B(n_92),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_53),
.C(n_64),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_15),
.A2(n_16),
.B1(n_53),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_28),
.B(n_33),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_17),
.A2(n_28),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_17),
.Y(n_164)
);

AOI22x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx3_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_22),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_23),
.Y(n_194)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_24),
.Y(n_172)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_30),
.Y(n_168)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

NAND2xp33_ASAP7_75t_SL g153 ( 
.A(n_32),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_43),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_34),
.B(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_42),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_43),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_50),
.B2(n_52),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx5_ASAP7_75t_SL g151 ( 
.A(n_52),
.Y(n_151)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_53),
.Y(n_175)
);

OR2x2_ASAP7_75t_SL g104 ( 
.A(n_54),
.B(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_54),
.Y(n_134)
);

AO22x2_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_57),
.Y(n_152)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_64),
.B(n_174),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_74),
.B(n_81),
.Y(n_64)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_65),
.Y(n_200)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_69),
.Y(n_191)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_73),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_74),
.A2(n_81),
.B(n_119),
.Y(n_183)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_75),
.B(n_85),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_75),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_77),
.Y(n_182)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_77),
.Y(n_202)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_78),
.Y(n_180)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx8_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_83),
.A2(n_147),
.B(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_135),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_101),
.B2(n_102),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_96),
.A2(n_161),
.B(n_163),
.Y(n_160)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_115),
.B(n_126),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_112),
.B2(n_113),
.Y(n_105)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_111),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_119),
.B(n_120),
.Y(n_115)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVxp33_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI32xp33_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_149),
.A3(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_148)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_134),
.Y(n_126)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_148),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_144),
.B(n_147),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_SL g149 ( 
.A(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_176),
.B(n_206),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_173),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_159),
.B(n_173),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_165),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_160),
.A2(n_165),
.B1(n_166),
.B2(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_197),
.B(n_205),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_184),
.B(n_196),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_195),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_195),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_186),
.Y(n_199)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_203),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_203),
.Y(n_205)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);


endmodule