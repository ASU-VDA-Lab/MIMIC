module fake_ibex_427_n_923 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_923);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_923;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_708;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_859;
wire n_259;
wire n_276;
wire n_470;
wire n_339;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_469;
wire n_323;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_732;
wire n_673;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_538;
wire n_464;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_636;
wire n_594;
wire n_710;
wire n_720;
wire n_490;
wire n_407;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_580;
wire n_543;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_857;
wire n_849;
wire n_765;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_472;
wire n_229;
wire n_209;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_704;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_869;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_392;
wire n_354;
wire n_206;
wire n_630;
wire n_567;
wire n_548;
wire n_516;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_444;
wire n_200;
wire n_562;
wire n_506;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_285;
wire n_247;
wire n_320;
wire n_379;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_890;
wire n_874;
wire n_816;
wire n_912;
wire n_921;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g178 ( 
.A(n_45),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_153),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_85),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_77),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_52),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_9),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_137),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_86),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_44),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_53),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_19),
.Y(n_189)
);

BUFx2_ASAP7_75t_SL g190 ( 
.A(n_24),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_139),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_67),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_72),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_113),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_120),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_155),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_38),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_98),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_150),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_146),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_78),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_136),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_94),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_80),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_56),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_177),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_90),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_142),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_87),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_11),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_121),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_133),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_89),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_40),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_61),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_176),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_123),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_99),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_115),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_48),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_124),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_143),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_169),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_160),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_75),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_39),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_166),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_126),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_81),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_104),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_74),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_30),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_28),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_58),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_55),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_70),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_63),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_20),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_158),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_154),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_165),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_156),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_68),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_49),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_128),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_101),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_161),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_23),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_119),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_145),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_174),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_91),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_28),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_9),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_122),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_51),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_57),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_42),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_96),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_130),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_138),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_46),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_149),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_95),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_16),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_31),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_148),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_173),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_32),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_50),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_62),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_73),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_60),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_6),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_127),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_54),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_131),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_141),
.B(n_102),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_66),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_2),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_140),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_37),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_33),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_13),
.Y(n_284)
);

INVxp67_ASAP7_75t_SL g285 ( 
.A(n_47),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_25),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_17),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_33),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_144),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_5),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_83),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_225),
.B(n_34),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_223),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_214),
.Y(n_294)
);

AND2x4_ASAP7_75t_L g295 ( 
.A(n_223),
.B(n_0),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_217),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_251),
.B(n_0),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_214),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_238),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_265),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_179),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_214),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_184),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_197),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_210),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_217),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_217),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_232),
.Y(n_308)
);

OAI21x1_ASAP7_75t_L g309 ( 
.A1(n_201),
.A2(n_82),
.B(n_172),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_217),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_233),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_248),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_214),
.B(n_1),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_230),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_245),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_245),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_254),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_214),
.Y(n_318)
);

OA21x2_ASAP7_75t_L g319 ( 
.A1(n_201),
.A2(n_84),
.B(n_171),
.Y(n_319)
);

XNOR2x1_ASAP7_75t_L g320 ( 
.A(n_190),
.B(n_2),
.Y(n_320)
);

AND2x4_ASAP7_75t_L g321 ( 
.A(n_266),
.B(n_3),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_245),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_245),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_273),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_273),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_199),
.Y(n_326)
);

AOI22x1_ASAP7_75t_SL g327 ( 
.A1(n_219),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_274),
.B(n_4),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_284),
.B(n_7),
.Y(n_329)
);

INVx5_ASAP7_75t_L g330 ( 
.A(n_273),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_286),
.B(n_7),
.Y(n_331)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_182),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_214),
.Y(n_333)
);

OAI21x1_ASAP7_75t_L g334 ( 
.A1(n_205),
.A2(n_88),
.B(n_168),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_205),
.Y(n_335)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_183),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_273),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_187),
.B(n_188),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_189),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_241),
.Y(n_340)
);

AND2x6_ASAP7_75t_L g341 ( 
.A(n_230),
.B(n_35),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_222),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_253),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_222),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_231),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_189),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_247),
.B(n_279),
.Y(n_347)
);

AND2x4_ASAP7_75t_L g348 ( 
.A(n_247),
.B(n_8),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_237),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_237),
.B(n_10),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_178),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_244),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_180),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_189),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_181),
.Y(n_355)
);

BUFx8_ASAP7_75t_SL g356 ( 
.A(n_219),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_244),
.B(n_10),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_185),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_189),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_186),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_235),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_257),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_257),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_279),
.Y(n_364)
);

AND2x6_ASAP7_75t_L g365 ( 
.A(n_277),
.B(n_36),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_277),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_281),
.B(n_12),
.Y(n_367)
);

AND2x4_ASAP7_75t_L g368 ( 
.A(n_281),
.B(n_14),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_191),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_193),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_198),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_294),
.Y(n_372)
);

BUFx10_ASAP7_75t_L g373 ( 
.A(n_295),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_294),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_298),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_298),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_368),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_293),
.B(n_200),
.Y(n_378)
);

AO21x2_ASAP7_75t_L g379 ( 
.A1(n_309),
.A2(n_334),
.B(n_313),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_318),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_318),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_333),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_296),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_348),
.B(n_202),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_333),
.Y(n_385)
);

OAI22xp33_ASAP7_75t_L g386 ( 
.A1(n_328),
.A2(n_288),
.B1(n_280),
.B2(n_290),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_301),
.B(n_304),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_300),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_302),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_332),
.B(n_269),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_305),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_332),
.B(n_283),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_348),
.B(n_369),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_296),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_341),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_364),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_340),
.B(n_287),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_364),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_321),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_305),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_369),
.B(n_371),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_321),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_369),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_369),
.Y(n_404)
);

NAND3xp33_ASAP7_75t_L g405 ( 
.A(n_295),
.B(n_207),
.C(n_203),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_364),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_371),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_336),
.B(n_351),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_341),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_371),
.Y(n_410)
);

NAND2xp33_ASAP7_75t_L g411 ( 
.A(n_341),
.B(n_365),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_296),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_306),
.Y(n_413)
);

OR2x6_ASAP7_75t_L g414 ( 
.A(n_361),
.B(n_208),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_362),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_306),
.Y(n_416)
);

NAND2xp33_ASAP7_75t_L g417 ( 
.A(n_341),
.B(n_291),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_362),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_353),
.B(n_211),
.Y(n_419)
);

NAND3xp33_ASAP7_75t_L g420 ( 
.A(n_297),
.B(n_289),
.C(n_213),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_306),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_363),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_363),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_336),
.B(n_212),
.Y(n_424)
);

NAND3xp33_ASAP7_75t_L g425 ( 
.A(n_343),
.B(n_224),
.C(n_220),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_343),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_314),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_306),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_366),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_307),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_335),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_307),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_335),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_342),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_342),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_344),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_347),
.B(n_234),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_355),
.B(n_239),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_356),
.Y(n_439)
);

BUFx6f_ASAP7_75t_SL g440 ( 
.A(n_370),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_344),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_345),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_345),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_349),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_349),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_352),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_352),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_307),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_303),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_358),
.B(n_243),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_370),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_292),
.A2(n_261),
.B1(n_259),
.B2(n_276),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_360),
.B(n_249),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_310),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g455 ( 
.A(n_308),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_311),
.B(n_192),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_312),
.B(n_250),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_317),
.Y(n_458)
);

INVxp33_ASAP7_75t_L g459 ( 
.A(n_356),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_310),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_310),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_310),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_341),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_315),
.Y(n_464)
);

OR2x2_ASAP7_75t_SL g465 ( 
.A(n_327),
.B(n_256),
.Y(n_465)
);

AND3x2_ASAP7_75t_L g466 ( 
.A(n_350),
.B(n_285),
.C(n_278),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_299),
.B(n_194),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_319),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_357),
.Y(n_469)
);

OR2x6_ASAP7_75t_L g470 ( 
.A(n_329),
.B(n_258),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_367),
.B(n_260),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_331),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_365),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_350),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_338),
.B(n_262),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_330),
.B(n_263),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_315),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_319),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_326),
.B(n_195),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g480 ( 
.A(n_330),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_313),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_330),
.B(n_264),
.Y(n_482)
);

AND2x2_ASAP7_75t_SL g483 ( 
.A(n_319),
.B(n_267),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_320),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_365),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_315),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_472),
.A2(n_229),
.B1(n_240),
.B2(n_365),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_451),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_L g489 ( 
.A1(n_469),
.A2(n_365),
.B1(n_268),
.B2(n_282),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_388),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_427),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_386),
.B(n_14),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_395),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g494 ( 
.A(n_386),
.B(n_391),
.Y(n_494)
);

AND2x6_ASAP7_75t_L g495 ( 
.A(n_395),
.B(n_271),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_373),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_455),
.B(n_196),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_457),
.B(n_204),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_457),
.B(n_206),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_400),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_390),
.B(n_221),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_409),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_426),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_423),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_373),
.Y(n_505)
);

INVxp67_ASAP7_75t_SL g506 ( 
.A(n_463),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_439),
.Y(n_507)
);

NAND2xp33_ASAP7_75t_L g508 ( 
.A(n_481),
.B(n_209),
.Y(n_508)
);

NAND2xp33_ASAP7_75t_L g509 ( 
.A(n_485),
.B(n_215),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_408),
.B(n_437),
.Y(n_510)
);

NOR2xp67_ASAP7_75t_SL g511 ( 
.A(n_463),
.B(n_216),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_475),
.B(n_218),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_446),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_415),
.Y(n_514)
);

BUFx6f_ASAP7_75t_SL g515 ( 
.A(n_414),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_475),
.B(n_227),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_405),
.B(n_399),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_449),
.B(n_228),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_404),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_397),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_392),
.B(n_226),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_470),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_470),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_473),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_458),
.B(n_242),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_440),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_474),
.B(n_402),
.Y(n_527)
);

INVx2_ASAP7_75t_SL g528 ( 
.A(n_377),
.Y(n_528)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_440),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_425),
.B(n_246),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_418),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_420),
.B(n_252),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_384),
.B(n_236),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_384),
.B(n_255),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_378),
.B(n_424),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_456),
.B(n_424),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_SL g537 ( 
.A(n_473),
.B(n_270),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_479),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_438),
.A2(n_359),
.B1(n_354),
.B2(n_346),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_471),
.B(n_272),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_467),
.B(n_275),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_422),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_429),
.B(n_15),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_466),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_438),
.B(n_278),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_393),
.B(n_330),
.Y(n_546)
);

NOR2x2_ASAP7_75t_L g547 ( 
.A(n_414),
.B(n_15),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_431),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_433),
.Y(n_549)
);

OAI21xp33_ASAP7_75t_L g550 ( 
.A1(n_419),
.A2(n_359),
.B(n_354),
.Y(n_550)
);

AND2x6_ASAP7_75t_SL g551 ( 
.A(n_414),
.B(n_18),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_434),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_419),
.B(n_339),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_396),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_450),
.B(n_339),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_435),
.B(n_18),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_387),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_453),
.B(n_346),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_372),
.B(n_346),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_466),
.B(n_379),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_372),
.B(n_374),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_436),
.B(n_441),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_442),
.B(n_443),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_444),
.B(n_354),
.Y(n_564)
);

INVxp67_ASAP7_75t_SL g565 ( 
.A(n_374),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_445),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_447),
.Y(n_567)
);

AO22x2_ASAP7_75t_L g568 ( 
.A1(n_484),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_375),
.A2(n_359),
.B1(n_337),
.B2(n_325),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_398),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_376),
.B(n_359),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_406),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_459),
.B(n_21),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_482),
.Y(n_574)
);

INVx5_ASAP7_75t_L g575 ( 
.A(n_480),
.Y(n_575)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_465),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_406),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_376),
.B(n_316),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_403),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_389),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_536),
.A2(n_411),
.B(n_417),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_528),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_535),
.B(n_483),
.Y(n_583)
);

AOI21xp5_ASAP7_75t_L g584 ( 
.A1(n_535),
.A2(n_468),
.B(n_478),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_494),
.A2(n_483),
.B1(n_468),
.B2(n_478),
.Y(n_585)
);

O2A1O1Ixp5_ASAP7_75t_L g586 ( 
.A1(n_512),
.A2(n_476),
.B(n_482),
.C(n_401),
.Y(n_586)
);

OAI21xp33_ASAP7_75t_L g587 ( 
.A1(n_527),
.A2(n_389),
.B(n_380),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_510),
.B(n_379),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_522),
.B(n_380),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_537),
.B(n_381),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_580),
.Y(n_591)
);

XOR2xp5_ASAP7_75t_L g592 ( 
.A(n_507),
.B(n_459),
.Y(n_592)
);

NOR3xp33_ASAP7_75t_L g593 ( 
.A(n_520),
.B(n_382),
.C(n_385),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_SL g594 ( 
.A(n_515),
.B(n_382),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_523),
.B(n_496),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_567),
.B(n_385),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_490),
.B(n_407),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g598 ( 
.A1(n_517),
.A2(n_410),
.B(n_486),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_537),
.B(n_316),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_503),
.Y(n_600)
);

OAI21x1_ASAP7_75t_L g601 ( 
.A1(n_561),
.A2(n_432),
.B(n_477),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_566),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_500),
.B(n_22),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_493),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_L g605 ( 
.A1(n_487),
.A2(n_488),
.B1(n_563),
.B2(n_562),
.Y(n_605)
);

NAND2x1p5_ASAP7_75t_L g606 ( 
.A(n_505),
.B(n_23),
.Y(n_606)
);

BUFx4f_ASAP7_75t_L g607 ( 
.A(n_492),
.Y(n_607)
);

NAND2x1p5_ASAP7_75t_L g608 ( 
.A(n_538),
.B(n_25),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_543),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_565),
.A2(n_416),
.B(n_464),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_SL g611 ( 
.A1(n_515),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_498),
.B(n_499),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_556),
.Y(n_613)
);

OAI21x1_ASAP7_75t_L g614 ( 
.A1(n_553),
.A2(n_462),
.B(n_461),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_498),
.B(n_29),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_506),
.A2(n_460),
.B(n_454),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_514),
.Y(n_617)
);

AOI21x1_ASAP7_75t_L g618 ( 
.A1(n_560),
.A2(n_454),
.B(n_448),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_574),
.A2(n_432),
.B(n_430),
.Y(n_619)
);

CKINVDCx10_ASAP7_75t_R g620 ( 
.A(n_557),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_499),
.B(n_31),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_518),
.A2(n_430),
.B(n_428),
.Y(n_622)
);

A2O1A1Ixp33_ASAP7_75t_L g623 ( 
.A1(n_545),
.A2(n_322),
.B(n_325),
.C(n_337),
.Y(n_623)
);

A2O1A1Ixp33_ASAP7_75t_L g624 ( 
.A1(n_548),
.A2(n_322),
.B(n_325),
.C(n_337),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_525),
.A2(n_412),
.B(n_416),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_502),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_524),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_540),
.A2(n_413),
.B(n_412),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_526),
.B(n_32),
.Y(n_629)
);

OAI21x1_ASAP7_75t_L g630 ( 
.A1(n_553),
.A2(n_413),
.B(n_421),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_540),
.A2(n_421),
.B(n_394),
.Y(n_631)
);

O2A1O1Ixp5_ASAP7_75t_L g632 ( 
.A1(n_516),
.A2(n_532),
.B(n_501),
.C(n_521),
.Y(n_632)
);

A2O1A1Ixp33_ASAP7_75t_L g633 ( 
.A1(n_549),
.A2(n_324),
.B(n_323),
.C(n_383),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_560),
.B(n_497),
.Y(n_634)
);

A2O1A1Ixp33_ASAP7_75t_L g635 ( 
.A1(n_552),
.A2(n_324),
.B(n_323),
.C(n_383),
.Y(n_635)
);

BUFx12f_ASAP7_75t_L g636 ( 
.A(n_551),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_533),
.B(n_41),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_575),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_508),
.A2(n_43),
.B(n_59),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_491),
.Y(n_640)
);

A2O1A1Ixp33_ASAP7_75t_L g641 ( 
.A1(n_531),
.A2(n_64),
.B(n_65),
.C(n_69),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_542),
.Y(n_642)
);

AO21x1_ASAP7_75t_L g643 ( 
.A1(n_555),
.A2(n_71),
.B(n_76),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_529),
.B(n_175),
.Y(n_644)
);

O2A1O1Ixp33_ASAP7_75t_L g645 ( 
.A1(n_530),
.A2(n_573),
.B(n_541),
.C(n_513),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_576),
.B(n_79),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_534),
.B(n_167),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_504),
.B(n_495),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_L g649 ( 
.A1(n_489),
.A2(n_92),
.B(n_93),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_L g650 ( 
.A1(n_558),
.A2(n_97),
.B(n_100),
.Y(n_650)
);

OAI21xp5_ASAP7_75t_L g651 ( 
.A1(n_578),
.A2(n_103),
.B(n_105),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_546),
.A2(n_106),
.B(n_107),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_495),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_559),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_568),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_578),
.A2(n_111),
.B(n_112),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_568),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_575),
.B(n_114),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_588),
.A2(n_509),
.B(n_571),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_612),
.B(n_575),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_583),
.A2(n_579),
.B(n_577),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_581),
.A2(n_554),
.B(n_572),
.Y(n_662)
);

OAI21xp5_ASAP7_75t_L g663 ( 
.A1(n_585),
.A2(n_564),
.B(n_570),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_600),
.B(n_575),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_617),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_592),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_642),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_654),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_631),
.A2(n_519),
.B(n_550),
.Y(n_669)
);

INVx5_ASAP7_75t_L g670 ( 
.A(n_653),
.Y(n_670)
);

O2A1O1Ixp33_ASAP7_75t_L g671 ( 
.A1(n_605),
.A2(n_539),
.B(n_547),
.C(n_569),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_L g672 ( 
.A1(n_632),
.A2(n_511),
.B(n_117),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_586),
.A2(n_116),
.B(n_118),
.Y(n_673)
);

AO31x2_ASAP7_75t_L g674 ( 
.A1(n_643),
.A2(n_125),
.A3(n_129),
.B(n_132),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_613),
.B(n_134),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_609),
.B(n_135),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_604),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_608),
.B(n_147),
.Y(n_678)
);

OAI21x1_ASAP7_75t_L g679 ( 
.A1(n_618),
.A2(n_151),
.B(n_152),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_607),
.B(n_595),
.Y(n_680)
);

NAND3xp33_ASAP7_75t_L g681 ( 
.A(n_603),
.B(n_157),
.C(n_159),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_591),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_619),
.A2(n_162),
.B(n_163),
.Y(n_683)
);

AOI221x1_ASAP7_75t_L g684 ( 
.A1(n_623),
.A2(n_164),
.B1(n_651),
.B2(n_650),
.C(n_649),
.Y(n_684)
);

BUFx12f_ASAP7_75t_L g685 ( 
.A(n_636),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_602),
.B(n_593),
.Y(n_686)
);

AOI21xp5_ASAP7_75t_L g687 ( 
.A1(n_610),
.A2(n_616),
.B(n_628),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_595),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_606),
.B(n_589),
.Y(n_689)
);

OR2x6_ASAP7_75t_L g690 ( 
.A(n_644),
.B(n_653),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_597),
.A2(n_645),
.B(n_637),
.Y(n_691)
);

AO31x2_ASAP7_75t_L g692 ( 
.A1(n_641),
.A2(n_624),
.A3(n_635),
.B(n_633),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_620),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_582),
.B(n_589),
.Y(n_694)
);

INVx5_ASAP7_75t_L g695 ( 
.A(n_591),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_638),
.B(n_644),
.Y(n_696)
);

NAND3x1_ASAP7_75t_L g697 ( 
.A(n_655),
.B(n_646),
.C(n_629),
.Y(n_697)
);

OAI21xp5_ASAP7_75t_L g698 ( 
.A1(n_587),
.A2(n_596),
.B(n_647),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_615),
.B(n_621),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_622),
.A2(n_625),
.B(n_598),
.Y(n_700)
);

AO31x2_ASAP7_75t_L g701 ( 
.A1(n_639),
.A2(n_656),
.A3(n_658),
.B(n_652),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_640),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_594),
.A2(n_611),
.B1(n_648),
.B2(n_638),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_604),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_626),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_626),
.B(n_627),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_627),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_588),
.A2(n_583),
.B(n_584),
.Y(n_708)
);

NOR2xp67_ASAP7_75t_L g709 ( 
.A(n_638),
.B(n_591),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_617),
.Y(n_710)
);

OAI21xp5_ASAP7_75t_L g711 ( 
.A1(n_584),
.A2(n_588),
.B(n_581),
.Y(n_711)
);

AOI21xp33_ASAP7_75t_L g712 ( 
.A1(n_612),
.A2(n_494),
.B(n_544),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_612),
.B(n_472),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_612),
.B(n_472),
.Y(n_714)
);

BUFx2_ASAP7_75t_L g715 ( 
.A(n_600),
.Y(n_715)
);

OAI21x1_ASAP7_75t_L g716 ( 
.A1(n_614),
.A2(n_601),
.B(n_630),
.Y(n_716)
);

OAI21xp5_ASAP7_75t_SL g717 ( 
.A1(n_608),
.A2(n_452),
.B(n_492),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_612),
.B(n_472),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_607),
.B(n_484),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_612),
.B(n_472),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_607),
.A2(n_304),
.B1(n_326),
.B2(n_301),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_588),
.A2(n_583),
.B(n_584),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_620),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_L g724 ( 
.A1(n_583),
.A2(n_607),
.B1(n_609),
.B2(n_596),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_617),
.Y(n_725)
);

AO31x2_ASAP7_75t_L g726 ( 
.A1(n_585),
.A2(n_643),
.A3(n_588),
.B(n_623),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_588),
.A2(n_583),
.B(n_584),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_612),
.B(n_472),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_583),
.A2(n_607),
.B1(n_609),
.B2(n_596),
.Y(n_729)
);

INVx5_ASAP7_75t_L g730 ( 
.A(n_653),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_588),
.A2(n_583),
.B(n_584),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_612),
.B(n_472),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_612),
.B(n_472),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_607),
.B(n_484),
.Y(n_734)
);

BUFx2_ASAP7_75t_SL g735 ( 
.A(n_600),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_612),
.B(n_472),
.Y(n_736)
);

CKINVDCx14_ASAP7_75t_R g737 ( 
.A(n_592),
.Y(n_737)
);

AO31x2_ASAP7_75t_L g738 ( 
.A1(n_585),
.A2(n_643),
.A3(n_588),
.B(n_623),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_612),
.B(n_472),
.Y(n_739)
);

O2A1O1Ixp5_ASAP7_75t_L g740 ( 
.A1(n_599),
.A2(n_590),
.B(n_632),
.C(n_634),
.Y(n_740)
);

OAI21x1_ASAP7_75t_L g741 ( 
.A1(n_614),
.A2(n_601),
.B(n_630),
.Y(n_741)
);

AOI21xp33_ASAP7_75t_L g742 ( 
.A1(n_697),
.A2(n_699),
.B(n_671),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_690),
.A2(n_724),
.B1(n_729),
.B2(n_739),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_717),
.A2(n_712),
.B1(n_732),
.B2(n_713),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_693),
.Y(n_745)
);

AO21x2_ASAP7_75t_L g746 ( 
.A1(n_731),
.A2(n_672),
.B(n_673),
.Y(n_746)
);

NAND2x1p5_ASAP7_75t_L g747 ( 
.A(n_670),
.B(n_730),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_710),
.Y(n_748)
);

O2A1O1Ixp33_ASAP7_75t_L g749 ( 
.A1(n_714),
.A2(n_720),
.B(n_736),
.C(n_728),
.Y(n_749)
);

BUFx12f_ASAP7_75t_L g750 ( 
.A(n_723),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_685),
.Y(n_751)
);

CKINVDCx11_ASAP7_75t_R g752 ( 
.A(n_666),
.Y(n_752)
);

OAI221xp5_ASAP7_75t_L g753 ( 
.A1(n_718),
.A2(n_733),
.B1(n_734),
.B2(n_719),
.C(n_721),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_725),
.B(n_665),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_680),
.A2(n_735),
.B1(n_688),
.B2(n_689),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_667),
.B(n_725),
.Y(n_756)
);

INVx1_ASAP7_75t_SL g757 ( 
.A(n_704),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_L g758 ( 
.A1(n_690),
.A2(n_660),
.B1(n_696),
.B2(n_703),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_668),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_694),
.B(n_696),
.Y(n_760)
);

AO31x2_ASAP7_75t_L g761 ( 
.A1(n_684),
.A2(n_700),
.A3(n_687),
.B(n_691),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_686),
.B(n_702),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_702),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_698),
.A2(n_669),
.B(n_662),
.Y(n_764)
);

NOR2x1_ASAP7_75t_R g765 ( 
.A(n_730),
.B(n_695),
.Y(n_765)
);

OR2x6_ASAP7_75t_L g766 ( 
.A(n_678),
.B(n_664),
.Y(n_766)
);

AND2x6_ASAP7_75t_L g767 ( 
.A(n_677),
.B(n_706),
.Y(n_767)
);

OAI21xp5_ASAP7_75t_L g768 ( 
.A1(n_661),
.A2(n_659),
.B(n_740),
.Y(n_768)
);

BUFx12f_ASAP7_75t_L g769 ( 
.A(n_695),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_695),
.B(n_682),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_682),
.B(n_737),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_709),
.B(n_675),
.Y(n_772)
);

AO21x1_ASAP7_75t_L g773 ( 
.A1(n_683),
.A2(n_663),
.B(n_679),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_709),
.A2(n_676),
.B1(n_681),
.B2(n_705),
.Y(n_774)
);

INVx8_ASAP7_75t_L g775 ( 
.A(n_707),
.Y(n_775)
);

A2O1A1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_726),
.A2(n_738),
.B(n_674),
.C(n_701),
.Y(n_776)
);

OAI21x1_ASAP7_75t_L g777 ( 
.A1(n_726),
.A2(n_738),
.B(n_701),
.Y(n_777)
);

INVx1_ASAP7_75t_SL g778 ( 
.A(n_692),
.Y(n_778)
);

OR2x6_ASAP7_75t_SL g779 ( 
.A(n_692),
.B(n_701),
.Y(n_779)
);

OAI21xp5_ASAP7_75t_L g780 ( 
.A1(n_708),
.A2(n_727),
.B(n_722),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_717),
.B(n_484),
.Y(n_781)
);

INVx1_ASAP7_75t_SL g782 ( 
.A(n_735),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_717),
.A2(n_657),
.B1(n_607),
.B2(n_605),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_712),
.A2(n_607),
.B1(n_657),
.B2(n_414),
.Y(n_784)
);

NAND4xp25_ASAP7_75t_L g785 ( 
.A(n_717),
.B(n_492),
.C(n_712),
.D(n_494),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_715),
.Y(n_786)
);

CKINVDCx6p67_ASAP7_75t_R g787 ( 
.A(n_685),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_690),
.A2(n_607),
.B1(n_583),
.B2(n_724),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_710),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_710),
.Y(n_790)
);

OR2x6_ASAP7_75t_L g791 ( 
.A(n_690),
.B(n_735),
.Y(n_791)
);

OA21x2_ASAP7_75t_L g792 ( 
.A1(n_711),
.A2(n_741),
.B(n_716),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_712),
.A2(n_607),
.B1(n_657),
.B2(n_414),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_693),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_748),
.Y(n_795)
);

AOI221xp5_ASAP7_75t_L g796 ( 
.A1(n_785),
.A2(n_753),
.B1(n_781),
.B2(n_749),
.C(n_742),
.Y(n_796)
);

BUFx2_ASAP7_75t_L g797 ( 
.A(n_767),
.Y(n_797)
);

OA21x2_ASAP7_75t_L g798 ( 
.A1(n_776),
.A2(n_780),
.B(n_764),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_744),
.B(n_756),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_782),
.B(n_744),
.Y(n_800)
);

CKINVDCx11_ASAP7_75t_R g801 ( 
.A(n_787),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_763),
.B(n_759),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_789),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_769),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_786),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_790),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_754),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_762),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_792),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_782),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_775),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_785),
.A2(n_783),
.B1(n_743),
.B2(n_788),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_783),
.A2(n_784),
.B1(n_793),
.B2(n_758),
.Y(n_813)
);

INVx1_ASAP7_75t_SL g814 ( 
.A(n_757),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_775),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_747),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_778),
.Y(n_817)
);

BUFx2_ASAP7_75t_L g818 ( 
.A(n_767),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_775),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_760),
.B(n_779),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_766),
.B(n_778),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_755),
.B(n_757),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_777),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_791),
.Y(n_824)
);

HB1xp67_ASAP7_75t_L g825 ( 
.A(n_791),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_761),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_768),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_L g828 ( 
.A1(n_812),
.A2(n_791),
.B1(n_774),
.B2(n_772),
.Y(n_828)
);

INVx4_ASAP7_75t_L g829 ( 
.A(n_797),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_795),
.Y(n_830)
);

OR2x2_ASAP7_75t_L g831 ( 
.A(n_799),
.B(n_770),
.Y(n_831)
);

INVxp67_ASAP7_75t_L g832 ( 
.A(n_810),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_820),
.B(n_746),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_809),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_820),
.B(n_746),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_805),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_808),
.B(n_771),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_803),
.B(n_806),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_803),
.B(n_806),
.Y(n_839)
);

INVxp67_ASAP7_75t_SL g840 ( 
.A(n_807),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_802),
.B(n_773),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_833),
.B(n_827),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_834),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_833),
.B(n_827),
.Y(n_844)
);

AND2x2_ASAP7_75t_SL g845 ( 
.A(n_829),
.B(n_818),
.Y(n_845)
);

OR2x2_ASAP7_75t_L g846 ( 
.A(n_835),
.B(n_821),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_841),
.B(n_817),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_838),
.B(n_796),
.Y(n_848)
);

OR2x2_ASAP7_75t_L g849 ( 
.A(n_831),
.B(n_821),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_830),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_841),
.B(n_823),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_836),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_839),
.B(n_826),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_842),
.B(n_844),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_850),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_843),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_842),
.B(n_844),
.Y(n_857)
);

HB1xp67_ASAP7_75t_L g858 ( 
.A(n_852),
.Y(n_858)
);

NOR2x1_ASAP7_75t_SL g859 ( 
.A(n_845),
.B(n_829),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_851),
.B(n_798),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_845),
.B(n_829),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_848),
.B(n_840),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_853),
.B(n_832),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_847),
.B(n_798),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_854),
.B(n_846),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_858),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_855),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_861),
.B(n_845),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_856),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_854),
.B(n_847),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_856),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_857),
.B(n_846),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_862),
.B(n_814),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_871),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_869),
.Y(n_875)
);

AOI21xp33_ASAP7_75t_SL g876 ( 
.A1(n_868),
.A2(n_745),
.B(n_794),
.Y(n_876)
);

INVx3_ASAP7_75t_L g877 ( 
.A(n_869),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_865),
.B(n_857),
.Y(n_878)
);

INVxp67_ASAP7_75t_SL g879 ( 
.A(n_866),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_872),
.B(n_860),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_871),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_866),
.B(n_860),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_867),
.Y(n_883)
);

O2A1O1Ixp33_ASAP7_75t_SL g884 ( 
.A1(n_868),
.A2(n_863),
.B(n_859),
.C(n_751),
.Y(n_884)
);

INVx1_ASAP7_75t_SL g885 ( 
.A(n_870),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_882),
.B(n_864),
.Y(n_886)
);

INVx1_ASAP7_75t_SL g887 ( 
.A(n_877),
.Y(n_887)
);

AOI21xp33_ASAP7_75t_L g888 ( 
.A1(n_876),
.A2(n_873),
.B(n_837),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_883),
.Y(n_889)
);

OR2x2_ASAP7_75t_L g890 ( 
.A(n_885),
.B(n_864),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_876),
.A2(n_873),
.B1(n_829),
.B2(n_849),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_889),
.B(n_879),
.Y(n_892)
);

NAND4xp25_ASAP7_75t_L g893 ( 
.A(n_891),
.B(n_884),
.C(n_813),
.D(n_804),
.Y(n_893)
);

NAND4xp25_ASAP7_75t_L g894 ( 
.A(n_888),
.B(n_804),
.C(n_828),
.D(n_822),
.Y(n_894)
);

NOR2x1_ASAP7_75t_L g895 ( 
.A(n_893),
.B(n_801),
.Y(n_895)
);

NOR3x1_ASAP7_75t_L g896 ( 
.A(n_894),
.B(n_890),
.C(n_824),
.Y(n_896)
);

NOR2x1_ASAP7_75t_L g897 ( 
.A(n_895),
.B(n_887),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_896),
.B(n_892),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_898),
.B(n_883),
.Y(n_899)
);

INVxp67_ASAP7_75t_L g900 ( 
.A(n_897),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_899),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_900),
.B(n_750),
.Y(n_902)
);

NOR4xp25_ASAP7_75t_L g903 ( 
.A(n_901),
.B(n_752),
.C(n_881),
.D(n_874),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_902),
.A2(n_800),
.B(n_881),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_902),
.Y(n_905)
);

XOR2x2_ASAP7_75t_L g906 ( 
.A(n_904),
.B(n_825),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_905),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_903),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_905),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_SL g910 ( 
.A1(n_905),
.A2(n_824),
.B1(n_815),
.B2(n_811),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_907),
.A2(n_877),
.B1(n_875),
.B2(n_886),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_909),
.B(n_877),
.Y(n_912)
);

OAI22x1_ASAP7_75t_L g913 ( 
.A1(n_908),
.A2(n_906),
.B1(n_910),
.B2(n_816),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_907),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_907),
.A2(n_765),
.B(n_874),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_907),
.Y(n_916)
);

AOI22xp33_ASAP7_75t_L g917 ( 
.A1(n_916),
.A2(n_875),
.B1(n_880),
.B2(n_878),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_914),
.A2(n_880),
.B1(n_878),
.B2(n_828),
.Y(n_918)
);

INVx2_ASAP7_75t_SL g919 ( 
.A(n_912),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_919),
.Y(n_920)
);

AO221x2_ASAP7_75t_L g921 ( 
.A1(n_920),
.A2(n_913),
.B1(n_911),
.B2(n_915),
.C(n_918),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_921),
.A2(n_917),
.B(n_765),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_922),
.A2(n_815),
.B(n_819),
.Y(n_923)
);


endmodule