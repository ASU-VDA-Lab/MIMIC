module fake_ariane_2924_n_132 (n_8, n_7, n_22, n_1, n_6, n_13, n_20, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_132);

input n_8;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;

output n_132;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_119;
wire n_124;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_120;
wire n_106;
wire n_53;
wire n_111;
wire n_115;
wire n_66;
wire n_71;
wire n_24;
wire n_109;
wire n_96;
wire n_49;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_30;
wire n_82;
wire n_42;
wire n_31;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_85;
wire n_130;
wire n_94;
wire n_101;
wire n_48;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_112;
wire n_45;
wire n_129;
wire n_126;
wire n_122;
wire n_52;
wire n_73;
wire n_77;
wire n_118;
wire n_93;
wire n_121;
wire n_61;
wire n_108;
wire n_102;
wire n_125;
wire n_43;
wire n_87;
wire n_81;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_116;
wire n_104;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_127;
wire n_35;
wire n_54;
wire n_25;

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_23),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_19),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_22),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_1),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

NAND3xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_1),
.C(n_2),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_28),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_3),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_30),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_36),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_26),
.Y(n_58)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_32),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_38),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

OAI21x1_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_46),
.B(n_47),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_42),
.B(n_45),
.C(n_49),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_43),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_52),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_51),
.B(n_46),
.C(n_50),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_53),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_53),
.B(n_50),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

AOI21x1_ASAP7_75t_SL g76 ( 
.A1(n_69),
.A2(n_60),
.B(n_59),
.Y(n_76)
);

CKINVDCx5p33_ASAP7_75t_R g77 ( 
.A(n_67),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_35),
.B1(n_29),
.B2(n_44),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_65),
.A2(n_56),
.B(n_63),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_39),
.B1(n_40),
.B2(n_31),
.Y(n_80)
);

AOI221x1_ASAP7_75t_SL g81 ( 
.A1(n_68),
.A2(n_52),
.B1(n_49),
.B2(n_33),
.C(n_9),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_59),
.B(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_55),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_63),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_50),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_50),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_56),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_86),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_78),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_81),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_96),
.A2(n_78),
.B1(n_88),
.B2(n_97),
.Y(n_105)
);

OR2x6_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_98),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_88),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_105),
.A2(n_97),
.B1(n_96),
.B2(n_91),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_90),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_105),
.A2(n_104),
.B(n_91),
.C(n_103),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_90),
.B1(n_48),
.B2(n_56),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_48),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_64),
.B(n_82),
.C(n_53),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

AOI211x1_ASAP7_75t_L g116 ( 
.A1(n_110),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_116)
);

NAND4xp25_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_79),
.C(n_9),
.D(n_60),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_107),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_112),
.B(n_53),
.Y(n_119)
);

NAND4xp25_ASAP7_75t_SL g120 ( 
.A(n_111),
.B(n_11),
.C(n_12),
.D(n_16),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_120),
.B(n_106),
.Y(n_121)
);

NAND2x1_ASAP7_75t_SL g122 ( 
.A(n_115),
.B(n_114),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_123),
.Y(n_124)
);

AND2x4_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_119),
.Y(n_125)
);

NOR3xp33_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_117),
.C(n_116),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_64),
.Y(n_127)
);

XNOR2x1_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_125),
.Y(n_128)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_125),
.B1(n_121),
.B2(n_122),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_129),
.A2(n_122),
.B1(n_48),
.B2(n_21),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_128),
.Y(n_131)
);

AOI31xp33_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_76),
.A3(n_48),
.B(n_20),
.Y(n_132)
);


endmodule