module fake_jpeg_17745_n_172 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_172);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_4),
.B(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx6p67_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_14),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_39),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_0),
.C(n_4),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_36),
.B(n_52),
.Y(n_83)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_0),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_22),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_40),
.A2(n_42),
.B1(n_43),
.B2(n_50),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_22),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_14),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_30),
.B(n_10),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

CKINVDCx12_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_28),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_48),
.Y(n_66)
);

INVx5_ASAP7_75t_SL g48 ( 
.A(n_28),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_55),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_26),
.A2(n_31),
.B1(n_29),
.B2(n_33),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_23),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_57),
.Y(n_69)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_32),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_58),
.B(n_63),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_32),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_32),
.Y(n_72)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_36),
.B(n_31),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_78),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_41),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_75),
.B(n_81),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_29),
.B1(n_26),
.B2(n_23),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_77),
.A2(n_82),
.B(n_53),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_19),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_19),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_80),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_41),
.B(n_21),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_20),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_48),
.A2(n_21),
.B1(n_25),
.B2(n_27),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_34),
.B(n_18),
.Y(n_84)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_74),
.A2(n_25),
.B1(n_27),
.B2(n_34),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_61),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_SL g123 ( 
.A(n_88),
.B(n_91),
.C(n_100),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_72),
.A2(n_34),
.B(n_41),
.C(n_53),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_83),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_97),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_59),
.A2(n_79),
.B1(n_78),
.B2(n_70),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_96),
.A2(n_106),
.B1(n_108),
.B2(n_86),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_58),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_68),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_94),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_68),
.A2(n_69),
.B(n_67),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_71),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_105),
.B(n_110),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_59),
.A2(n_67),
.B1(n_84),
.B2(n_80),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_64),
.A2(n_60),
.B1(n_71),
.B2(n_66),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_64),
.A2(n_60),
.B1(n_65),
.B2(n_75),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_109),
.A2(n_61),
.B1(n_76),
.B2(n_104),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_76),
.Y(n_110)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_113),
.A2(n_119),
.B1(n_129),
.B2(n_130),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_76),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_116),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_76),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_102),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_121),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_103),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_90),
.C(n_97),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_132),
.C(n_126),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_131),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_92),
.B(n_101),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_127),
.Y(n_143)
);

BUFx24_ASAP7_75t_SL g128 ( 
.A(n_92),
.Y(n_128)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_90),
.A2(n_93),
.B1(n_109),
.B2(n_88),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_101),
.B(n_93),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_100),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_91),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_98),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_135),
.B(n_138),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_89),
.B(n_110),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_89),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_147),
.Y(n_156)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_113),
.C(n_117),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_124),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_123),
.B1(n_122),
.B2(n_133),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_146),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_118),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_118),
.C(n_135),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_154),
.Y(n_160)
);

BUFx12_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_157),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_156),
.A2(n_148),
.B1(n_136),
.B2(n_145),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_162),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_150),
.B(n_143),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_153),
.C(n_155),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_151),
.C(n_158),
.Y(n_165)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_155),
.C(n_149),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_165),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_161),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_167),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_160),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_137),
.B1(n_168),
.B2(n_169),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);


endmodule