module fake_jpeg_22030_n_338 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_19;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_42),
.Y(n_61)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_22),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_48),
.Y(n_72)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_24),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_60),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_50),
.Y(n_78)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_53),
.Y(n_86)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_21),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_58),
.B(n_63),
.Y(n_93)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_30),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_64),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_18),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_32),
.B(n_28),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_31),
.Y(n_82)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_70),
.Y(n_98)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_71),
.B(n_73),
.Y(n_114)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_15),
.B1(n_16),
.B2(n_24),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_74),
.A2(n_92),
.B1(n_70),
.B2(n_71),
.Y(n_109)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_79),
.Y(n_119)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_81),
.A2(n_84),
.B1(n_87),
.B2(n_88),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_82),
.B(n_50),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_47),
.A2(n_15),
.B1(n_16),
.B2(n_28),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_67),
.A2(n_15),
.B1(n_16),
.B2(n_28),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_65),
.A2(n_15),
.B1(n_16),
.B2(n_24),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_90),
.A2(n_63),
.B1(n_58),
.B2(n_43),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_95),
.A2(n_105),
.B1(n_106),
.B2(n_117),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_36),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_102),
.Y(n_125)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_101),
.Y(n_122)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_78),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_118),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_L g104 ( 
.A1(n_68),
.A2(n_55),
.B1(n_38),
.B2(n_24),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_104),
.A2(n_26),
.B1(n_91),
.B2(n_57),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_89),
.A2(n_49),
.B1(n_46),
.B2(n_59),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_49),
.B1(n_46),
.B2(n_59),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_68),
.A2(n_61),
.B(n_64),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_107),
.A2(n_51),
.B(n_21),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_90),
.A2(n_34),
.B1(n_60),
.B2(n_44),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_109),
.B1(n_112),
.B2(n_79),
.Y(n_127)
);

FAx1_ASAP7_75t_SL g110 ( 
.A(n_77),
.B(n_42),
.CI(n_66),
.CON(n_110),
.SN(n_110)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_110),
.B(n_115),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_77),
.B(n_42),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_116),
.C(n_21),
.Y(n_124)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_93),
.B(n_42),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_17),
.B1(n_31),
.B2(n_53),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_69),
.B(n_48),
.Y(n_118)
);

OAI22x1_ASAP7_75t_SL g121 ( 
.A1(n_94),
.A2(n_83),
.B1(n_55),
.B2(n_73),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_121),
.A2(n_127),
.B1(n_147),
.B2(n_106),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_124),
.A2(n_135),
.B(n_145),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_103),
.B(n_80),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_129),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_32),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_131),
.Y(n_153)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_135),
.B(n_125),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_107),
.A2(n_18),
.B(n_87),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_138),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_99),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_137),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_119),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_94),
.A2(n_17),
.B(n_31),
.C(n_55),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_139),
.A2(n_116),
.B(n_113),
.Y(n_152)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_142),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

OAI32xp33_ASAP7_75t_L g143 ( 
.A1(n_108),
.A2(n_18),
.A3(n_37),
.B1(n_39),
.B2(n_31),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_113),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_109),
.A2(n_75),
.B1(n_81),
.B2(n_26),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_144),
.A2(n_146),
.B1(n_112),
.B2(n_117),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_113),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_95),
.A2(n_39),
.B1(n_37),
.B2(n_17),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_148),
.B(n_156),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_145),
.A2(n_110),
.B(n_116),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_151),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g177 ( 
.A1(n_152),
.A2(n_151),
.B1(n_163),
.B2(n_159),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_154),
.A2(n_166),
.B1(n_146),
.B2(n_121),
.Y(n_178)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_160),
.Y(n_174)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_157),
.B(n_159),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_158),
.A2(n_97),
.B1(n_111),
.B2(n_57),
.Y(n_197)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_171),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_140),
.B(n_110),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_141),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_110),
.B(n_96),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_163),
.A2(n_139),
.B1(n_141),
.B2(n_100),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_125),
.A2(n_123),
.B(n_134),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_123),
.C(n_145),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_121),
.A2(n_112),
.B1(n_111),
.B2(n_101),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_170),
.A2(n_144),
.B1(n_147),
.B2(n_139),
.Y(n_181)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_127),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_99),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_124),
.B(n_96),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_173),
.B(n_136),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_175),
.B(n_195),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_177),
.A2(n_178),
.B(n_188),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_180),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_181),
.A2(n_190),
.B1(n_192),
.B2(n_198),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_133),
.C(n_130),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_150),
.C(n_180),
.Y(n_217)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_186),
.Y(n_211)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_153),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_131),
.Y(n_187)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_187),
.Y(n_214)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_158),
.A2(n_138),
.B1(n_139),
.B2(n_143),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_191),
.B(n_17),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_172),
.A2(n_139),
.B1(n_115),
.B2(n_111),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

OAI32xp33_ASAP7_75t_L g195 ( 
.A1(n_161),
.A2(n_139),
.A3(n_97),
.B1(n_17),
.B2(n_31),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_26),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_196),
.A2(n_156),
.B(n_148),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_197),
.B(n_169),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_170),
.A2(n_99),
.B1(n_120),
.B2(n_27),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_164),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_199),
.A2(n_157),
.B1(n_167),
.B2(n_149),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_201),
.A2(n_205),
.B(n_208),
.Y(n_232)
);

INVxp33_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_203),
.A2(n_218),
.B1(n_219),
.B2(n_223),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_168),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_177),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_200),
.A2(n_168),
.B(n_162),
.Y(n_205)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_207),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_189),
.A2(n_152),
.B(n_149),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_190),
.A2(n_154),
.B1(n_166),
.B2(n_171),
.Y(n_210)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_210),
.Y(n_242)
);

OA21x2_ASAP7_75t_L g212 ( 
.A1(n_197),
.A2(n_152),
.B(n_169),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_212),
.A2(n_29),
.B(n_27),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_189),
.A2(n_167),
.B(n_173),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_215),
.A2(n_196),
.B(n_30),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_174),
.Y(n_216)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_216),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_177),
.C(n_193),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_187),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_181),
.A2(n_198),
.B1(n_183),
.B2(n_179),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_220),
.A2(n_226),
.B1(n_184),
.B2(n_186),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_224),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_178),
.A2(n_120),
.B1(n_30),
.B2(n_29),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_227),
.A2(n_229),
.B1(n_231),
.B2(n_237),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_176),
.Y(n_228)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_228),
.Y(n_254)
);

HAxp5_ASAP7_75t_SL g229 ( 
.A(n_214),
.B(n_199),
.CON(n_229),
.SN(n_229)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_202),
.C(n_205),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_223),
.A2(n_188),
.B1(n_195),
.B2(n_177),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_236),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_192),
.C(n_196),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_240),
.C(n_241),
.Y(n_255)
);

OAI32xp33_ASAP7_75t_L g238 ( 
.A1(n_209),
.A2(n_22),
.A3(n_120),
.B1(n_2),
.B2(n_3),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_244),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_214),
.A2(n_29),
.B1(n_27),
.B2(n_25),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_239),
.A2(n_226),
.B1(n_225),
.B2(n_210),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_22),
.C(n_25),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_22),
.C(n_25),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_224),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_22),
.C(n_20),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_247),
.C(n_221),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_218),
.C(n_220),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_211),
.Y(n_249)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_249),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_234),
.B(n_204),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_250),
.B(n_251),
.Y(n_283)
);

XOR2x2_ASAP7_75t_SL g251 ( 
.A(n_237),
.B(n_202),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_203),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_252),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_207),
.Y(n_253)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_260),
.C(n_265),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_243),
.Y(n_259)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_259),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_213),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_264),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_235),
.B(n_209),
.Y(n_262)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_262),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_231),
.B(n_206),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_245),
.Y(n_266)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_266),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_232),
.A2(n_212),
.B(n_201),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_267),
.A2(n_233),
.B(n_240),
.Y(n_272)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_232),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_268),
.A2(n_206),
.B1(n_242),
.B2(n_247),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_14),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_275),
.A2(n_277),
.B1(n_281),
.B2(n_251),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_257),
.A2(n_230),
.B1(n_246),
.B2(n_212),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_276),
.A2(n_280),
.B1(n_284),
.B2(n_262),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_263),
.A2(n_248),
.B1(n_241),
.B2(n_239),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_278),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_254),
.A2(n_238),
.B1(n_236),
.B2(n_20),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_267),
.A2(n_20),
.B1(n_19),
.B2(n_2),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_249),
.A2(n_19),
.B(n_1),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_260),
.C(n_285),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_290),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_276),
.B(n_256),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_287),
.A2(n_289),
.B(n_296),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_288),
.A2(n_298),
.B1(n_297),
.B2(n_5),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_255),
.C(n_250),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_270),
.C(n_255),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_291),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_256),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_292),
.B(n_297),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_265),
.C(n_19),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_294),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_14),
.C(n_1),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_272),
.C(n_274),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_299),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_0),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_282),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_0),
.C(n_1),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_284),
.Y(n_302)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_302),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_282),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_306),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_289),
.A2(n_280),
.B(n_281),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_307),
.A2(n_308),
.B(n_8),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_287),
.A2(n_2),
.B(n_4),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_309),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_311),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_4),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_304),
.B(n_4),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_313),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_6),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_314),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_305),
.B(n_6),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_316),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_7),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_8),
.C(n_9),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_321),
.B(n_302),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_324),
.C(n_325),
.Y(n_329)
);

AOI21xp33_ASAP7_75t_L g323 ( 
.A1(n_317),
.A2(n_301),
.B(n_312),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_323),
.A2(n_316),
.B(n_10),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_320),
.A2(n_9),
.B(n_10),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_327),
.A2(n_318),
.B(n_319),
.Y(n_330)
);

OA21x2_ASAP7_75t_L g332 ( 
.A1(n_330),
.A2(n_331),
.B(n_326),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_332),
.B(n_329),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_328),
.C(n_10),
.Y(n_335)
);

O2A1O1Ixp33_ASAP7_75t_SL g336 ( 
.A1(n_335),
.A2(n_13),
.B(n_10),
.C(n_11),
.Y(n_336)
);

MAJx2_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_9),
.C(n_12),
.Y(n_337)
);

OA21x2_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_12),
.B(n_317),
.Y(n_338)
);


endmodule