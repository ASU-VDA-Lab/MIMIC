module real_jpeg_6383_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_17;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_0),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_0),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_0),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_0),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_0),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_0),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_0),
.B(n_213),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_0),
.B(n_282),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_1),
.B(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_1),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_1),
.B(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_1),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_1),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_1),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_1),
.B(n_224),
.Y(n_223)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_2),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_3),
.B(n_37),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_3),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_3),
.B(n_251),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_3),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_3),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_3),
.B(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_3),
.B(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_3),
.B(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_4),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_5),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_5),
.B(n_31),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_5),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_5),
.B(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_5),
.B(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_5),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_5),
.B(n_431),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_5),
.B(n_444),
.Y(n_443)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_7),
.Y(n_200)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_7),
.Y(n_214)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_7),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_8),
.B(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_8),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_8),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_8),
.B(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_8),
.B(n_412),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_8),
.B(n_427),
.Y(n_426)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_9),
.Y(n_101)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_9),
.Y(n_112)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_9),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_10),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_10),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_10),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_10),
.B(n_115),
.Y(n_114)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_12),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_12),
.Y(n_229)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_12),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_12),
.Y(n_311)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_13),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_13),
.Y(n_151)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_13),
.Y(n_429)
);

BUFx5_ASAP7_75t_L g444 ( 
.A(n_13),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_14),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_14),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_14),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g150 ( 
.A(n_14),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_14),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_14),
.B(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_14),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_15),
.B(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_15),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_15),
.B(n_269),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_15),
.B(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_15),
.B(n_446),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_183),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_181),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_157),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_19),
.B(n_157),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_105),
.C(n_121),
.Y(n_19)
);

FAx1_ASAP7_75t_SL g489 ( 
.A(n_20),
.B(n_105),
.CI(n_121),
.CON(n_489),
.SN(n_489)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_61),
.B1(n_103),
.B2(n_104),
.Y(n_20)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_21),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_43),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_22),
.B(n_43),
.C(n_104),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.C(n_38),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_23),
.B(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_28),
.C(n_32),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_24),
.B(n_51),
.C(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_24),
.A2(n_32),
.B1(n_73),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_24),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_24),
.A2(n_130),
.B1(n_136),
.B2(n_302),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_24),
.A2(n_136),
.B1(n_395),
.B2(n_396),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_25),
.B(n_69),
.Y(n_68)
);

OR2x2_ASAP7_75t_SL g146 ( 
.A(n_25),
.B(n_147),
.Y(n_146)
);

OR2x2_ASAP7_75t_SL g175 ( 
.A(n_25),
.B(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_28),
.A2(n_134),
.B1(n_135),
.B2(n_137),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_28),
.Y(n_134)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx6_ASAP7_75t_L g314 ( 
.A(n_31),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_32),
.A2(n_67),
.B1(n_68),
.B2(n_73),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_32),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_32),
.B(n_63),
.C(n_68),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_32),
.B(n_327),
.C(n_332),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_32),
.A2(n_73),
.B1(n_391),
.B2(n_392),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_33),
.Y(n_196)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_33),
.Y(n_419)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_34),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_35),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_36),
.A2(n_38),
.B1(n_39),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_36),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_38),
.A2(n_39),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_38),
.A2(n_39),
.B1(n_152),
.B2(n_153),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_39),
.B(n_139),
.C(n_152),
.Y(n_138)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_41),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_41),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_42),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_48),
.B1(n_49),
.B2(n_60),
.Y(n_43)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_44),
.B(n_51),
.C(n_54),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_47),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_54),
.B2(n_59),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_50),
.A2(n_51),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_53),
.Y(n_398)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_58),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g287 ( 
.A(n_58),
.Y(n_287)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_74),
.C(n_87),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_62),
.B(n_363),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_67),
.A2(n_68),
.B1(n_114),
.B2(n_116),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_67),
.B(n_108),
.C(n_114),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_67),
.A2(n_68),
.B1(n_130),
.B2(n_302),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_68),
.B(n_130),
.C(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_71),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g283 ( 
.A(n_72),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_72),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_74),
.B(n_87),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.C(n_81),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_75),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_75),
.A2(n_126),
.B1(n_250),
.B2(n_255),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_75),
.B(n_114),
.C(n_250),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_78),
.B(n_81),
.Y(n_127)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_79),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_80),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_80),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_84),
.Y(n_412)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_85),
.Y(n_385)
);

INVx5_ASAP7_75t_L g402 ( 
.A(n_85),
.Y(n_402)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_86),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_98),
.B2(n_102),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_89)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_97),
.C(n_98),
.Y(n_120)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_93),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_94),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_94),
.B(n_281),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_94),
.B(n_281),
.C(n_284),
.Y(n_294)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_101),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_117),
.B2(n_118),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_106),
.B(n_119),
.C(n_120),
.Y(n_159)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_113),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_112),
.Y(n_218)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_114),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_114),
.A2(n_116),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_114),
.A2(n_116),
.B1(n_249),
.B2(n_256),
.Y(n_248)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_138),
.C(n_154),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_122),
.A2(n_123),
.B1(n_365),
.B2(n_366),
.Y(n_364)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_129),
.C(n_133),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_124),
.A2(n_125),
.B1(n_129),
.B2(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_129),
.Y(n_348)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_130),
.Y(n_302)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_133),
.B(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_135),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_136),
.B(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_138),
.B(n_154),
.Y(n_365)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_140),
.B(n_355),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_146),
.C(n_149),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_142),
.B(n_150),
.Y(n_297)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_146),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_146),
.Y(n_296)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx24_ASAP7_75t_SL g492 ( 
.A(n_157),
.Y(n_492)
);

FAx1_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_159),
.CI(n_160),
.CON(n_157),
.SN(n_157)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_170),
.B2(n_180),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_169),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_170),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_177),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_174),
.A2(n_175),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_175),
.B(n_223),
.C(n_228),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_487),
.B(n_490),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

AO21x2_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_358),
.B(n_367),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_342),
.B(n_357),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_317),
.B(n_341),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_188),
.B(n_485),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_289),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_189),
.B(n_289),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_247),
.C(n_276),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_190),
.B(n_340),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_219),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_191),
.B(n_220),
.C(n_231),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_203),
.C(n_209),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_192),
.B(n_337),
.Y(n_336)
);

BUFx24_ASAP7_75t_SL g493 ( 
.A(n_192),
.Y(n_493)
);

FAx1_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_197),
.CI(n_201),
.CON(n_192),
.SN(n_192)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_193),
.B(n_197),
.C(n_201),
.Y(n_288)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_195),
.B(n_241),
.Y(n_240)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_203),
.A2(n_209),
.B1(n_210),
.B2(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_203),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_204),
.B(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_215),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_211),
.A2(n_212),
.B1(n_215),
.B2(n_216),
.Y(n_335)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_214),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_214),
.Y(n_438)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_231),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_227),
.B1(n_228),
.B2(n_230),
.Y(n_222)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_223),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_223),
.A2(n_230),
.B1(n_262),
.B2(n_263),
.Y(n_403)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_239),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_232),
.A2(n_233),
.B(n_234),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_232),
.B(n_240),
.C(n_242),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_238),
.Y(n_234)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_238),
.B(n_419),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_243),
.B(n_387),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_243),
.B(n_401),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_243),
.B(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx6_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_247),
.B(n_276),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_257),
.C(n_259),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_248),
.A2(n_257),
.B1(n_258),
.B2(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_248),
.Y(n_322)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_249),
.Y(n_256)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_250),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_259),
.B(n_321),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_267),
.C(n_272),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_260),
.A2(n_261),
.B1(n_474),
.B2(n_475),
.Y(n_473)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx8_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_267),
.A2(n_268),
.B1(n_272),
.B2(n_273),
.Y(n_475)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_288),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_278),
.B(n_279),
.C(n_288),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_284),
.Y(n_279)
);

INVx8_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_290),
.B(n_292),
.C(n_316),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_303),
.B1(n_315),
.B2(n_316),
.Y(n_291)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_292),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_299),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_294),
.B(n_295),
.C(n_299),
.Y(n_350)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_297),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_303),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_304),
.B(n_306),
.C(n_307),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_308),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_312),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_310),
.B(n_312),
.C(n_353),
.Y(n_352)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_339),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_318),
.B(n_339),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_323),
.C(n_336),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_319),
.A2(n_320),
.B1(n_480),
.B2(n_481),
.Y(n_479)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g480 ( 
.A(n_323),
.B(n_336),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_326),
.C(n_335),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_324),
.B(n_467),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_326),
.B(n_335),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_327),
.A2(n_328),
.B1(n_332),
.B2(n_333),
.Y(n_392)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_343),
.B(n_358),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_344),
.B(n_345),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_345),
.B(n_359),
.Y(n_358)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_345),
.B(n_359),
.Y(n_486)
);

FAx1_ASAP7_75t_SL g345 ( 
.A(n_346),
.B(n_349),
.CI(n_356),
.CON(n_345),
.SN(n_345)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_350),
.B(n_352),
.C(n_354),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_354),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_360),
.B(n_362),
.C(n_364),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_364),
.Y(n_361)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_365),
.Y(n_366)
);

OAI31xp33_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_483),
.A3(n_484),
.B(n_486),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_369),
.A2(n_477),
.B(n_482),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_370),
.A2(n_462),
.B(n_476),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_371),
.A2(n_414),
.B(n_461),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_372),
.B(n_404),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_372),
.B(n_404),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_393),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_390),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_374),
.B(n_390),
.C(n_393),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_381),
.C(n_386),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_375),
.A2(n_376),
.B1(n_381),
.B2(n_382),
.Y(n_406)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx8_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

BUFx8_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g405 ( 
.A(n_386),
.B(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_394),
.B(n_399),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_394),
.B(n_471),
.C(n_472),
.Y(n_470)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx6_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_403),
.Y(n_399)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_400),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_403),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_407),
.C(n_413),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_405),
.B(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_407),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_407),
.A2(n_413),
.B1(n_453),
.B2(n_459),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_411),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_408),
.Y(n_451)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_411),
.Y(n_452)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_413),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_415),
.A2(n_455),
.B(n_460),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_416),
.A2(n_440),
.B(n_454),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_417),
.A2(n_424),
.B(n_439),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_420),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_419),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_422),
.Y(n_420)
);

INVx4_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_425),
.B(n_435),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_425),
.B(n_435),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_426),
.A2(n_430),
.B(n_434),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_426),
.B(n_430),
.Y(n_434)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_434),
.A2(n_442),
.B1(n_448),
.B2(n_449),
.Y(n_441)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_434),
.Y(n_448)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx8_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_441),
.B(n_450),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_441),
.B(n_450),
.Y(n_454)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_442),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_443),
.B(n_445),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_443),
.A2(n_445),
.B(n_448),
.Y(n_456)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_451),
.A2(n_452),
.B(n_453),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_457),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_456),
.B(n_457),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_464),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_463),
.B(n_464),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_465),
.A2(n_466),
.B1(n_468),
.B2(n_469),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_465),
.B(n_470),
.C(n_473),
.Y(n_478)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_473),
.Y(n_469)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_479),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_478),
.B(n_479),
.Y(n_482)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_480),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_489),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_488),
.B(n_489),
.Y(n_490)
);

BUFx24_ASAP7_75t_SL g494 ( 
.A(n_489),
.Y(n_494)
);


endmodule