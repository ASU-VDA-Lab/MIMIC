module fake_jpeg_646_n_156 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_156);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_156;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_19),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

AND2x6_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_15),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_62),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx4f_ASAP7_75t_SL g63 ( 
.A(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_41),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_48),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_71),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_47),
.Y(n_67)
);

CKINVDCx12_ASAP7_75t_R g70 ( 
.A(n_62),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_42),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_75),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_58),
.B(n_52),
.Y(n_75)
);

OR2x2_ASAP7_75t_SL g76 ( 
.A(n_67),
.B(n_64),
.Y(n_76)
);

BUFx8_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_80),
.B(n_86),
.Y(n_96)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_65),
.A2(n_56),
.B1(n_54),
.B2(n_49),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_88),
.B1(n_18),
.B2(n_38),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_51),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_90),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_68),
.A2(n_56),
.B1(n_54),
.B2(n_49),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_84),
.Y(n_106)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_50),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_92),
.B(n_94),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_45),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_98),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_43),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_89),
.A2(n_46),
.B1(n_43),
.B2(n_2),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_95),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_0),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_76),
.A2(n_46),
.B1(n_2),
.B2(n_3),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_105),
.B1(n_5),
.B2(n_6),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_1),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_104),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_1),
.Y(n_104)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_88),
.B(n_4),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_107),
.B(n_4),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_111),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_21),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_102),
.C(n_14),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_100),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_114),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_7),
.Y(n_114)
);

AND2x6_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_23),
.Y(n_115)
);

NOR3xp33_ASAP7_75t_SL g132 ( 
.A(n_115),
.B(n_29),
.C(n_39),
.Y(n_132)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_91),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_102),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_105),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_118)
);

AOI221xp5_ASAP7_75t_L g127 ( 
.A1(n_118),
.A2(n_121),
.B1(n_122),
.B2(n_106),
.C(n_99),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g120 ( 
.A(n_93),
.B(n_22),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_12),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_9),
.B(n_10),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_106),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_28),
.B(n_36),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_125),
.A2(n_30),
.B(n_32),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_116),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_132),
.C(n_135),
.Y(n_141)
);

AOI21xp33_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_130),
.B(n_131),
.Y(n_143)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_137),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_124),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_136),
.A2(n_109),
.B1(n_120),
.B2(n_113),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_140),
.C(n_120),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_110),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_139),
.B(n_142),
.Y(n_145)
);

XOR2x2_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_115),
.Y(n_140)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_143),
.Y(n_144)
);

FAx1_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_147),
.CI(n_135),
.CON(n_149),
.SN(n_149)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_145),
.B(n_146),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_141),
.A2(n_128),
.B1(n_123),
.B2(n_125),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_144),
.B1(n_147),
.B2(n_140),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_148),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_129),
.Y(n_153)
);

NAND4xp25_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_132),
.C(n_137),
.D(n_16),
.Y(n_154)
);

AOI31xp33_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_26),
.A3(n_14),
.B(n_13),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_139),
.Y(n_156)
);


endmodule