module fake_jpeg_15978_n_94 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_94);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_94;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_5),
.B(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_1),
.B(n_7),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_6),
.B(n_3),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_22),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_17),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_25),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_22),
.B(n_19),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_32),
.B(n_36),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_23),
.B(n_19),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_27),
.A2(n_10),
.B1(n_13),
.B2(n_9),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_25),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_46),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_11),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_37),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_32),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_54),
.B1(n_60),
.B2(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_52),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_47),
.A2(n_37),
.B(n_14),
.C(n_12),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_16),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_58),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_20),
.B1(n_27),
.B2(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_43),
.B(n_13),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_30),
.B(n_10),
.C(n_24),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_62),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_54),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_65),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_66),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_72),
.C(n_75),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_49),
.C(n_52),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_49),
.B(n_58),
.Y(n_74)
);

AO21x1_ASAP7_75t_L g77 ( 
.A1(n_74),
.A2(n_68),
.B(n_62),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_67),
.C(n_64),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_77),
.A2(n_81),
.B(n_76),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_9),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_80),
.Y(n_84)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_40),
.B(n_50),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_72),
.C(n_69),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_82),
.A2(n_83),
.B(n_15),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_28),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_2),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_87),
.B(n_88),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_2),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_26),
.C(n_33),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

OAI221xp5_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_91),
.B1(n_34),
.B2(n_35),
.C(n_26),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_34),
.Y(n_94)
);


endmodule