module fake_jpeg_2439_n_226 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_226);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx3_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_20),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

CKINVDCx11_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_24),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_1),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_10),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_14),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_2),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_9),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_8),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_37),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_27),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_55),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_81),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_0),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_80),
.B(n_70),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx5_ASAP7_75t_SL g94 ( 
.A(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_79),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_60),
.B1(n_61),
.B2(n_69),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_91),
.B1(n_93),
.B2(n_72),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_82),
.A2(n_60),
.B1(n_61),
.B2(n_69),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_85),
.A2(n_74),
.B1(n_66),
.B2(n_71),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_92),
.A2(n_95),
.B1(n_84),
.B2(n_79),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_83),
.A2(n_67),
.B1(n_58),
.B2(n_54),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_85),
.A2(n_74),
.B1(n_66),
.B2(n_71),
.Y(n_95)
);

AO22x1_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_53),
.B1(n_67),
.B2(n_73),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_79),
.B(n_73),
.C(n_57),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

INVxp33_ASAP7_75t_SL g131 ( 
.A(n_102),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_96),
.A2(n_83),
.B1(n_59),
.B2(n_76),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_107),
.B1(n_113),
.B2(n_117),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_80),
.B(n_53),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_117),
.B(n_75),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_59),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_68),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_111),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_78),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_108),
.B(n_109),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_79),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_94),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_83),
.B1(n_77),
.B2(n_76),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_89),
.B(n_65),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_94),
.Y(n_128)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_116),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_77),
.C(n_62),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_119),
.B(n_128),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_93),
.B1(n_91),
.B2(n_90),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_123),
.A2(n_127),
.B1(n_138),
.B2(n_132),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_107),
.B1(n_104),
.B2(n_103),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_90),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_130),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_94),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_48),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_1),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_135),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_51),
.Y(n_135)
);

NOR3xp33_ASAP7_75t_SL g136 ( 
.A(n_115),
.B(n_75),
.C(n_3),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_139),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_75),
.B1(n_3),
.B2(n_4),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_2),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_140),
.A2(n_160),
.B1(n_11),
.B2(n_12),
.Y(n_169)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_144),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_50),
.C(n_49),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_147),
.C(n_125),
.Y(n_164)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

NOR3xp33_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_162),
.C(n_136),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_46),
.Y(n_147)
);

OAI32xp33_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_161),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_43),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_156),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_122),
.Y(n_150)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_5),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_152),
.B(n_153),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_119),
.B(n_6),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_135),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_155),
.B(n_163),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_122),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_126),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_158),
.Y(n_183)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_120),
.A2(n_41),
.B1(n_39),
.B2(n_36),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_159),
.A2(n_118),
.B(n_29),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_35),
.B1(n_34),
.B2(n_32),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_128),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_133),
.B(n_31),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_118),
.B(n_11),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_164),
.B(n_165),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_150),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_175),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_181),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_143),
.B(n_28),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_172),
.C(n_176),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_26),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_13),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_25),
.C(n_14),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_13),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_182),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_24),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_161),
.C(n_160),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_145),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_15),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_17),
.Y(n_184)
);

NOR3xp33_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_145),
.C(n_146),
.Y(n_190)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_183),
.Y(n_185)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_185),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_166),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_194),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_21),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_174),
.A2(n_159),
.B1(n_156),
.B2(n_162),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_191),
.A2(n_179),
.B1(n_178),
.B2(n_181),
.Y(n_202)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_197),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_174),
.A2(n_168),
.B(n_180),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_186),
.B(n_171),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_201),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_164),
.C(n_172),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_203),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_176),
.C(n_170),
.Y(n_203)
);

OA21x2_ASAP7_75t_SL g204 ( 
.A1(n_192),
.A2(n_19),
.B(n_20),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_205),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_19),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_207),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_198),
.A2(n_192),
.B1(n_206),
.B2(n_189),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_211),
.Y(n_216)
);

FAx1_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_187),
.CI(n_194),
.CON(n_211),
.SN(n_211)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_200),
.A2(n_189),
.B1(n_193),
.B2(n_22),
.Y(n_212)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_212),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_213),
.B(n_201),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_217),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_211),
.B(n_203),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_218),
.Y(n_220)
);

AOI21x1_ASAP7_75t_L g221 ( 
.A1(n_220),
.A2(n_208),
.B(n_216),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_221),
.B(n_209),
.Y(n_222)
);

A2O1A1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_222),
.A2(n_214),
.B(n_209),
.C(n_219),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_223),
.A2(n_193),
.B(n_22),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_23),
.C(n_208),
.Y(n_225)
);

INVxp33_ASAP7_75t_L g226 ( 
.A(n_225),
.Y(n_226)
);


endmodule