module fake_jpeg_15915_n_157 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_157);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_157;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_5),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx6f_ASAP7_75t_SL g58 ( 
.A(n_28),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_31),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_10),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_71),
.Y(n_79)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_76),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_61),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_78),
.Y(n_102)
);

AO22x1_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_46),
.B1(n_63),
.B2(n_56),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_80),
.A2(n_47),
.B1(n_49),
.B2(n_51),
.Y(n_107)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_86),
.A2(n_62),
.B1(n_46),
.B2(n_63),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_89),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_79),
.A2(n_55),
.B(n_50),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_95),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_57),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_93),
.B(n_94),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_57),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_62),
.Y(n_95)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_60),
.B1(n_56),
.B2(n_48),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_98),
.A2(n_107),
.B1(n_84),
.B2(n_2),
.Y(n_112)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_0),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_75),
.B(n_59),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_6),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_52),
.B1(n_2),
.B2(n_3),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_108),
.A2(n_112),
.B1(n_8),
.B2(n_9),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_114),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_100),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_117),
.A2(n_118),
.B(n_105),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_104),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_121),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_111),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_124),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_113),
.A2(n_110),
.B(n_102),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_125),
.A2(n_126),
.B1(n_117),
.B2(n_96),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_127),
.B(n_98),
.Y(n_135)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_125),
.B1(n_123),
.B2(n_115),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_132),
.A2(n_134),
.B1(n_90),
.B2(n_9),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_120),
.C(n_109),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_133),
.B(n_99),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_127),
.A2(n_96),
.B1(n_97),
.B2(n_116),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_135),
.A2(n_137),
.B(n_131),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_128),
.A2(n_101),
.B(n_103),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_136),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_139),
.A2(n_141),
.B1(n_8),
.B2(n_11),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_140),
.A2(n_133),
.B(n_137),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_144),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_12),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_12),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_145),
.B(n_14),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_13),
.B(n_15),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_150),
.B(n_16),
.Y(n_151)
);

OAI321xp33_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_17),
.A3(n_19),
.B1(n_20),
.B2(n_21),
.C(n_23),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_152),
.A2(n_26),
.B(n_27),
.Y(n_153)
);

AO21x1_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_29),
.B(n_32),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_33),
.C(n_35),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_38),
.C(n_39),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_156),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_157)
);


endmodule