module fake_netlist_1_8034_n_26 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_26);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_26;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
INVx1_ASAP7_75t_L g9 ( .A(n_7), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_5), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_0), .Y(n_11) );
AND2x4_ASAP7_75t_L g12 ( .A(n_4), .B(n_6), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
BUFx3_ASAP7_75t_L g14 ( .A(n_12), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_11), .Y(n_15) );
NOR2xp67_ASAP7_75t_L g16 ( .A(n_9), .B(n_1), .Y(n_16) );
NAND2x1p5_ASAP7_75t_L g17 ( .A(n_16), .B(n_12), .Y(n_17) );
NOR2x1_ASAP7_75t_SL g18 ( .A(n_14), .B(n_10), .Y(n_18) );
AND2x2_ASAP7_75t_L g19 ( .A(n_18), .B(n_14), .Y(n_19) );
OR2x2_ASAP7_75t_L g20 ( .A(n_19), .B(n_17), .Y(n_20) );
HB1xp67_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
AOI211xp5_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_15), .B(n_12), .C(n_13), .Y(n_22) );
NOR2x1_ASAP7_75t_L g23 ( .A(n_22), .B(n_1), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
OAI21x1_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_2), .B(n_3), .Y(n_25) );
INVxp67_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
endmodule