module fake_jpeg_2488_n_438 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_438);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_438;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_SL g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_49),
.B(n_57),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_5),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_50),
.B(n_64),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_51),
.Y(n_143)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx5_ASAP7_75t_SL g112 ( 
.A(n_52),
.Y(n_112)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_55),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_56),
.Y(n_131)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_58),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_59),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_60),
.Y(n_140)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_15),
.B(n_12),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_62),
.B(n_66),
.Y(n_103)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_63),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_18),
.B(n_12),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_67),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_16),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_68),
.B(n_70),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_69),
.Y(n_133)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_71),
.B(n_77),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

BUFx4f_ASAP7_75t_SL g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx2_ASAP7_75t_SL g145 ( 
.A(n_73),
.Y(n_145)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g116 ( 
.A(n_74),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_76),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_20),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_35),
.B(n_9),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_79),
.B(n_80),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_34),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_84),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_23),
.B(n_8),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_87),
.Y(n_153)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_29),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_43),
.B(n_6),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_93),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_22),
.Y(n_92)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_94),
.Y(n_139)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_95),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_40),
.B1(n_47),
.B2(n_30),
.Y(n_113)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_98),
.Y(n_106)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_28),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_65),
.A2(n_21),
.B1(n_30),
.B2(n_47),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_102),
.A2(n_135),
.B1(n_146),
.B2(n_96),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_90),
.A2(n_28),
.B1(n_47),
.B2(n_31),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_115),
.A2(n_130),
.B1(n_137),
.B2(n_144),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_88),
.A2(n_33),
.B1(n_17),
.B2(n_36),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_119),
.A2(n_152),
.B1(n_55),
.B2(n_63),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_123),
.B(n_78),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_48),
.B(n_26),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_132),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_91),
.A2(n_28),
.B1(n_45),
.B2(n_19),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_54),
.B(n_26),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_99),
.A2(n_23),
.B1(n_42),
.B2(n_17),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_76),
.A2(n_19),
.B1(n_39),
.B2(n_38),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_56),
.A2(n_25),
.B1(n_39),
.B2(n_38),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_60),
.A2(n_42),
.B1(n_17),
.B2(n_45),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_67),
.A2(n_31),
.B1(n_25),
.B2(n_15),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_150),
.A2(n_151),
.B1(n_156),
.B2(n_52),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_72),
.A2(n_40),
.B1(n_37),
.B2(n_6),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_58),
.A2(n_37),
.B1(n_6),
.B2(n_2),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_73),
.B(n_0),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_0),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_75),
.A2(n_37),
.B1(n_6),
.B2(n_2),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_111),
.Y(n_158)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_158),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_122),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_159),
.B(n_169),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_73),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_160),
.B(n_178),
.Y(n_206)
);

NAND2x1_ASAP7_75t_SL g161 ( 
.A(n_124),
.B(n_52),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_161),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_162),
.B(n_163),
.Y(n_220)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_166),
.Y(n_233)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

INVx4_ASAP7_75t_SL g203 ( 
.A(n_167),
.Y(n_203)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_111),
.Y(n_168)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_168),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_103),
.B(n_55),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_171),
.Y(n_229)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

OAI21xp33_ASAP7_75t_L g173 ( 
.A1(n_124),
.A2(n_126),
.B(n_132),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_173),
.B(n_179),
.Y(n_228)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_131),
.Y(n_176)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_110),
.Y(n_177)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_177),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_101),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_124),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_107),
.B(n_154),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_183),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_181),
.B(n_182),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_110),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_140),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_185),
.Y(n_227)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_108),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_187),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_120),
.B(n_98),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_92),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_188),
.B(n_190),
.Y(n_231)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_108),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_189),
.B(n_191),
.Y(n_232)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_140),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_120),
.B(n_155),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_192),
.B(n_193),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_106),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_112),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_194),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_120),
.B(n_0),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_195),
.B(n_201),
.Y(n_235)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_114),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_149),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_149),
.Y(n_198)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_138),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_112),
.B1(n_142),
.B2(n_183),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_105),
.A2(n_93),
.B1(n_59),
.B2(n_82),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_200),
.A2(n_148),
.B(n_133),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_106),
.A2(n_51),
.B1(n_87),
.B2(n_85),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_123),
.B(n_0),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_116),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_109),
.C(n_114),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_204),
.B(n_209),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_109),
.C(n_127),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_184),
.A2(n_102),
.B1(n_118),
.B2(n_141),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_211),
.A2(n_219),
.B1(n_177),
.B2(n_165),
.Y(n_246)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_213),
.A2(n_148),
.B1(n_133),
.B2(n_167),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_184),
.A2(n_118),
.B1(n_141),
.B2(n_128),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_215),
.A2(n_222),
.B1(n_201),
.B2(n_183),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_162),
.A2(n_153),
.B1(n_125),
.B2(n_104),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_187),
.A2(n_153),
.B1(n_125),
.B2(n_127),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_117),
.C(n_121),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_225),
.B(n_237),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_161),
.B(n_117),
.C(n_121),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_238),
.B(n_143),
.Y(n_258)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_239),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_202),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_247),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_241),
.A2(n_243),
.B1(n_244),
.B2(n_265),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_236),
.A2(n_170),
.B1(n_163),
.B2(n_182),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_236),
.A2(n_170),
.B1(n_163),
.B2(n_195),
.Y(n_244)
);

MAJx2_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_158),
.C(n_186),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_236),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_246),
.A2(n_215),
.B1(n_222),
.B2(n_210),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_234),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_248),
.A2(n_252),
.B(n_254),
.Y(n_270)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_207),
.Y(n_249)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_204),
.B(n_196),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_250),
.B(n_256),
.Y(n_283)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_251),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_228),
.A2(n_189),
.B(n_105),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_231),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_253),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_220),
.A2(n_100),
.B(n_116),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_206),
.B(n_100),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_255),
.B(n_259),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_172),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_217),
.B(n_175),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_257),
.B(n_263),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_267),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_209),
.B(n_192),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_205),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_261),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_199),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_205),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_264),
.Y(n_279)
);

OA21x2_ASAP7_75t_L g265 ( 
.A1(n_220),
.A2(n_219),
.B(n_211),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_208),
.B(n_190),
.Y(n_266)
);

AOI32xp33_ASAP7_75t_L g278 ( 
.A1(n_266),
.A2(n_227),
.A3(n_210),
.B1(n_214),
.B2(n_223),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_225),
.B(n_136),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_237),
.C(n_224),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_272),
.C(n_273),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_208),
.C(n_235),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_235),
.C(n_220),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_275),
.B(n_258),
.Y(n_314)
);

NOR2xp67_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_216),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_276),
.B(n_245),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_278),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_281),
.A2(n_289),
.B1(n_246),
.B2(n_221),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_252),
.A2(n_229),
.B(n_213),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_285),
.A2(n_254),
.B(n_244),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_242),
.A2(n_229),
.B1(n_214),
.B2(n_226),
.Y(n_289)
);

MAJx2_ASAP7_75t_L g290 ( 
.A(n_262),
.B(n_226),
.C(n_218),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_291),
.C(n_293),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_262),
.B(n_218),
.C(n_221),
.Y(n_291)
);

OAI32xp33_ASAP7_75t_L g292 ( 
.A1(n_242),
.A2(n_266),
.A3(n_256),
.B1(n_257),
.B2(n_250),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_292),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_247),
.B(n_212),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_285),
.A2(n_253),
.B(n_265),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_295),
.B(n_301),
.Y(n_323)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_292),
.Y(n_296)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_296),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_297),
.A2(n_203),
.B1(n_143),
.B2(n_138),
.Y(n_338)
);

NAND2x1p5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_243),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_299),
.B(n_310),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_280),
.B(n_255),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_300),
.B(n_315),
.Y(n_334)
);

AOI32xp33_ASAP7_75t_L g301 ( 
.A1(n_286),
.A2(n_290),
.A3(n_283),
.B1(n_293),
.B2(n_288),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_302),
.Y(n_336)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_283),
.Y(n_303)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_303),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_240),
.Y(n_305)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_284),
.A2(n_265),
.B1(n_241),
.B2(n_267),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_307),
.A2(n_308),
.B1(n_309),
.B2(n_313),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_284),
.A2(n_265),
.B1(n_287),
.B2(n_277),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_270),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_279),
.Y(n_311)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_311),
.Y(n_339)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_279),
.Y(n_312)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_312),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_316),
.Y(n_320)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_271),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_273),
.B(n_245),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_268),
.C(n_272),
.Y(n_319)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_274),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_317),
.B(n_233),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_307),
.A2(n_269),
.B1(n_259),
.B2(n_287),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_318),
.A2(n_330),
.B1(n_333),
.B2(n_335),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_319),
.B(n_325),
.C(n_327),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_320),
.B(n_74),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_298),
.B(n_291),
.Y(n_325)
);

AO21x2_ASAP7_75t_SL g326 ( 
.A1(n_295),
.A2(n_306),
.B(n_296),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_326),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_298),
.B(n_277),
.C(n_269),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_306),
.A2(n_270),
.B1(n_282),
.B2(n_274),
.Y(n_330)
);

OAI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_294),
.A2(n_282),
.B1(n_271),
.B2(n_274),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_331),
.A2(n_310),
.B1(n_317),
.B2(n_305),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_304),
.B(n_249),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_332),
.B(n_341),
.C(n_166),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_294),
.A2(n_251),
.B1(n_239),
.B2(n_198),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_308),
.A2(n_176),
.B1(n_197),
.B2(n_185),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_338),
.A2(n_297),
.B(n_299),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_340),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_304),
.B(n_223),
.C(n_203),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_342),
.A2(n_345),
.B1(n_361),
.B2(n_362),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_322),
.B(n_303),
.Y(n_343)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_343),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_322),
.B(n_314),
.Y(n_346)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_346),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_326),
.A2(n_299),
.B(n_129),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_348),
.A2(n_362),
.B(n_330),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_350),
.B(n_359),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_336),
.B(n_136),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_351),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_337),
.B(n_0),
.Y(n_353)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_353),
.Y(n_373)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_339),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_354),
.B(n_355),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_318),
.B(n_129),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_326),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_356),
.B(n_357),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_334),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_325),
.B(n_93),
.C(n_59),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_358),
.B(n_320),
.Y(n_366)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_328),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_360),
.Y(n_365)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_328),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_326),
.A2(n_69),
.B(n_81),
.Y(n_362)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_363),
.Y(n_385)
);

AO21x1_ASAP7_75t_L g364 ( 
.A1(n_348),
.A2(n_321),
.B(n_323),
.Y(n_364)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_364),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_366),
.Y(n_382)
);

XNOR2x1_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_329),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_372),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_357),
.B(n_327),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_374),
.B(n_378),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_344),
.B(n_332),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_375),
.B(n_344),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_377),
.A2(n_347),
.B1(n_356),
.B2(n_349),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_343),
.Y(n_378)
);

A2O1A1O1Ixp25_ASAP7_75t_L g379 ( 
.A1(n_346),
.A2(n_329),
.B(n_319),
.C(n_341),
.D(n_324),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_379),
.A2(n_350),
.B(n_347),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_381),
.B(n_384),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_370),
.B(n_368),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_375),
.B(n_354),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_386),
.B(n_393),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_388),
.A2(n_352),
.B1(n_335),
.B2(n_373),
.Y(n_405)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_376),
.Y(n_389)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_389),
.Y(n_401)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_365),
.Y(n_390)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_390),
.Y(n_406)
);

OAI221xp5_ASAP7_75t_L g395 ( 
.A1(n_391),
.A2(n_364),
.B1(n_376),
.B2(n_363),
.C(n_352),
.Y(n_395)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_365),
.Y(n_392)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_392),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_367),
.B(n_359),
.C(n_358),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_391),
.B(n_367),
.C(n_372),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_394),
.B(n_396),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_395),
.B(n_371),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_382),
.B(n_342),
.C(n_349),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_383),
.B(n_349),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_397),
.B(n_399),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_387),
.B(n_355),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_387),
.B(n_361),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_400),
.B(n_404),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_380),
.B(n_333),
.Y(n_404)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_405),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_397),
.A2(n_389),
.B(n_385),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_408),
.A2(n_409),
.B(n_415),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g409 ( 
.A(n_401),
.B(n_373),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_403),
.B(n_388),
.C(n_393),
.Y(n_410)
);

OR2x2_ASAP7_75t_L g421 ( 
.A(n_410),
.B(n_396),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_402),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_412),
.B(n_360),
.Y(n_422)
);

AOI21xp33_ASAP7_75t_L g415 ( 
.A1(n_406),
.A2(n_385),
.B(n_379),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_416),
.A2(n_371),
.B(n_404),
.Y(n_425)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_398),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_417),
.B(n_399),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_410),
.B(n_407),
.Y(n_418)
);

AOI21xp33_ASAP7_75t_L g426 ( 
.A1(n_418),
.A2(n_420),
.B(n_422),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_414),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_421),
.B(n_425),
.C(n_411),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_423),
.B(n_424),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_408),
.A2(n_394),
.B(n_369),
.Y(n_424)
);

NOR2xp67_ASAP7_75t_L g431 ( 
.A(n_427),
.B(n_429),
.Y(n_431)
);

NOR2xp67_ASAP7_75t_L g428 ( 
.A(n_419),
.B(n_413),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_428),
.A2(n_409),
.B(n_351),
.Y(n_432)
);

BUFx24_ASAP7_75t_SL g429 ( 
.A(n_421),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_432),
.A2(n_433),
.B(n_426),
.Y(n_434)
);

A2O1A1O1Ixp25_ASAP7_75t_L g433 ( 
.A1(n_430),
.A2(n_353),
.B(n_340),
.C(n_4),
.D(n_3),
.Y(n_433)
);

OAI21xp33_ASAP7_75t_L g436 ( 
.A1(n_434),
.A2(n_435),
.B(n_4),
.Y(n_436)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_431),
.B(n_1),
.Y(n_435)
);

AO221x1_ASAP7_75t_L g437 ( 
.A1(n_436),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.C(n_212),
.Y(n_437)
);

NOR3xp33_ASAP7_75t_SL g438 ( 
.A(n_437),
.B(n_1),
.C(n_3),
.Y(n_438)
);


endmodule