module fake_jpeg_11617_n_374 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_374);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_374;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_SL g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_10),
.B(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_3),
.B(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx9p33_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_40),
.B(n_41),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_53),
.B(n_65),
.Y(n_117)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

BUFx4f_ASAP7_75t_SL g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_7),
.B1(n_15),
.B2(n_12),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_56),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_135)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_26),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_63),
.B(n_85),
.Y(n_109)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_64),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_21),
.B(n_16),
.Y(n_65)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_21),
.B(n_16),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_73),
.B(n_78),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_75),
.Y(n_146)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_76),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_30),
.B(n_11),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_79),
.Y(n_158)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_82),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_18),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_88),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_30),
.B(n_11),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_90),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

BUFx2_ASAP7_75t_SL g139 ( 
.A(n_91),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_31),
.B(n_10),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_93),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_31),
.B(n_7),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_94),
.B(n_95),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_99),
.Y(n_115)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_98),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_18),
.B(n_0),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_23),
.B(n_0),
.C(n_1),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_101),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g101 ( 
.A1(n_33),
.A2(n_0),
.B(n_2),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_102),
.B(n_104),
.Y(n_153)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_5),
.Y(n_136)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_80),
.A2(n_66),
.B1(n_83),
.B2(n_27),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_105),
.A2(n_118),
.B1(n_124),
.B2(n_132),
.Y(n_168)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_58),
.A2(n_32),
.B1(n_48),
.B2(n_47),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_106),
.A2(n_139),
.B(n_140),
.C(n_125),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_69),
.A2(n_27),
.B1(n_48),
.B2(n_47),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_72),
.A2(n_32),
.B1(n_36),
.B2(n_22),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_119),
.A2(n_140),
.B1(n_125),
.B2(n_148),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_59),
.A2(n_49),
.B1(n_33),
.B2(n_39),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_120),
.A2(n_133),
.B1(n_159),
.B2(n_160),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_69),
.A2(n_36),
.B1(n_103),
.B2(n_99),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g131 ( 
.A1(n_98),
.A2(n_49),
.B(n_4),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_131),
.A2(n_98),
.B(n_121),
.C(n_101),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_81),
.A2(n_39),
.B1(n_35),
.B2(n_28),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_60),
.A2(n_35),
.B1(n_28),
.B2(n_26),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_160),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_136),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_96),
.A2(n_43),
.B1(n_26),
.B2(n_6),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_144),
.A2(n_154),
.B1(n_155),
.B2(n_108),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_54),
.A2(n_71),
.B1(n_94),
.B2(n_90),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_89),
.A2(n_77),
.B1(n_87),
.B2(n_86),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_55),
.B(n_5),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_157),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_95),
.B(n_6),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_74),
.A2(n_79),
.B1(n_82),
.B2(n_84),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_56),
.A2(n_26),
.B1(n_6),
.B2(n_43),
.Y(n_160)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_163),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_117),
.B(n_111),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_164),
.B(n_169),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_6),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_165),
.B(n_186),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_121),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_166),
.B(n_167),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_110),
.B(n_43),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_126),
.Y(n_170)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_170),
.Y(n_221)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_135),
.A2(n_43),
.B1(n_106),
.B2(n_112),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_172),
.A2(n_183),
.B1(n_194),
.B2(n_201),
.Y(n_214)
);

NAND2xp33_ASAP7_75t_SL g173 ( 
.A(n_121),
.B(n_115),
.Y(n_173)
);

OAI21xp33_ASAP7_75t_L g227 ( 
.A1(n_173),
.A2(n_192),
.B(n_204),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_121),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_174),
.B(n_176),
.Y(n_233)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_107),
.Y(n_175)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_175),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_153),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_107),
.Y(n_177)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_114),
.Y(n_178)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_178),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_128),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_179),
.B(n_188),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_181),
.A2(n_200),
.B1(n_205),
.B2(n_208),
.Y(n_235)
);

BUFx8_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_182),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_106),
.A2(n_115),
.B1(n_142),
.B2(n_148),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_190),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_109),
.B(n_116),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_185),
.B(n_187),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_150),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_127),
.B(n_138),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_145),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_122),
.B(n_131),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_189),
.B(n_191),
.Y(n_249)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_150),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_122),
.B(n_106),
.Y(n_191)
);

NAND2xp33_ASAP7_75t_SL g192 ( 
.A(n_119),
.B(n_143),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_108),
.A2(n_137),
.B1(n_161),
.B2(n_141),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_195),
.A2(n_194),
.B1(n_162),
.B2(n_192),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_122),
.B(n_123),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_197),
.B(n_206),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_129),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_198),
.B(n_199),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_123),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_141),
.A2(n_129),
.B1(n_142),
.B2(n_149),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_149),
.A2(n_147),
.B1(n_151),
.B2(n_158),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_126),
.A2(n_130),
.B1(n_147),
.B2(n_151),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_202),
.A2(n_195),
.B1(n_191),
.B2(n_170),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_113),
.B(n_158),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_207),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_130),
.A2(n_45),
.B1(n_80),
.B2(n_83),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_110),
.B(n_117),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_146),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_126),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_146),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_209),
.B(n_212),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_121),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_169),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_119),
.A2(n_45),
.B1(n_80),
.B2(n_83),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_211),
.B(n_168),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_134),
.A2(n_121),
.B(n_112),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_213),
.A2(n_182),
.B1(n_170),
.B2(n_208),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_217),
.A2(n_224),
.B1(n_238),
.B2(n_202),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_179),
.B(n_206),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_219),
.B(n_231),
.Y(n_252)
);

NOR2x1_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_165),
.Y(n_222)
);

NOR2x1_ASAP7_75t_L g280 ( 
.A(n_222),
.B(n_226),
.Y(n_280)
);

NOR2x1_ASAP7_75t_R g226 ( 
.A(n_173),
.B(n_174),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_187),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_230),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_186),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_176),
.B(n_164),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_172),
.A2(n_166),
.B1(n_212),
.B2(n_194),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_201),
.A2(n_162),
.B1(n_163),
.B2(n_207),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_242),
.A2(n_244),
.B1(n_214),
.B2(n_239),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_180),
.B(n_203),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_245),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_171),
.A2(n_209),
.B1(n_190),
.B2(n_175),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_180),
.B(n_196),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_246),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_197),
.B(n_178),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_188),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_251),
.A2(n_222),
.B(n_226),
.Y(n_300)
);

FAx1_ASAP7_75t_SL g254 ( 
.A(n_243),
.B(n_204),
.CI(n_184),
.CON(n_254),
.SN(n_254)
);

FAx1_ASAP7_75t_SL g293 ( 
.A(n_254),
.B(n_226),
.CI(n_223),
.CON(n_293),
.SN(n_293)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_215),
.Y(n_255)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_255),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_199),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_256),
.Y(n_281)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_215),
.Y(n_257)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_257),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_215),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_258),
.B(n_268),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_259),
.A2(n_235),
.B(n_234),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_238),
.A2(n_217),
.B1(n_249),
.B2(n_230),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_260),
.A2(n_267),
.B1(n_272),
.B2(n_246),
.Y(n_297)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_215),
.Y(n_261)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_261),
.Y(n_301)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_228),
.Y(n_262)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_262),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_219),
.B(n_177),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_274),
.C(n_247),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_265),
.B(n_276),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_249),
.A2(n_182),
.B1(n_208),
.B2(n_227),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_228),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_182),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_270),
.Y(n_295)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_232),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_271),
.B(n_275),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_216),
.A2(n_214),
.B1(n_242),
.B2(n_248),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_273),
.A2(n_277),
.B1(n_216),
.B2(n_220),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_216),
.B(n_248),
.C(n_233),
.Y(n_274)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_221),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_240),
.B(n_229),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_213),
.A2(n_225),
.B1(n_233),
.B2(n_239),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_240),
.B(n_245),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_278),
.B(n_279),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_248),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_248),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_283),
.B(n_274),
.C(n_264),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_285),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_273),
.A2(n_216),
.B1(n_223),
.B2(n_213),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_286),
.A2(n_296),
.B1(n_297),
.B2(n_300),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_253),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_291),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_289),
.B(n_280),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_253),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_252),
.B(n_231),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_293),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_252),
.B(n_225),
.Y(n_294)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_294),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_277),
.A2(n_236),
.B1(n_222),
.B2(n_218),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_303),
.A2(n_258),
.B1(n_261),
.B2(n_257),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_305),
.B(n_307),
.C(n_310),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_263),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_280),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_299),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_311),
.B(n_318),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_283),
.B(n_279),
.C(n_260),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_284),
.Y(n_325)
);

NAND3xp33_ASAP7_75t_L g313 ( 
.A(n_292),
.B(n_266),
.C(n_276),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_313),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_287),
.B(n_278),
.Y(n_314)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_314),
.Y(n_328)
);

AOI322xp5_ASAP7_75t_SL g315 ( 
.A1(n_294),
.A2(n_236),
.A3(n_254),
.B1(n_265),
.B2(n_267),
.C1(n_280),
.C2(n_272),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_315),
.Y(n_327)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_302),
.Y(n_317)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_317),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_281),
.B(n_241),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_319),
.B(n_321),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_320),
.B(n_286),
.Y(n_330)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_302),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_316),
.A2(n_297),
.B(n_300),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_322),
.B(n_323),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_316),
.A2(n_284),
.B(n_288),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_325),
.B(n_329),
.C(n_330),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_303),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_304),
.A2(n_291),
.B1(n_296),
.B2(n_285),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_331),
.A2(n_311),
.B1(n_312),
.B2(n_298),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_306),
.A2(n_288),
.B(n_295),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_333),
.B(n_295),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_334),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_336),
.A2(n_346),
.B1(n_332),
.B2(n_322),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_337),
.B(n_347),
.Y(n_354)
);

NOR3xp33_ASAP7_75t_SL g339 ( 
.A(n_328),
.B(n_304),
.C(n_282),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_339),
.B(n_340),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_324),
.B(n_335),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_326),
.B(n_325),
.C(n_305),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_342),
.B(n_343),
.C(n_329),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_326),
.B(n_307),
.C(n_310),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_344),
.B(n_345),
.Y(n_353)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_335),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_327),
.A2(n_318),
.B(n_308),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_332),
.A2(n_308),
.B1(n_301),
.B2(n_298),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_348),
.A2(n_355),
.B1(n_353),
.B2(n_354),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_349),
.B(n_352),
.Y(n_356)
);

OAI31xp33_ASAP7_75t_L g351 ( 
.A1(n_338),
.A2(n_331),
.A3(n_323),
.B(n_309),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_351),
.A2(n_327),
.B(n_282),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_342),
.B(n_330),
.C(n_333),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_347),
.A2(n_301),
.B1(n_290),
.B2(n_317),
.Y(n_355)
);

A2O1A1Ixp33_ASAP7_75t_SL g357 ( 
.A1(n_351),
.A2(n_290),
.B(n_251),
.C(n_339),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_358),
.B(n_360),
.Y(n_363)
);

AOI31xp67_ASAP7_75t_SL g359 ( 
.A1(n_350),
.A2(n_293),
.A3(n_336),
.B(n_254),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_359),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_352),
.A2(n_343),
.B(n_341),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_361),
.B(n_349),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_362),
.A2(n_355),
.B(n_357),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_356),
.B(n_354),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_365),
.B(n_299),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_363),
.A2(n_341),
.B(n_357),
.Y(n_366)
);

OR2x2_ASAP7_75t_L g369 ( 
.A(n_366),
.B(n_367),
.Y(n_369)
);

INVxp33_ASAP7_75t_SL g370 ( 
.A(n_368),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_369),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_371),
.B(n_372),
.C(n_364),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_370),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_373),
.B(n_321),
.Y(n_374)
);


endmodule