module fake_netlist_1_10010_n_36 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_36);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_36;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx3_ASAP7_75t_L g10 ( .A(n_3), .Y(n_10) );
OR2x2_ASAP7_75t_L g11 ( .A(n_7), .B(n_0), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_0), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_6), .Y(n_13) );
INVx3_ASAP7_75t_L g14 ( .A(n_2), .Y(n_14) );
INVx3_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
AOI22xp5_ASAP7_75t_L g16 ( .A1(n_10), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_16) );
INVx8_ASAP7_75t_L g17 ( .A(n_10), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_10), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_14), .Y(n_19) );
AOI21x1_ASAP7_75t_L g20 ( .A1(n_18), .A2(n_13), .B(n_11), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_17), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_17), .Y(n_22) );
BUFx2_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_22), .B(n_19), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_24), .B(n_22), .Y(n_25) );
AND2x4_ASAP7_75t_SL g26 ( .A(n_23), .B(n_16), .Y(n_26) );
A2O1A1Ixp33_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_13), .B(n_11), .C(n_14), .Y(n_27) );
OAI32xp33_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_15), .A3(n_14), .B1(n_12), .B2(n_20), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
CKINVDCx20_ASAP7_75t_R g30 ( .A(n_28), .Y(n_30) );
NAND2x1_ASAP7_75t_SL g31 ( .A(n_29), .B(n_4), .Y(n_31) );
AO22x2_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_5), .B1(n_8), .B2(n_9), .Y(n_32) );
INVx1_ASAP7_75t_SL g33 ( .A(n_31), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
HB1xp67_ASAP7_75t_L g35 ( .A(n_34), .Y(n_35) );
AOI22x1_ASAP7_75t_L g36 ( .A1(n_35), .A2(n_32), .B1(n_34), .B2(n_33), .Y(n_36) );
endmodule