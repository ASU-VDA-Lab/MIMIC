module fake_jpeg_23295_n_51 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_51);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_51;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx11_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

AOI22xp5_ASAP7_75t_L g9 ( 
.A1(n_3),
.A2(n_4),
.B1(n_5),
.B2(n_1),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx4_ASAP7_75t_SL g11 ( 
.A(n_4),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_9),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_17),
.B(n_20),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g18 ( 
.A1(n_11),
.A2(n_14),
.B1(n_7),
.B2(n_9),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_18),
.A2(n_23),
.B1(n_10),
.B2(n_13),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_1),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_13),
.C(n_10),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_12),
.B(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_7),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_29),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_17),
.C(n_22),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_19),
.B1(n_21),
.B2(n_24),
.Y(n_36)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_35),
.C(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_31),
.B1(n_25),
.B2(n_30),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_28),
.B(n_25),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_40),
.C(n_27),
.Y(n_42)
);

FAx1_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_8),
.CI(n_15),
.CON(n_44),
.SN(n_44)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_36),
.C(n_32),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_42),
.C(n_8),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_44),
.B(n_15),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_45),
.A2(n_47),
.B(n_41),
.Y(n_48)
);

BUFx24_ASAP7_75t_SL g50 ( 
.A(n_48),
.Y(n_50)
);

INVxp33_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

AOI21x1_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_49),
.B(n_44),
.Y(n_51)
);


endmodule