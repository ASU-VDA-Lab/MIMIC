module real_aes_12797_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_635;
wire n_287;
wire n_503;
wire n_673;
wire n_386;
wire n_905;
wire n_518;
wire n_254;
wire n_792;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_537;
wire n_551;
wire n_320;
wire n_884;
wire n_560;
wire n_660;
wire n_260;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_932;
wire n_235;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_478;
wire n_356;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_938;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_931;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_656;
wire n_316;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_298;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_922;
wire n_926;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_237;
wire n_797;
wire n_862;
INVx2_ASAP7_75t_SL g582 ( .A(n_0), .Y(n_582) );
AOI21xp33_ASAP7_75t_L g933 ( .A1(n_1), .A2(n_537), .B(n_934), .Y(n_933) );
CKINVDCx5p33_ASAP7_75t_R g699 ( .A(n_2), .Y(n_699) );
OA21x2_ASAP7_75t_L g157 ( .A1(n_3), .A2(n_50), .B(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g172 ( .A(n_3), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g680 ( .A(n_4), .B(n_230), .Y(n_680) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_5), .B(n_224), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_6), .B(n_149), .Y(n_148) );
NAND2xp33_ASAP7_75t_L g204 ( .A(n_7), .B(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g648 ( .A(n_8), .B(n_210), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_9), .B(n_247), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_10), .B(n_185), .Y(n_242) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_11), .A2(n_65), .B1(n_550), .B2(n_551), .Y(n_549) );
INVx1_ASAP7_75t_L g551 ( .A(n_11), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_12), .B(n_152), .Y(n_675) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_13), .Y(n_169) );
INVx1_ASAP7_75t_L g137 ( .A(n_14), .Y(n_137) );
BUFx3_ASAP7_75t_L g141 ( .A(n_14), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_15), .B(n_209), .Y(n_682) );
A2O1A1Ixp33_ASAP7_75t_L g325 ( .A1(n_16), .A2(n_276), .B(n_326), .C(n_328), .Y(n_325) );
BUFx10_ASAP7_75t_L g121 ( .A(n_17), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_18), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_19), .B(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_20), .B(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_21), .B(n_232), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g316 ( .A1(n_22), .A2(n_206), .B(n_317), .C(n_318), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g668 ( .A(n_23), .Y(n_668) );
NAND3xp33_ASAP7_75t_L g628 ( .A(n_24), .B(n_270), .C(n_626), .Y(n_628) );
AND2x2_ASAP7_75t_L g220 ( .A(n_25), .B(n_219), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_26), .B(n_149), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_27), .B(n_209), .Y(n_248) );
AND2x2_ASAP7_75t_L g537 ( .A(n_28), .B(n_538), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_29), .A2(n_74), .B1(n_186), .B2(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g164 ( .A(n_30), .Y(n_164) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_31), .A2(n_75), .B1(n_522), .B2(n_523), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_31), .Y(n_522) );
INVx1_ASAP7_75t_L g155 ( .A(n_32), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_33), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g939 ( .A(n_34), .Y(n_939) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_35), .B(n_186), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_36), .B(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g110 ( .A(n_37), .Y(n_110) );
AND3x2_ASAP7_75t_L g937 ( .A(n_37), .B(n_111), .C(n_544), .Y(n_937) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_38), .B(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_39), .B(n_276), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_40), .B(n_209), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_41), .B(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g702 ( .A(n_42), .B(n_135), .Y(n_702) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_43), .Y(n_327) );
AND2x4_ASAP7_75t_L g163 ( .A(n_44), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_45), .B(n_209), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_46), .B(n_219), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_47), .B(n_209), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g184 ( .A1(n_48), .A2(n_87), .B1(n_185), .B2(n_186), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_49), .A2(n_548), .B1(n_549), .B2(n_552), .Y(n_547) );
CKINVDCx5p33_ASAP7_75t_R g552 ( .A(n_49), .Y(n_552) );
INVx1_ASAP7_75t_L g171 ( .A(n_50), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g644 ( .A(n_51), .Y(n_644) );
A2O1A1Ixp33_ASAP7_75t_L g579 ( .A1(n_52), .A2(n_580), .B(n_581), .C(n_583), .Y(n_579) );
INVx1_ASAP7_75t_L g158 ( .A(n_53), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_54), .B(n_209), .Y(n_703) );
AND2x4_ASAP7_75t_L g108 ( .A(n_55), .B(n_109), .Y(n_108) );
INVx3_ASAP7_75t_L g666 ( .A(n_56), .Y(n_666) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_57), .Y(n_115) );
NOR2xp67_ASAP7_75t_L g531 ( .A(n_57), .B(n_77), .Y(n_531) );
AND2x2_ASAP7_75t_L g263 ( .A(n_58), .B(n_210), .Y(n_263) );
INVx1_ASAP7_75t_L g109 ( .A(n_59), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_60), .B(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_61), .B(n_593), .Y(n_598) );
NAND2x1_ASAP7_75t_L g275 ( .A(n_62), .B(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_63), .B(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g678 ( .A(n_64), .Y(n_678) );
INVx1_ASAP7_75t_L g550 ( .A(n_65), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_66), .B(n_139), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_67), .B(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g112 ( .A(n_68), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_69), .B(n_185), .Y(n_622) );
CKINVDCx5p33_ASAP7_75t_R g639 ( .A(n_70), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_71), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_72), .B(n_270), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_73), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g523 ( .A(n_75), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_76), .B(n_255), .Y(n_262) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_77), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_78), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_79), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_80), .B(n_247), .Y(n_271) );
NAND2xp33_ASAP7_75t_SL g146 ( .A(n_81), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g134 ( .A(n_82), .B(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g573 ( .A(n_83), .Y(n_573) );
CKINVDCx5p33_ASAP7_75t_R g645 ( .A(n_84), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_85), .B(n_139), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_86), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g144 ( .A(n_88), .Y(n_144) );
BUFx3_ASAP7_75t_L g152 ( .A(n_88), .Y(n_152) );
INVx1_ASAP7_75t_L g181 ( .A(n_88), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_89), .B(n_261), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_90), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_91), .B(n_185), .Y(n_697) );
INVx1_ASAP7_75t_L g664 ( .A(n_92), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g611 ( .A(n_93), .B(n_245), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_94), .B(n_210), .Y(n_614) );
NAND2xp33_ASAP7_75t_L g198 ( .A(n_95), .B(n_199), .Y(n_198) );
OAI21xp5_ASAP7_75t_L g122 ( .A1(n_96), .A2(n_123), .B(n_532), .Y(n_122) );
INVx1_ASAP7_75t_L g534 ( .A(n_96), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_97), .B(n_597), .Y(n_596) );
CKINVDCx5p33_ASAP7_75t_R g660 ( .A(n_98), .Y(n_660) );
INVx1_ASAP7_75t_L g656 ( .A(n_99), .Y(n_656) );
CKINVDCx5p33_ASAP7_75t_R g641 ( .A(n_100), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_101), .B(n_135), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_102), .B(n_593), .Y(n_592) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_118), .B(n_938), .Y(n_103) );
BUFx5_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
BUFx10_ASAP7_75t_L g940 ( .A(n_105), .Y(n_940) );
AND2x4_ASAP7_75t_L g105 ( .A(n_106), .B(n_113), .Y(n_105) );
NOR3xp33_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .C(n_111), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_110), .B(n_531), .Y(n_530) );
BUFx2_ASAP7_75t_L g559 ( .A(n_110), .Y(n_559) );
AND2x2_ASAP7_75t_L g543 ( .A(n_111), .B(n_544), .Y(n_543) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g529 ( .A(n_112), .Y(n_529) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AO21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_122), .B(n_540), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_120), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx3_ASAP7_75t_L g545 ( .A(n_121), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_121), .B(n_937), .Y(n_936) );
OR2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_525), .Y(n_123) );
AOI21xp33_ASAP7_75t_SL g532 ( .A1(n_124), .A2(n_533), .B(n_537), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_520), .B1(n_521), .B2(n_524), .Y(n_124) );
INVx2_ASAP7_75t_L g524 ( .A(n_125), .Y(n_524) );
AO22x2_ASAP7_75t_L g554 ( .A1(n_125), .A2(n_555), .B1(n_556), .B2(n_560), .Y(n_554) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_403), .Y(n_125) );
NOR4xp25_ASAP7_75t_L g126 ( .A(n_127), .B(n_303), .C(n_349), .D(n_389), .Y(n_126) );
OAI21xp33_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_212), .B(n_280), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_165), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_129), .B(n_380), .Y(n_423) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g483 ( .A(n_130), .B(n_380), .Y(n_483) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_131), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_131), .B(n_296), .Y(n_494) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g290 ( .A(n_132), .B(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g294 ( .A(n_132), .Y(n_294) );
AND2x2_ASAP7_75t_L g365 ( .A(n_132), .B(n_192), .Y(n_365) );
AND2x2_ASAP7_75t_L g393 ( .A(n_132), .B(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g417 ( .A(n_132), .B(n_332), .Y(n_417) );
AND2x2_ASAP7_75t_L g447 ( .A(n_132), .B(n_332), .Y(n_447) );
AO31x2_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_145), .A3(n_153), .B(n_159), .Y(n_132) );
AO21x1_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_138), .B(n_142), .Y(n_133) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g147 ( .A(n_136), .Y(n_147) );
INVx1_ASAP7_75t_L g199 ( .A(n_136), .Y(n_199) );
INVx2_ASAP7_75t_L g230 ( .A(n_136), .Y(n_230) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g226 ( .A(n_137), .Y(n_226) );
INVx2_ASAP7_75t_L g274 ( .A(n_139), .Y(n_274) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g191 ( .A(n_140), .Y(n_191) );
INVx2_ASAP7_75t_L g197 ( .A(n_140), .Y(n_197) );
INVx2_ASAP7_75t_L g261 ( .A(n_140), .Y(n_261) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_141), .Y(n_150) );
INVx2_ASAP7_75t_L g187 ( .A(n_141), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_142), .A2(n_229), .B(n_231), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_142), .A2(n_244), .B(n_246), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_142), .A2(n_269), .B(n_271), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_142), .A2(n_611), .B(n_612), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g679 ( .A1(n_142), .A2(n_680), .B(n_681), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_142), .A2(n_696), .B(n_697), .Y(n_695) );
BUFx10_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g626 ( .A(n_143), .Y(n_626) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx3_ASAP7_75t_L g584 ( .A(n_144), .Y(n_584) );
AO21x1_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_148), .B(n_151), .Y(n_145) );
INVx2_ASAP7_75t_L g247 ( .A(n_147), .Y(n_247) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g185 ( .A(n_150), .Y(n_185) );
INVx2_ASAP7_75t_L g203 ( .A(n_150), .Y(n_203) );
INVx2_ASAP7_75t_L g232 ( .A(n_150), .Y(n_232) );
INVx3_ASAP7_75t_L g572 ( .A(n_150), .Y(n_572) );
INVx3_ASAP7_75t_L g638 ( .A(n_150), .Y(n_638) );
INVx2_ASAP7_75t_L g701 ( .A(n_150), .Y(n_701) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_151), .A2(n_241), .B(n_242), .Y(n_240) );
O2A1O1Ixp5_ASAP7_75t_L g698 ( .A1(n_151), .A2(n_699), .B(n_700), .C(n_702), .Y(n_698) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g200 ( .A(n_152), .Y(n_200) );
INVx2_ASAP7_75t_L g207 ( .A(n_152), .Y(n_207) );
AOI211x1_ASAP7_75t_L g221 ( .A1(n_152), .A2(n_220), .B(n_222), .C(n_228), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_152), .B(n_658), .Y(n_657) );
NOR3xp33_ASAP7_75t_L g663 ( .A(n_152), .B(n_658), .C(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_154), .A2(n_160), .B(n_162), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
INVxp33_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx2_ASAP7_75t_L g161 ( .A(n_157), .Y(n_161) );
INVx1_ASAP7_75t_L g211 ( .A(n_157), .Y(n_211) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_157), .Y(n_219) );
INVx1_ASAP7_75t_L g173 ( .A(n_158), .Y(n_173) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx3_ASAP7_75t_L g193 ( .A(n_161), .Y(n_193) );
OAI21x1_ASAP7_75t_L g194 ( .A1(n_162), .A2(n_195), .B(n_201), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_162), .A2(n_218), .B(n_220), .Y(n_217) );
OAI21x1_ASAP7_75t_L g239 ( .A1(n_162), .A2(n_240), .B(n_243), .Y(n_239) );
OAI21x1_ASAP7_75t_L g606 ( .A1(n_162), .A2(n_607), .B(n_610), .Y(n_606) );
OAI21x1_ASAP7_75t_L g672 ( .A1(n_162), .A2(n_673), .B(n_679), .Y(n_672) );
BUFx6f_ASAP7_75t_SL g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g177 ( .A(n_163), .Y(n_177) );
INVx1_ASAP7_75t_L g252 ( .A(n_163), .Y(n_252) );
INVx2_ASAP7_75t_L g278 ( .A(n_163), .Y(n_278) );
INVx3_ASAP7_75t_L g658 ( .A(n_163), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_165), .B(n_393), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_165), .B(n_338), .Y(n_420) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_192), .Y(n_165) );
AND2x2_ASAP7_75t_L g293 ( .A(n_166), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g289 ( .A(n_167), .Y(n_289) );
AND2x2_ASAP7_75t_L g331 ( .A(n_167), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g339 ( .A(n_167), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g360 ( .A(n_167), .Y(n_360) );
AND2x2_ASAP7_75t_L g380 ( .A(n_167), .B(n_192), .Y(n_380) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_167), .Y(n_416) );
INVxp67_ASAP7_75t_L g446 ( .A(n_167), .Y(n_446) );
OR2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_174), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_170), .B(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g323 ( .A(n_170), .Y(n_323) );
AO21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_173), .Y(n_170) );
AOI21x1_ASAP7_75t_L g183 ( .A1(n_171), .A2(n_172), .B(n_173), .Y(n_183) );
OAI22xp5_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_184), .B1(n_188), .B2(n_190), .Y(n_174) );
NAND3xp33_ASAP7_75t_L g175 ( .A(n_176), .B(n_178), .C(n_182), .Y(n_175) );
NAND3xp33_ASAP7_75t_L g188 ( .A(n_176), .B(n_182), .C(n_189), .Y(n_188) );
BUFx2_ASAP7_75t_L g647 ( .A(n_176), .Y(n_647) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
OAI21xp33_ASAP7_75t_L g585 ( .A1(n_177), .A2(n_323), .B(n_578), .Y(n_585) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_179), .B(n_658), .Y(n_661) );
NOR3xp33_ASAP7_75t_L g665 ( .A(n_179), .B(n_658), .C(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g328 ( .A(n_180), .Y(n_328) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
BUFx3_ASAP7_75t_L g189 ( .A(n_181), .Y(n_189) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_182), .Y(n_652) );
NOR2xp33_ASAP7_75t_SL g667 ( .A(n_182), .B(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_186), .B(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g205 ( .A(n_187), .Y(n_205) );
INVx1_ASAP7_75t_L g270 ( .A(n_187), .Y(n_270) );
INVx2_ASAP7_75t_L g257 ( .A(n_189), .Y(n_257) );
O2A1O1Ixp5_ASAP7_75t_L g272 ( .A1(n_189), .A2(n_273), .B(n_274), .C(n_275), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_189), .A2(n_608), .B(n_609), .Y(n_607) );
INVx1_ASAP7_75t_L g291 ( .A(n_192), .Y(n_291) );
INVx1_ASAP7_75t_L g296 ( .A(n_192), .Y(n_296) );
INVx1_ASAP7_75t_L g340 ( .A(n_192), .Y(n_340) );
AND2x2_ASAP7_75t_L g518 ( .A(n_192), .B(n_427), .Y(n_518) );
OAI21x1_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_208), .Y(n_192) );
OAI21x1_ASAP7_75t_L g671 ( .A1(n_193), .A2(n_672), .B(n_682), .Y(n_671) );
OAI21x1_ASAP7_75t_L g693 ( .A1(n_193), .A2(n_694), .B(n_703), .Y(n_693) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_198), .B(n_200), .Y(n_195) );
INVx2_ASAP7_75t_L g593 ( .A(n_197), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_197), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g597 ( .A(n_199), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_200), .A2(n_260), .B(n_262), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_204), .B(n_206), .Y(n_201) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_207), .B(n_678), .Y(n_677) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_209), .Y(n_619) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_213), .B(n_233), .Y(n_212) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g361 ( .A(n_214), .B(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g367 ( .A(n_214), .B(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_214), .B(n_353), .Y(n_388) );
AND2x2_ASAP7_75t_L g412 ( .A(n_214), .B(n_298), .Y(n_412) );
BUFx3_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
OR2x2_ASAP7_75t_L g335 ( .A(n_215), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g489 ( .A(n_215), .B(n_433), .Y(n_489) );
AND2x2_ASAP7_75t_L g495 ( .A(n_215), .B(n_314), .Y(n_495) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g287 ( .A(n_216), .Y(n_287) );
AND2x2_ASAP7_75t_L g307 ( .A(n_216), .B(n_285), .Y(n_307) );
INVx2_ASAP7_75t_L g344 ( .A(n_216), .Y(n_344) );
INVx1_ASAP7_75t_L g376 ( .A(n_216), .Y(n_376) );
AND2x2_ASAP7_75t_L g383 ( .A(n_216), .B(n_336), .Y(n_383) );
AND2x2_ASAP7_75t_L g419 ( .A(n_216), .B(n_375), .Y(n_419) );
BUFx2_ASAP7_75t_L g458 ( .A(n_216), .Y(n_458) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_216), .Y(n_481) );
OR2x6_ASAP7_75t_L g216 ( .A(n_217), .B(n_221), .Y(n_216) );
INVxp67_ASAP7_75t_SL g218 ( .A(n_219), .Y(n_218) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_219), .Y(n_238) );
NOR2xp67_ASAP7_75t_SL g251 ( .A(n_219), .B(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g710 ( .A(n_219), .Y(n_710) );
OAI21xp5_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_227), .Y(n_222) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g245 ( .A(n_225), .Y(n_245) );
INVx2_ASAP7_75t_L g276 ( .A(n_225), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_225), .B(n_319), .Y(n_318) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_225), .Y(n_575) );
INVx3_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_226), .Y(n_255) );
INVx2_ASAP7_75t_L g580 ( .A(n_230), .Y(n_580) );
INVxp67_ASAP7_75t_L g643 ( .A(n_232), .Y(n_643) );
INVxp67_ASAP7_75t_L g674 ( .A(n_232), .Y(n_674) );
AOI22xp33_ASAP7_75t_SL g399 ( .A1(n_233), .A2(n_337), .B1(n_378), .B2(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
OR2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_264), .Y(n_234) );
INVx4_ASAP7_75t_L g298 ( .A(n_235), .Y(n_298) );
NAND2xp33_ASAP7_75t_SL g351 ( .A(n_235), .B(n_352), .Y(n_351) );
OAI32xp33_ASAP7_75t_L g496 ( .A1(n_235), .A2(n_381), .A3(n_497), .B1(n_498), .B2(n_500), .Y(n_496) );
OR2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_249), .Y(n_235) );
INVx2_ASAP7_75t_L g348 ( .A(n_236), .Y(n_348) );
OAI21x1_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_239), .B(n_248), .Y(n_236) );
OAI21x1_ASAP7_75t_L g266 ( .A1(n_237), .A2(n_267), .B(n_279), .Y(n_266) );
OAI21xp5_ASAP7_75t_L g285 ( .A1(n_237), .A2(n_239), .B(n_248), .Y(n_285) );
OAI21x1_ASAP7_75t_L g605 ( .A1(n_237), .A2(n_606), .B(n_614), .Y(n_605) );
OAI21x1_ASAP7_75t_L g714 ( .A1(n_237), .A2(n_635), .B(n_715), .Y(n_714) );
OAI21x1_ASAP7_75t_L g740 ( .A1(n_237), .A2(n_606), .B(n_614), .Y(n_740) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NOR2x1_ASAP7_75t_SL g599 ( .A(n_238), .B(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g640 ( .A(n_245), .Y(n_640) );
AND2x4_ASAP7_75t_L g286 ( .A(n_249), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g306 ( .A(n_249), .Y(n_306) );
INVx2_ASAP7_75t_L g336 ( .A(n_249), .Y(n_336) );
AND2x2_ASAP7_75t_L g362 ( .A(n_249), .B(n_348), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_249), .B(n_265), .Y(n_368) );
AND2x4_ASAP7_75t_L g249 ( .A(n_250), .B(n_258), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_253), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_251), .A2(n_259), .B(n_263), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_256), .B(n_257), .Y(n_253) );
INVx1_ASAP7_75t_L g317 ( .A(n_255), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_255), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g613 ( .A(n_255), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_255), .B(n_656), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g595 ( .A1(n_257), .A2(n_596), .B(n_598), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_261), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g450 ( .A(n_264), .B(n_383), .Y(n_450) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_264), .Y(n_499) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_265), .Y(n_310) );
AND2x2_ASAP7_75t_L g353 ( .A(n_265), .B(n_348), .Y(n_353) );
AND2x2_ASAP7_75t_L g432 ( .A(n_265), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g302 ( .A(n_266), .Y(n_302) );
INVx1_ASAP7_75t_L g347 ( .A(n_266), .Y(n_347) );
OAI21xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_272), .B(n_277), .Y(n_267) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx2_ASAP7_75t_SL g321 ( .A(n_278), .Y(n_321) );
INVx1_ASAP7_75t_L g629 ( .A(n_278), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_288), .B1(n_292), .B2(n_297), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_286), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_283), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g478 ( .A(n_283), .Y(n_478) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g385 ( .A(n_284), .B(n_301), .Y(n_385) );
OAI22xp33_ASAP7_75t_L g504 ( .A1(n_284), .A2(n_391), .B1(n_471), .B2(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g443 ( .A(n_285), .B(n_336), .Y(n_443) );
AND2x2_ASAP7_75t_L g406 ( .A(n_286), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g428 ( .A(n_286), .B(n_429), .Y(n_428) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_286), .Y(n_487) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_287), .Y(n_474) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_289), .Y(n_370) );
AND2x2_ASAP7_75t_L g425 ( .A(n_289), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g435 ( .A(n_289), .B(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g475 ( .A(n_289), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_289), .B(n_476), .Y(n_491) );
AND2x2_ASAP7_75t_L g330 ( .A(n_290), .B(n_331), .Y(n_330) );
INVx3_ASAP7_75t_L g454 ( .A(n_290), .Y(n_454) );
AOI33xp33_ASAP7_75t_L g488 ( .A1(n_290), .A2(n_298), .A3(n_371), .B1(n_489), .B2(n_490), .B3(n_495), .Y(n_488) );
NAND2x1p5_ASAP7_75t_L g311 ( .A(n_292), .B(n_312), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g350 ( .A1(n_292), .A2(n_351), .B1(n_354), .B2(n_361), .Y(n_350) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
AND2x2_ASAP7_75t_L g449 ( .A(n_293), .B(n_426), .Y(n_449) );
AND2x4_ASAP7_75t_L g517 ( .A(n_293), .B(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g379 ( .A(n_294), .B(n_314), .Y(n_379) );
INVx1_ASAP7_75t_L g476 ( .A(n_294), .Y(n_476) );
BUFx3_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVxp67_ASAP7_75t_SL g357 ( .A(n_296), .Y(n_357) );
NOR2x1_ASAP7_75t_L g395 ( .A(n_297), .B(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g472 ( .A(n_297), .Y(n_472) );
AND2x4_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
OAI21xp33_ASAP7_75t_L g515 ( .A1(n_298), .A2(n_479), .B(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g334 ( .A(n_300), .B(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g397 ( .A(n_300), .B(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_300), .B(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g375 ( .A(n_302), .Y(n_375) );
A2O1A1Ixp33_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_308), .B(n_311), .C(n_329), .Y(n_303) );
NAND2x1_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_305), .A2(n_513), .B1(n_515), .B2(n_519), .Y(n_512) );
INVx4_ASAP7_75t_R g305 ( .A(n_306), .Y(n_305) );
OAI32xp33_ASAP7_75t_L g477 ( .A1(n_306), .A2(n_478), .A3(n_479), .B1(n_480), .B2(n_482), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_306), .B(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g309 ( .A(n_307), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g479 ( .A(n_312), .B(n_454), .Y(n_479) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_314), .Y(n_338) );
BUFx2_ASAP7_75t_L g372 ( .A(n_314), .Y(n_372) );
INVx1_ASAP7_75t_L g394 ( .A(n_314), .Y(n_394) );
NAND2x1p5_ASAP7_75t_L g314 ( .A(n_315), .B(n_324), .Y(n_314) );
NAND2x1p5_ASAP7_75t_L g332 ( .A(n_315), .B(n_324), .Y(n_332) );
OA21x2_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_320), .B(n_322), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_317), .A2(n_593), .B1(n_663), .B2(n_665), .Y(n_662) );
OR2x2_ASAP7_75t_L g324 ( .A(n_320), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g600 ( .A(n_321), .Y(n_600) );
INVxp67_ASAP7_75t_L g646 ( .A(n_323), .Y(n_646) );
INVx1_ASAP7_75t_L g576 ( .A(n_328), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g591 ( .A1(n_328), .A2(n_592), .B(n_594), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_333), .B1(n_337), .B2(n_341), .Y(n_329) );
AOI222xp33_ASAP7_75t_L g421 ( .A1(n_330), .A2(n_422), .B1(n_428), .B2(n_430), .C1(n_435), .C2(n_437), .Y(n_421) );
AND2x2_ASAP7_75t_L g364 ( .A(n_331), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g359 ( .A(n_332), .B(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g427 ( .A(n_332), .Y(n_427) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OAI22xp33_ASAP7_75t_L g413 ( .A1(n_334), .A2(n_414), .B1(n_418), .B2(n_420), .Y(n_413) );
INVx2_ASAP7_75t_L g434 ( .A(n_335), .Y(n_434) );
AND2x4_ASAP7_75t_SL g343 ( .A(n_336), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
AND2x4_ASAP7_75t_SL g386 ( .A(n_339), .B(n_379), .Y(n_386) );
INVx1_ASAP7_75t_L g471 ( .A(n_339), .Y(n_471) );
AND2x2_ASAP7_75t_L g426 ( .A(n_340), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
INVx1_ASAP7_75t_L g398 ( .A(n_343), .Y(n_398) );
INVx1_ASAP7_75t_L g438 ( .A(n_343), .Y(n_438) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_SL g407 ( .A(n_346), .Y(n_407) );
INVx1_ASAP7_75t_L g463 ( .A(n_346), .Y(n_463) );
OR2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
BUFx2_ASAP7_75t_L g493 ( .A(n_347), .Y(n_493) );
INVx1_ASAP7_75t_L g433 ( .A(n_348), .Y(n_433) );
NAND3xp33_ASAP7_75t_L g349 ( .A(n_350), .B(n_363), .C(n_377), .Y(n_349) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_353), .B(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
OR2x2_ASAP7_75t_L g453 ( .A(n_358), .B(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g466 ( .A(n_359), .B(n_365), .Y(n_466) );
INVx1_ASAP7_75t_L g392 ( .A(n_360), .Y(n_392) );
AND2x2_ASAP7_75t_L g373 ( .A(n_362), .B(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_362), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g464 ( .A(n_362), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_366), .B1(n_369), .B2(n_373), .Y(n_363) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g402 ( .A(n_368), .Y(n_402) );
OAI22xp33_ASAP7_75t_L g490 ( .A1(n_368), .A2(n_491), .B1(n_492), .B2(n_494), .Y(n_490) );
AND2x4_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_375), .Y(n_429) );
OR2x2_ASAP7_75t_L g514 ( .A(n_375), .B(n_376), .Y(n_514) );
AOI32xp33_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_381), .A3(n_384), .B1(n_386), .B2(n_387), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
INVx2_ASAP7_75t_L g409 ( .A(n_380), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_380), .B(n_393), .Y(n_497) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND3xp33_ASAP7_75t_SL g508 ( .A(n_384), .B(n_464), .C(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g461 ( .A(n_386), .Y(n_461) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OAI21xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_395), .B(n_399), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_393), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_397), .A2(n_470), .B1(n_472), .B2(n_473), .Y(n_469) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_404), .B(n_467), .Y(n_403) );
NAND4xp25_ASAP7_75t_L g404 ( .A(n_405), .B(n_421), .C(n_439), .D(n_451), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_408), .B1(n_410), .B2(n_412), .C(n_413), .Y(n_405) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g511 ( .A(n_409), .B(n_417), .Y(n_511) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_417), .Y(n_414) );
OR2x2_ASAP7_75t_L g500 ( .A(n_415), .B(n_454), .Y(n_500) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g436 ( .A(n_417), .Y(n_436) );
OR2x2_ASAP7_75t_L g470 ( .A(n_417), .B(n_471), .Y(n_470) );
OR2x2_ASAP7_75t_L g507 ( .A(n_417), .B(n_481), .Y(n_507) );
INVx1_ASAP7_75t_L g440 ( .A(n_418), .Y(n_440) );
INVxp67_ASAP7_75t_SL g502 ( .A(n_420), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g519 ( .A(n_425), .B(n_476), .Y(n_519) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_434), .Y(n_431) );
INVx1_ASAP7_75t_L g505 ( .A(n_432), .Y(n_505) );
OAI32xp33_ASAP7_75t_L g460 ( .A1(n_437), .A2(n_461), .A3(n_462), .B1(n_464), .B2(n_465), .Y(n_460) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
O2A1O1Ixp33_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_441), .B(n_444), .C(n_448), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g459 ( .A(n_443), .Y(n_459) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
AND2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
INVx1_ASAP7_75t_L g509 ( .A(n_450), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_455), .B(n_460), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_459), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NAND4xp25_ASAP7_75t_L g467 ( .A(n_468), .B(n_484), .C(n_501), .D(n_512), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_477), .Y(n_468) );
NAND3xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .C(n_476), .Y(n_473) );
AOI322xp5_ASAP7_75t_L g501 ( .A1(n_478), .A2(n_502), .A3(n_503), .B1(n_504), .B2(n_506), .C1(n_508), .C2(n_510), .Y(n_501) );
OAI21xp33_ASAP7_75t_L g485 ( .A1(n_479), .A2(n_486), .B(n_488), .Y(n_485) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_481), .Y(n_503) );
INVx2_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
NOR2xp33_ASAP7_75t_SL g484 ( .A(n_485), .B(n_496), .Y(n_484) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_521), .Y(n_520) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_SL g536 ( .A(n_526), .Y(n_536) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_527), .Y(n_539) );
INVx2_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
NOR2x1p5_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_531), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
OAI21xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_546), .B(n_933), .Y(n_540) );
BUFx8_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
OR2x6_ASAP7_75t_L g542 ( .A(n_543), .B(n_545), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_553), .B1(n_554), .B2(n_932), .Y(n_546) );
INVx1_ASAP7_75t_L g932 ( .A(n_547), .Y(n_932) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVxp67_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
BUFx8_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
BUFx6f_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND3x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_836), .C(n_882), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_562), .B(n_780), .Y(n_561) );
NAND3xp33_ASAP7_75t_SL g562 ( .A(n_563), .B(n_717), .C(n_752), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_601), .B1(n_704), .B2(n_711), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_586), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x4_ASAP7_75t_L g832 ( .A(n_567), .B(n_604), .Y(n_832) );
AND2x4_ASAP7_75t_L g845 ( .A(n_567), .B(n_740), .Y(n_845) );
AND2x2_ASAP7_75t_L g876 ( .A(n_567), .B(n_761), .Y(n_876) );
HB1xp67_ASAP7_75t_L g909 ( .A(n_567), .Y(n_909) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OR2x6_ASAP7_75t_L g729 ( .A(n_568), .B(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_SL g741 ( .A(n_568), .B(n_708), .Y(n_741) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g707 ( .A(n_569), .Y(n_707) );
OAI21x1_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_577), .B(n_585), .Y(n_569) );
AOI21x1_ASAP7_75t_SL g570 ( .A1(n_571), .A2(n_574), .B(n_576), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
AOI22x1_ASAP7_75t_L g635 ( .A1(n_576), .A2(n_584), .B1(n_636), .B2(n_642), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_580), .A2(n_643), .B1(n_644), .B2(n_645), .Y(n_642) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AOI21x1_ASAP7_75t_L g621 ( .A1(n_584), .A2(n_622), .B(n_623), .Y(n_621) );
OR2x2_ASAP7_75t_L g821 ( .A(n_586), .B(n_822), .Y(n_821) );
OR2x2_ASAP7_75t_L g842 ( .A(n_586), .B(n_729), .Y(n_842) );
BUFx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g749 ( .A(n_587), .Y(n_749) );
AND2x2_ASAP7_75t_L g756 ( .A(n_587), .B(n_708), .Y(n_756) );
INVx2_ASAP7_75t_L g761 ( .A(n_587), .Y(n_761) );
AND2x2_ASAP7_75t_L g776 ( .A(n_587), .B(n_777), .Y(n_776) );
AND2x4_ASAP7_75t_L g786 ( .A(n_587), .B(n_616), .Y(n_786) );
OR2x2_ASAP7_75t_L g802 ( .A(n_587), .B(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g831 ( .A(n_587), .Y(n_831) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND2x1_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
OAI21x1_ASAP7_75t_SL g590 ( .A1(n_591), .A2(n_595), .B(n_599), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_631), .B1(n_683), .B2(n_687), .Y(n_601) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g869 ( .A(n_603), .B(n_870), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_615), .Y(n_603) );
BUFx3_ASAP7_75t_L g685 ( .A(n_604), .Y(n_685) );
AND2x2_ASAP7_75t_L g774 ( .A(n_604), .B(n_749), .Y(n_774) );
INVx1_ASAP7_75t_L g777 ( .A(n_604), .Y(n_777) );
AND2x2_ASAP7_75t_L g891 ( .A(n_604), .B(n_707), .Y(n_891) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
HB1xp67_ASAP7_75t_L g813 ( .A(n_605), .Y(n_813) );
INVxp67_ASAP7_75t_L g627 ( .A(n_613), .Y(n_627) );
HB1xp67_ASAP7_75t_L g789 ( .A(n_615), .Y(n_789) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_616), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_616), .B(n_707), .Y(n_822) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g730 ( .A(n_617), .Y(n_730) );
INVxp67_ASAP7_75t_SL g803 ( .A(n_617), .Y(n_803) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI21x1_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_620), .B(n_630), .Y(n_618) );
OA21x2_ASAP7_75t_L g708 ( .A1(n_620), .A2(n_630), .B(n_709), .Y(n_708) );
OAI21x1_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_624), .B(n_629), .Y(n_620) );
OAI21xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_627), .B(n_628), .Y(n_624) );
OAI21xp5_ASAP7_75t_L g694 ( .A1(n_629), .A2(n_695), .B(n_698), .Y(n_694) );
INVx2_ASAP7_75t_L g782 ( .A(n_631), .Y(n_782) );
OR2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_649), .Y(n_631) );
INVx1_ASAP7_75t_L g747 ( .A(n_632), .Y(n_747) );
INVx1_ASAP7_75t_L g779 ( .A(n_632), .Y(n_779) );
BUFx3_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g765 ( .A(n_633), .Y(n_765) );
AO31x2_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_646), .A3(n_647), .B(n_648), .Y(n_633) );
AO31x2_ASAP7_75t_L g797 ( .A1(n_634), .A2(n_646), .A3(n_647), .B(n_648), .Y(n_797) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OAI22x1_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_639), .B1(n_640), .B2(n_641), .Y(n_636) );
INVxp67_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g715 ( .A(n_648), .Y(n_715) );
INVx1_ASAP7_75t_L g915 ( .A(n_649), .Y(n_915) );
INVxp67_ASAP7_75t_SL g926 ( .A(n_649), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_669), .Y(n_649) );
NOR2x1_ASAP7_75t_L g690 ( .A(n_650), .B(n_691), .Y(n_690) );
BUFx2_ASAP7_75t_L g751 ( .A(n_650), .Y(n_751) );
INVx1_ASAP7_75t_L g793 ( .A(n_650), .Y(n_793) );
AND2x2_ASAP7_75t_L g852 ( .A(n_650), .B(n_670), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_650), .B(n_716), .Y(n_874) );
INVx3_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g712 ( .A(n_651), .B(n_670), .Y(n_712) );
AO21x2_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B(n_667), .Y(n_651) );
AO21x1_ASAP7_75t_L g725 ( .A1(n_652), .A2(n_653), .B(n_667), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_662), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_657), .B1(n_659), .B2(n_661), .Y(n_654) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_670), .Y(n_689) );
INVx3_ASAP7_75t_L g721 ( .A(n_670), .Y(n_721) );
INVx2_ASAP7_75t_L g734 ( .A(n_670), .Y(n_734) );
AND2x2_ASAP7_75t_L g738 ( .A(n_670), .B(n_714), .Y(n_738) );
INVx1_ASAP7_75t_L g762 ( .A(n_670), .Y(n_762) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OAI21xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_675), .B(n_676), .Y(n_673) );
INVxp67_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_685), .B(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g800 ( .A(n_685), .Y(n_800) );
OR2x2_ASAP7_75t_L g841 ( .A(n_685), .B(n_842), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_690), .Y(n_687) );
OR2x2_ASAP7_75t_L g921 ( .A(n_688), .B(n_922), .Y(n_921) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g737 ( .A(n_691), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_691), .B(n_721), .Y(n_770) );
NOR2xp67_ASAP7_75t_L g880 ( .A(n_691), .B(n_720), .Y(n_880) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx3_ASAP7_75t_L g716 ( .A(n_692), .Y(n_716) );
AND2x2_ASAP7_75t_L g723 ( .A(n_692), .B(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g835 ( .A(n_692), .B(n_714), .Y(n_835) );
INVx1_ASAP7_75t_L g858 ( .A(n_692), .Y(n_858) );
INVx3_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AOI211xp5_ASAP7_75t_L g717 ( .A1(n_706), .A2(n_718), .B(n_726), .C(n_742), .Y(n_717) );
AND2x2_ASAP7_75t_L g866 ( .A(n_706), .B(n_830), .Y(n_866) );
NAND2xp5_ASAP7_75t_SL g919 ( .A(n_706), .B(n_761), .Y(n_919) );
AND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
INVx1_ASAP7_75t_L g745 ( .A(n_707), .Y(n_745) );
AND2x4_ASAP7_75t_L g755 ( .A(n_707), .B(n_740), .Y(n_755) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
AOI32xp33_ASAP7_75t_L g843 ( .A1(n_711), .A2(n_785), .A3(n_844), .B1(n_846), .B2(n_848), .Y(n_843) );
AND2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
AND2x2_ASAP7_75t_L g834 ( .A(n_712), .B(n_835), .Y(n_834) );
INVx2_ASAP7_75t_L g735 ( .A(n_713), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_713), .B(n_793), .Y(n_809) );
AND2x2_ASAP7_75t_L g862 ( .A(n_713), .B(n_751), .Y(n_862) );
AND2x2_ASAP7_75t_L g925 ( .A(n_713), .B(n_926), .Y(n_925) );
AND2x4_ASAP7_75t_L g713 ( .A(n_714), .B(n_716), .Y(n_713) );
INVx1_ASAP7_75t_L g772 ( .A(n_714), .Y(n_772) );
OR2x2_ASAP7_75t_L g796 ( .A(n_716), .B(n_797), .Y(n_796) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
AOI21xp33_ASAP7_75t_SL g815 ( .A1(n_719), .A2(n_773), .B(n_814), .Y(n_815) );
OR2x2_ASAP7_75t_L g719 ( .A(n_720), .B(n_722), .Y(n_719) );
BUFx2_ASAP7_75t_L g860 ( .A(n_720), .Y(n_860) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_721), .B(n_779), .Y(n_778) );
OR2x2_ASAP7_75t_L g825 ( .A(n_721), .B(n_797), .Y(n_825) );
INVx1_ASAP7_75t_L g759 ( .A(n_722), .Y(n_759) );
OR2x2_ASAP7_75t_L g805 ( .A(n_722), .B(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g764 ( .A(n_723), .Y(n_764) );
HB1xp67_ASAP7_75t_L g826 ( .A(n_723), .Y(n_826) );
AND2x2_ASAP7_75t_L g867 ( .A(n_723), .B(n_765), .Y(n_867) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g733 ( .A(n_725), .B(n_734), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_725), .B(n_772), .Y(n_771) );
OAI22xp33_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_731), .B1(n_736), .B2(n_739), .Y(n_726) );
INVxp67_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NAND2x1p5_ASAP7_75t_L g775 ( .A(n_728), .B(n_776), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_728), .A2(n_898), .B1(n_900), .B2(n_902), .Y(n_897) );
INVx2_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
OR2x2_ASAP7_75t_L g818 ( .A(n_729), .B(n_761), .Y(n_818) );
AND2x2_ASAP7_75t_L g746 ( .A(n_730), .B(n_740), .Y(n_746) );
INVx2_ASAP7_75t_L g931 ( .A(n_731), .Y(n_931) );
OR2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_735), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g839 ( .A(n_733), .B(n_840), .Y(n_839) );
AND2x2_ASAP7_75t_L g848 ( .A(n_733), .B(n_835), .Y(n_848) );
AND2x2_ASAP7_75t_L g887 ( .A(n_733), .B(n_779), .Y(n_887) );
AND2x2_ASAP7_75t_L g906 ( .A(n_733), .B(n_870), .Y(n_906) );
INVx1_ASAP7_75t_L g753 ( .A(n_735), .Y(n_753) );
OAI321xp33_ASAP7_75t_L g923 ( .A1(n_736), .A2(n_812), .A3(n_846), .B1(n_924), .B2(n_927), .C(n_930), .Y(n_923) );
NAND2xp5_ASAP7_75t_SL g736 ( .A(n_737), .B(n_738), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_737), .B(n_879), .Y(n_922) );
INVx1_ASAP7_75t_L g806 ( .A(n_738), .Y(n_806) );
AND2x4_ASAP7_75t_L g872 ( .A(n_738), .B(n_873), .Y(n_872) );
INVx3_ASAP7_75t_L g893 ( .A(n_739), .Y(n_893) );
OR2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
AND2x4_ASAP7_75t_L g785 ( .A(n_740), .B(n_786), .Y(n_785) );
INVx2_ASAP7_75t_L g767 ( .A(n_741), .Y(n_767) );
NOR4xp25_ASAP7_75t_L g742 ( .A(n_743), .B(n_747), .C(n_748), .D(n_750), .Y(n_742) );
NAND2x1_ASAP7_75t_L g783 ( .A(n_743), .B(n_784), .Y(n_783) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g865 ( .A1(n_744), .A2(n_819), .B1(n_866), .B2(n_867), .Y(n_865) );
AND2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
OAI322xp33_ASAP7_75t_L g904 ( .A1(n_747), .A2(n_905), .A3(n_907), .B1(n_913), .B2(n_916), .C1(n_917), .C2(n_921), .Y(n_904) );
AND2x2_ASAP7_75t_L g864 ( .A(n_748), .B(n_832), .Y(n_864) );
BUFx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
AND2x2_ASAP7_75t_L g847 ( .A(n_749), .B(n_803), .Y(n_847) );
INVx1_ASAP7_75t_L g870 ( .A(n_749), .Y(n_870) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
NOR2x1_ASAP7_75t_L g819 ( .A(n_751), .B(n_796), .Y(n_819) );
AOI211xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_754), .B(n_757), .C(n_768), .Y(n_752) );
AND2x2_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
INVx1_ASAP7_75t_L g828 ( .A(n_755), .Y(n_828) );
NOR2x1_ASAP7_75t_L g928 ( .A(n_755), .B(n_929), .Y(n_928) );
INVx2_ASAP7_75t_L g814 ( .A(n_756), .Y(n_814) );
O2A1O1Ixp33_ASAP7_75t_SL g757 ( .A1(n_758), .A2(n_760), .B(n_763), .C(n_766), .Y(n_757) );
INVxp67_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
OR2x2_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
AND2x2_ASAP7_75t_L g920 ( .A(n_761), .B(n_891), .Y(n_920) );
INVx2_ASAP7_75t_L g795 ( .A(n_762), .Y(n_795) );
OR2x6_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
INVx2_ASAP7_75t_L g840 ( .A(n_765), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_765), .B(n_852), .Y(n_851) );
NAND2xp33_ASAP7_75t_SL g902 ( .A(n_766), .B(n_903), .Y(n_902) );
INVx2_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
OAI32xp33_ASAP7_75t_L g768 ( .A1(n_767), .A2(n_769), .A3(n_773), .B1(n_775), .B2(n_778), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_767), .B(n_870), .Y(n_916) );
OR2x2_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
INVx2_ASAP7_75t_L g879 ( .A(n_771), .Y(n_879) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
OR2x2_ASAP7_75t_L g850 ( .A(n_777), .B(n_822), .Y(n_850) );
NAND3xp33_ASAP7_75t_L g780 ( .A(n_781), .B(n_798), .C(n_816), .Y(n_780) );
AOI22xp5_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_783), .B1(n_787), .B2(n_790), .Y(n_781) );
INVx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
O2A1O1Ixp5_ASAP7_75t_L g827 ( .A1(n_786), .A2(n_828), .B(n_829), .C(n_833), .Y(n_827) );
HB1xp67_ASAP7_75t_L g885 ( .A(n_786), .Y(n_885) );
INVx1_ASAP7_75t_L g929 ( .A(n_786), .Y(n_929) );
INVxp67_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVxp67_ASAP7_75t_SL g788 ( .A(n_789), .Y(n_788) );
INVx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_792), .B(n_794), .Y(n_791) );
INVx1_ASAP7_75t_L g896 ( .A(n_792), .Y(n_896) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
AND2x2_ASAP7_75t_L g901 ( .A(n_793), .B(n_858), .Y(n_901) );
INVx1_ASAP7_75t_L g808 ( .A(n_794), .Y(n_808) );
NOR2x1p5_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .Y(n_794) );
INVx1_ASAP7_75t_L g859 ( .A(n_797), .Y(n_859) );
AOI221xp5_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_804), .B1(n_807), .B2(n_810), .C(n_815), .Y(n_798) );
INVx1_ASAP7_75t_L g854 ( .A(n_799), .Y(n_854) );
AND2x2_ASAP7_75t_L g799 ( .A(n_800), .B(n_801), .Y(n_799) );
INVx2_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
OR2x2_ASAP7_75t_L g889 ( .A(n_802), .B(n_890), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_804), .B(n_885), .Y(n_884) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .Y(n_807) );
INVx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
OR2x2_ASAP7_75t_L g811 ( .A(n_812), .B(n_814), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
AND2x2_ASAP7_75t_L g881 ( .A(n_813), .B(n_847), .Y(n_881) );
AOI221xp5_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_819), .B1(n_820), .B2(n_823), .C(n_827), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
AND2x2_ASAP7_75t_L g823 ( .A(n_824), .B(n_826), .Y(n_823) );
AND2x4_ASAP7_75t_L g900 ( .A(n_824), .B(n_901), .Y(n_900) );
INVx2_ASAP7_75t_SL g824 ( .A(n_825), .Y(n_824) );
OR2x2_ASAP7_75t_L g899 ( .A(n_825), .B(n_874), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_830), .B(n_832), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx3_ASAP7_75t_R g903 ( .A(n_832), .Y(n_903) );
INVx2_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
NOR4xp25_ASAP7_75t_L g836 ( .A(n_837), .B(n_849), .C(n_853), .D(n_868), .Y(n_836) );
OAI21xp33_ASAP7_75t_SL g837 ( .A1(n_838), .A2(n_841), .B(n_843), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
AOI21xp33_ASAP7_75t_SL g849 ( .A1(n_841), .A2(n_850), .B(n_851), .Y(n_849) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
OAI21xp5_ASAP7_75t_L g930 ( .A1(n_845), .A2(n_881), .B(n_931), .Y(n_930) );
BUFx3_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
OAI221xp5_ASAP7_75t_SL g853 ( .A1(n_854), .A2(n_855), .B1(n_861), .B2(n_863), .C(n_865), .Y(n_853) );
OAI221xp5_ASAP7_75t_L g868 ( .A1(n_855), .A2(n_869), .B1(n_871), .B2(n_875), .C(n_877), .Y(n_868) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
AND2x2_ASAP7_75t_L g856 ( .A(n_857), .B(n_860), .Y(n_856) );
INVx1_ASAP7_75t_L g895 ( .A(n_857), .Y(n_895) );
AND2x4_ASAP7_75t_L g914 ( .A(n_857), .B(n_915), .Y(n_914) );
AND2x2_ASAP7_75t_L g857 ( .A(n_858), .B(n_859), .Y(n_857) );
INVx1_ASAP7_75t_L g911 ( .A(n_858), .Y(n_911) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVxp67_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
NAND4xp25_ASAP7_75t_L g892 ( .A(n_870), .B(n_893), .C(n_894), .D(n_896), .Y(n_892) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVxp67_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_878), .B(n_881), .Y(n_877) );
AND2x2_ASAP7_75t_L g878 ( .A(n_879), .B(n_880), .Y(n_878) );
NOR3xp33_ASAP7_75t_L g882 ( .A(n_883), .B(n_904), .C(n_923), .Y(n_882) );
NAND4xp25_ASAP7_75t_L g883 ( .A(n_884), .B(n_886), .C(n_892), .D(n_897), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_887), .B(n_888), .Y(n_886) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
HB1xp67_ASAP7_75t_L g912 ( .A(n_891), .Y(n_912) );
INVx1_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
INVx1_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
NOR2xp33_ASAP7_75t_SL g907 ( .A(n_908), .B(n_912), .Y(n_907) );
NOR2xp33_ASAP7_75t_L g908 ( .A(n_909), .B(n_910), .Y(n_908) );
INVx2_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
NOR2xp33_ASAP7_75t_L g917 ( .A(n_918), .B(n_920), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
BUFx6f_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
NOR2xp33_ASAP7_75t_R g938 ( .A(n_939), .B(n_940), .Y(n_938) );
endmodule