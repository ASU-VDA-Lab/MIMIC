module fake_jpeg_7149_n_138 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_138);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_138;

wire n_117;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_1),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_23),
.B(n_25),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_13),
.Y(n_31)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g28 ( 
.A(n_16),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_34),
.Y(n_46)
);

AND2x2_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_13),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_21),
.A2(n_17),
.B1(n_11),
.B2(n_20),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_19),
.B1(n_10),
.B2(n_17),
.Y(n_41)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_35),
.B(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_39),
.B(n_44),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_22),
.B(n_28),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_49),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_35),
.B(n_23),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVxp33_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_48),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_47),
.B(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_22),
.B1(n_21),
.B2(n_25),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_40),
.B1(n_38),
.B2(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_46),
.B(n_31),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_46),
.B(n_19),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_10),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_32),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_24),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_63),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_24),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_68),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_67),
.B1(n_61),
.B2(n_63),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_48),
.B1(n_47),
.B2(n_36),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

NOR4xp25_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_47),
.C(n_27),
.D(n_29),
.Y(n_69)
);

NAND3xp33_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_68),
.C(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_73),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_75),
.Y(n_87)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_30),
.Y(n_74)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_24),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_30),
.Y(n_76)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

OAI221xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_86),
.B1(n_24),
.B2(n_30),
.C(n_32),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_73),
.A2(n_61),
.B(n_52),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_81),
.B(n_12),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_52),
.B(n_27),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_30),
.B1(n_36),
.B2(n_29),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_36),
.B1(n_26),
.B2(n_12),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_36),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_25),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_26),
.C(n_30),
.Y(n_91)
);

OA21x2_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_69),
.B(n_71),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_93),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_94),
.C(n_101),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_96),
.B(n_100),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_79),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_95),
.A2(n_99),
.B1(n_83),
.B2(n_87),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_32),
.Y(n_96)
);

OAI322xp33_ASAP7_75t_L g97 ( 
.A1(n_77),
.A2(n_24),
.A3(n_33),
.B1(n_32),
.B2(n_15),
.C1(n_14),
.C2(n_20),
.Y(n_97)
);

NOR3xp33_ASAP7_75t_SL g106 ( 
.A(n_97),
.B(n_14),
.C(n_33),
.Y(n_106)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_33),
.C(n_32),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_102),
.A2(n_104),
.B1(n_105),
.B2(n_95),
.Y(n_115)
);

OAI21x1_ASAP7_75t_L g104 ( 
.A1(n_99),
.A2(n_82),
.B(n_85),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_14),
.B1(n_15),
.B2(n_33),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_108),
.Y(n_114)
);

NOR3xp33_ASAP7_75t_SL g108 ( 
.A(n_90),
.B(n_5),
.C(n_8),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_1),
.C(n_2),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_5),
.C(n_8),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_101),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_106),
.Y(n_120)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_109),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_115),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_107),
.A2(n_98),
.B1(n_90),
.B2(n_91),
.Y(n_113)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_117),
.Y(n_123)
);

BUFx24_ASAP7_75t_SL g117 ( 
.A(n_108),
.Y(n_117)
);

FAx1_ASAP7_75t_SL g119 ( 
.A(n_113),
.B(n_110),
.CI(n_103),
.CON(n_119),
.SN(n_119)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_114),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_121),
.C(n_116),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_5),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_118),
.A2(n_122),
.B(n_119),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_124),
.A2(n_128),
.B(n_9),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_127),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_126),
.A2(n_121),
.B(n_120),
.Y(n_129)
);

AOI31xp33_ASAP7_75t_SL g127 ( 
.A1(n_119),
.A2(n_4),
.A3(n_6),
.B(n_7),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_7),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_132),
.C(n_9),
.Y(n_133)
);

NOR3xp33_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_1),
.C(n_2),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_9),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_135),
.C(n_3),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_2),
.B(n_3),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_2),
.C(n_3),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_137),
.Y(n_138)
);


endmodule