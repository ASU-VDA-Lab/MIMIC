module fake_netlist_5_893_n_1121 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1121);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1121;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_419;
wire n_380;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_316;
wire n_785;
wire n_389;
wire n_855;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_968;
wire n_912;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_718;
wire n_671;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_1120;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_859;
wire n_864;
wire n_1110;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_946;
wire n_417;
wire n_932;
wire n_1048;
wire n_612;
wire n_1001;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_509;
wire n_568;
wire n_936;
wire n_373;
wire n_820;
wire n_947;
wire n_757;
wire n_1090;
wire n_307;
wire n_633;
wire n_530;
wire n_439;
wire n_1024;
wire n_1063;
wire n_556;
wire n_1107;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1032;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_1104;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_992;
wire n_1049;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_519;
wire n_406;
wire n_470;
wire n_919;
wire n_782;
wire n_908;
wire n_1108;
wire n_325;
wire n_449;
wire n_1073;
wire n_1100;
wire n_862;
wire n_900;
wire n_1016;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_976;
wire n_1096;
wire n_1095;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_660;
wire n_223;
wire n_1114;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_696;
wire n_255;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_1062;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_974;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_1119;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_829;
wire n_928;
wire n_749;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_342;
wire n_517;
wire n_482;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_1069;
wire n_236;
wire n_1075;
wire n_388;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_1113;
wire n_652;
wire n_778;
wire n_1111;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_201;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_781;
wire n_711;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_1015;
wire n_1000;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_846;
wire n_586;
wire n_748;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_332;
wire n_1101;
wire n_1053;
wire n_273;
wire n_585;
wire n_349;
wire n_1106;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_963;
wire n_745;
wire n_1052;
wire n_954;
wire n_627;
wire n_1116;
wire n_767;
wire n_206;
wire n_993;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_1059;
wire n_1084;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_647;
wire n_480;
wire n_607;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_707;
wire n_710;
wire n_679;
wire n_795;
wire n_695;
wire n_857;
wire n_832;
wire n_1072;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_207;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_768;
wire n_996;
wire n_921;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_1109;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_202;
wire n_1080;
wire n_266;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_868;
wire n_803;
wire n_1092;
wire n_238;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_890;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_187),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_126),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_21),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_158),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_194),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_182),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_48),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_92),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_186),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_10),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_106),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_10),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_195),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_185),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_181),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_120),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_17),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_15),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_31),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_17),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_141),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_184),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_68),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_133),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_155),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_105),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_108),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_53),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_12),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_166),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_113),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_50),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_28),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_16),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_139),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_136),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_96),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_173),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_149),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_159),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_111),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_190),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_49),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_145),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_9),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_160),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_23),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_125),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_94),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_22),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_104),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_63),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_188),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_167),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_142),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_117),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_51),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_66),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_99),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_154),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_196),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_112),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_138),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_191),
.Y(n_267)
);

BUFx10_ASAP7_75t_L g268 ( 
.A(n_9),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_89),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_47),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_228),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_212),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_247),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_199),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_214),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_261),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_201),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_214),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_247),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_219),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_209),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_264),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_214),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_204),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_237),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_253),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_205),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_206),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_268),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_216),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_208),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_216),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_211),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_258),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_263),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_258),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_220),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_214),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_223),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_200),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_232),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_202),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_213),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_248),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_203),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_210),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_250),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_215),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_217),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_218),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_221),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_224),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_214),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_226),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_227),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_236),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_268),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_230),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_233),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_266),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_235),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_275),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_318),
.A2(n_300),
.B1(n_302),
.B2(n_298),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_290),
.B(n_207),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_292),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_301),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_274),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_277),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_272),
.Y(n_330)
);

AND2x6_ASAP7_75t_L g331 ( 
.A(n_275),
.B(n_260),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_303),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_271),
.B(n_222),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_280),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_278),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_284),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_278),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_285),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_281),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_286),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_283),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_283),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_294),
.B(n_207),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_295),
.B(n_287),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_299),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_299),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_306),
.Y(n_347)
);

AND2x4_ASAP7_75t_L g348 ( 
.A(n_296),
.B(n_242),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_307),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_314),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_R g351 ( 
.A(n_288),
.B(n_229),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_314),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_291),
.B(n_225),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_310),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_312),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_277),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_317),
.B(n_313),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_293),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_319),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_320),
.B(n_225),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_304),
.B(n_265),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_322),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_309),
.B(n_265),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_276),
.B(n_260),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_321),
.B(n_231),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_321),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_311),
.B(n_251),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_315),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_308),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_316),
.B(n_308),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_273),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_282),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_289),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_297),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_298),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_300),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_R g377 ( 
.A(n_302),
.B(n_234),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_305),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_305),
.B(n_252),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_318),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_323),
.Y(n_381)
);

INVxp33_ASAP7_75t_L g382 ( 
.A(n_324),
.Y(n_382)
);

INVx2_ASAP7_75t_SL g383 ( 
.A(n_365),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_341),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_323),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_353),
.B(n_238),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_361),
.B(n_239),
.Y(n_387)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_341),
.Y(n_388)
);

NAND3xp33_ASAP7_75t_L g389 ( 
.A(n_325),
.B(n_262),
.C(n_260),
.Y(n_389)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_341),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_335),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_335),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_L g393 ( 
.A1(n_325),
.A2(n_343),
.B1(n_360),
.B2(n_348),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_367),
.B(n_363),
.Y(n_394)
);

OR2x6_ASAP7_75t_L g395 ( 
.A(n_372),
.B(n_260),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_337),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_337),
.Y(n_397)
);

BUFx10_ASAP7_75t_L g398 ( 
.A(n_344),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_369),
.B(n_273),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_345),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_345),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_341),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_370),
.B(n_279),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_350),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_341),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_350),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_352),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_333),
.B(n_240),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_343),
.B(n_241),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_L g410 ( 
.A1(n_360),
.A2(n_348),
.B1(n_357),
.B2(n_326),
.Y(n_410)
);

NAND2xp33_ASAP7_75t_SL g411 ( 
.A(n_374),
.B(n_279),
.Y(n_411)
);

AND2x2_ASAP7_75t_SL g412 ( 
.A(n_379),
.B(n_214),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_374),
.B(n_270),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_342),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_352),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_342),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_357),
.B(n_243),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_366),
.Y(n_418)
);

OR2x6_ASAP7_75t_L g419 ( 
.A(n_372),
.B(n_32),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_377),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_342),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_359),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_368),
.B(n_244),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_342),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_364),
.B(n_269),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g426 ( 
.A(n_366),
.B(n_245),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_368),
.B(n_351),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_342),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_346),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_339),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_327),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_346),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_368),
.B(n_267),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_365),
.B(n_246),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_328),
.B(n_259),
.Y(n_435)
);

AOI22x1_ASAP7_75t_L g436 ( 
.A1(n_348),
.A2(n_257),
.B1(n_256),
.B2(n_255),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_359),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_328),
.B(n_254),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_346),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_346),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_346),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_359),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_354),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_L g444 ( 
.A1(n_332),
.A2(n_214),
.B1(n_249),
.B2(n_2),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_354),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_336),
.B(n_0),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_354),
.B(n_33),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_354),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_354),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_371),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_355),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_379),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_355),
.Y(n_453)
);

INVxp33_ASAP7_75t_L g454 ( 
.A(n_376),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_362),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_422),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_394),
.B(n_362),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_381),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_422),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_437),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_426),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_418),
.B(n_330),
.Y(n_462)
);

NAND2x1p5_ASAP7_75t_L g463 ( 
.A(n_452),
.B(n_372),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_420),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_410),
.B(n_329),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_417),
.B(n_329),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_381),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_383),
.B(n_336),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_431),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_437),
.B(n_362),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_418),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_431),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_385),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_442),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_442),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_383),
.B(n_358),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_448),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_452),
.B(n_330),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_412),
.B(n_358),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_434),
.B(n_362),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_385),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_420),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_448),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_393),
.B(n_362),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_386),
.B(n_347),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_391),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_451),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_391),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_430),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_451),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_417),
.B(n_356),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_450),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_419),
.B(n_334),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_448),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_392),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_448),
.Y(n_496)
);

OAI221xp5_ASAP7_75t_L g497 ( 
.A1(n_444),
.A2(n_349),
.B1(n_338),
.B2(n_340),
.C(n_334),
.Y(n_497)
);

NAND3xp33_ASAP7_75t_L g498 ( 
.A(n_425),
.B(n_379),
.C(n_372),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_387),
.B(n_331),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_409),
.B(n_373),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_448),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_382),
.A2(n_371),
.B1(n_378),
.B2(n_375),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_419),
.B(n_338),
.Y(n_503)
);

AND2x6_ASAP7_75t_L g504 ( 
.A(n_421),
.B(n_372),
.Y(n_504)
);

AND2x6_ASAP7_75t_L g505 ( 
.A(n_421),
.B(n_373),
.Y(n_505)
);

INVx4_ASAP7_75t_L g506 ( 
.A(n_384),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_395),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_453),
.Y(n_508)
);

NAND2xp33_ASAP7_75t_L g509 ( 
.A(n_436),
.B(n_331),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_453),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_409),
.B(n_454),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_411),
.Y(n_512)
);

AO22x2_ASAP7_75t_L g513 ( 
.A1(n_446),
.A2(n_378),
.B1(n_375),
.B2(n_380),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_419),
.B(n_340),
.Y(n_514)
);

OAI22xp33_ASAP7_75t_SL g515 ( 
.A1(n_419),
.A2(n_373),
.B1(n_1),
.B2(n_2),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_427),
.B(n_376),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_450),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_426),
.B(n_376),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_412),
.B(n_331),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_397),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_392),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_395),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_397),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_399),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_412),
.B(n_331),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_419),
.B(n_376),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_423),
.A2(n_433),
.B1(n_413),
.B2(n_435),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_401),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_401),
.Y(n_529)
);

INVx8_ASAP7_75t_L g530 ( 
.A(n_395),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_398),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_403),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_404),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_404),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_395),
.Y(n_535)
);

NAND2xp33_ASAP7_75t_L g536 ( 
.A(n_436),
.B(n_331),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_398),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_415),
.Y(n_538)
);

OAI21xp33_ASAP7_75t_SL g539 ( 
.A1(n_519),
.A2(n_395),
.B(n_408),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_456),
.Y(n_540)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_469),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_456),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_532),
.B(n_376),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_457),
.B(n_415),
.Y(n_544)
);

OR2x6_ASAP7_75t_L g545 ( 
.A(n_530),
.B(n_438),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_484),
.A2(n_389),
.B1(n_455),
.B2(n_449),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_479),
.A2(n_455),
.B1(n_449),
.B2(n_445),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_518),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_469),
.B(n_443),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_459),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_485),
.B(n_424),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_510),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_471),
.B(n_424),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_478),
.B(n_429),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_491),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_469),
.B(n_443),
.Y(n_556)
);

BUFx2_ASAP7_75t_L g557 ( 
.A(n_517),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_466),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_478),
.B(n_429),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_524),
.B(n_398),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_459),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_472),
.B(n_384),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_460),
.B(n_396),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_465),
.B(n_396),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_460),
.B(n_474),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_475),
.B(n_400),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_528),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_472),
.B(n_493),
.Y(n_568)
);

NOR3xp33_ASAP7_75t_SL g569 ( 
.A(n_502),
.B(n_389),
.C(n_447),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_528),
.B(n_400),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_472),
.B(n_384),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_529),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_529),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_511),
.A2(n_449),
.B1(n_445),
.B2(n_443),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_493),
.A2(n_445),
.B1(n_441),
.B2(n_440),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_533),
.Y(n_576)
);

INVx5_ASAP7_75t_L g577 ( 
.A(n_507),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_533),
.B(n_406),
.Y(n_578)
);

BUFx5_ASAP7_75t_L g579 ( 
.A(n_504),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_461),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_503),
.B(n_384),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_492),
.A2(n_441),
.B1(n_440),
.B2(n_432),
.Y(n_582)
);

AND3x2_ASAP7_75t_SL g583 ( 
.A(n_515),
.B(n_0),
.C(n_1),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_500),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_473),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_503),
.A2(n_432),
.B1(n_414),
.B2(n_428),
.Y(n_586)
);

INVxp67_ASAP7_75t_L g587 ( 
.A(n_512),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_473),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_534),
.B(n_406),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_534),
.B(n_407),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_480),
.B(n_407),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_462),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_477),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_526),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_482),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_458),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_526),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_514),
.A2(n_402),
.B1(n_428),
.B2(n_416),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_462),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_520),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_487),
.B(n_402),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_514),
.B(n_384),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_489),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_523),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_595),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_542),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_558),
.A2(n_516),
.B1(n_498),
.B2(n_527),
.Y(n_607)
);

NOR2x1_ASAP7_75t_L g608 ( 
.A(n_541),
.B(n_468),
.Y(n_608)
);

BUFx2_ASAP7_75t_L g609 ( 
.A(n_557),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_561),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_594),
.A2(n_525),
.B1(n_507),
.B2(n_535),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_548),
.B(n_476),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_R g613 ( 
.A(n_555),
.B(n_464),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_564),
.A2(n_508),
.B1(n_490),
.B2(n_522),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_577),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_540),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_R g617 ( 
.A(n_560),
.B(n_531),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_552),
.B(n_507),
.Y(n_618)
);

INVx5_ASAP7_75t_L g619 ( 
.A(n_577),
.Y(n_619)
);

AO22x1_ASAP7_75t_L g620 ( 
.A1(n_543),
.A2(n_537),
.B1(n_505),
.B2(n_535),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_584),
.A2(n_513),
.B1(n_538),
.B2(n_497),
.Y(n_621)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_577),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_603),
.B(n_513),
.Y(n_623)
);

O2A1O1Ixp33_ASAP7_75t_L g624 ( 
.A1(n_587),
.A2(n_463),
.B(n_536),
.C(n_509),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_552),
.B(n_535),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_592),
.B(n_530),
.Y(n_626)
);

INVx5_ASAP7_75t_L g627 ( 
.A(n_545),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_541),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_599),
.B(n_477),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_597),
.A2(n_505),
.B1(n_504),
.B2(n_481),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_580),
.B(n_470),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_550),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_569),
.A2(n_567),
.B1(n_573),
.B2(n_572),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_600),
.B(n_467),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g635 ( 
.A(n_549),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_551),
.B(n_505),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_604),
.B(n_505),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_576),
.B(n_504),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_545),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_568),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_566),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_566),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_565),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g644 ( 
.A1(n_565),
.A2(n_598),
.B1(n_586),
.B2(n_575),
.Y(n_644)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_549),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_556),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_544),
.B(n_504),
.Y(n_647)
);

OR2x2_ASAP7_75t_L g648 ( 
.A(n_545),
.B(n_486),
.Y(n_648)
);

AO22x1_ASAP7_75t_L g649 ( 
.A1(n_583),
.A2(n_499),
.B1(n_495),
.B2(n_521),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_585),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_544),
.B(n_488),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_570),
.Y(n_652)
);

NOR2xp67_ASAP7_75t_L g653 ( 
.A(n_539),
.B(n_501),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_582),
.B(n_501),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_556),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_581),
.B(n_506),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_554),
.B(n_506),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_602),
.B(n_477),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_596),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_593),
.Y(n_660)
);

CKINVDCx11_ASAP7_75t_R g661 ( 
.A(n_588),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_593),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_562),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_570),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_605),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_606),
.Y(n_666)
);

OR2x2_ASAP7_75t_L g667 ( 
.A(n_609),
.B(n_559),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_619),
.Y(n_668)
);

OAI21xp5_ASAP7_75t_L g669 ( 
.A1(n_647),
.A2(n_546),
.B(n_574),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_619),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_625),
.B(n_571),
.Y(n_671)
);

INVx5_ASAP7_75t_L g672 ( 
.A(n_615),
.Y(n_672)
);

O2A1O1Ixp5_ASAP7_75t_L g673 ( 
.A1(n_620),
.A2(n_591),
.B(n_590),
.C(n_589),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_610),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_643),
.B(n_591),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_616),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_L g677 ( 
.A1(n_612),
.A2(n_547),
.B1(n_553),
.B2(n_601),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_635),
.B(n_601),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_619),
.Y(n_679)
);

BUFx2_ASAP7_75t_L g680 ( 
.A(n_613),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_659),
.Y(n_681)
);

INVxp67_ASAP7_75t_SL g682 ( 
.A(n_615),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_623),
.B(n_578),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_645),
.Y(n_684)
);

INVx4_ASAP7_75t_L g685 ( 
.A(n_615),
.Y(n_685)
);

OAI22xp5_ASAP7_75t_L g686 ( 
.A1(n_607),
.A2(n_590),
.B1(n_589),
.B2(n_578),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_655),
.B(n_563),
.Y(n_687)
);

NAND2x1p5_ASAP7_75t_L g688 ( 
.A(n_622),
.B(n_483),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_641),
.B(n_579),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_642),
.A2(n_563),
.B1(n_579),
.B2(n_416),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_617),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_632),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_612),
.Y(n_693)
);

BUFx4_ASAP7_75t_SL g694 ( 
.A(n_639),
.Y(n_694)
);

O2A1O1Ixp33_ASAP7_75t_SL g695 ( 
.A1(n_638),
.A2(n_579),
.B(n_428),
.C(n_416),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_652),
.Y(n_696)
);

HB1xp67_ASAP7_75t_L g697 ( 
.A(n_646),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_664),
.B(n_579),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_650),
.Y(n_699)
);

INVx1_ASAP7_75t_SL g700 ( 
.A(n_661),
.Y(n_700)
);

INVx4_ASAP7_75t_L g701 ( 
.A(n_622),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_628),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_631),
.B(n_579),
.Y(n_703)
);

INVx3_ASAP7_75t_SL g704 ( 
.A(n_627),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_640),
.B(n_483),
.Y(n_705)
);

BUFx12f_ASAP7_75t_L g706 ( 
.A(n_628),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_627),
.Y(n_707)
);

INVx4_ASAP7_75t_L g708 ( 
.A(n_628),
.Y(n_708)
);

BUFx12f_ASAP7_75t_L g709 ( 
.A(n_627),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_634),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_662),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_633),
.Y(n_712)
);

NAND2xp33_ASAP7_75t_L g713 ( 
.A(n_644),
.B(n_483),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_651),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_633),
.B(n_494),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_614),
.B(n_3),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_648),
.Y(n_717)
);

INVx5_ASAP7_75t_L g718 ( 
.A(n_660),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_660),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_SL g720 ( 
.A(n_654),
.B(n_494),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_656),
.Y(n_721)
);

BUFx12f_ASAP7_75t_L g722 ( 
.A(n_663),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_621),
.Y(n_723)
);

OAI21x1_ASAP7_75t_L g724 ( 
.A1(n_673),
.A2(n_624),
.B(n_653),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_681),
.B(n_608),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_666),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_706),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_718),
.Y(n_728)
);

OAI21x1_ASAP7_75t_SL g729 ( 
.A1(n_712),
.A2(n_621),
.B(n_637),
.Y(n_729)
);

NOR2xp67_ASAP7_75t_L g730 ( 
.A(n_691),
.B(n_626),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_681),
.B(n_649),
.Y(n_731)
);

BUFx2_ASAP7_75t_L g732 ( 
.A(n_697),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_666),
.Y(n_733)
);

OAI21x1_ASAP7_75t_L g734 ( 
.A1(n_689),
.A2(n_653),
.B(n_636),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_696),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_696),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_714),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_707),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_723),
.A2(n_618),
.B1(n_663),
.B2(n_657),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_683),
.B(n_663),
.Y(n_740)
);

INVx4_ASAP7_75t_L g741 ( 
.A(n_672),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_714),
.B(n_611),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_716),
.A2(n_629),
.B1(n_658),
.B2(n_656),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_718),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_706),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_710),
.B(n_658),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_674),
.Y(n_747)
);

OAI21x1_ASAP7_75t_L g748 ( 
.A1(n_689),
.A2(n_630),
.B(n_405),
.Y(n_748)
);

AOI21xp5_ASAP7_75t_SL g749 ( 
.A1(n_686),
.A2(n_496),
.B(n_494),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_687),
.B(n_34),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_699),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_699),
.Y(n_752)
);

OR2x2_ASAP7_75t_L g753 ( 
.A(n_675),
.B(n_402),
.Y(n_753)
);

NOR2x1_ASAP7_75t_SL g754 ( 
.A(n_715),
.B(n_496),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_721),
.B(n_35),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_670),
.Y(n_756)
);

OAI22xp5_ASAP7_75t_L g757 ( 
.A1(n_707),
.A2(n_496),
.B1(n_414),
.B2(n_405),
.Y(n_757)
);

CKINVDCx6p67_ASAP7_75t_R g758 ( 
.A(n_672),
.Y(n_758)
);

OAI21xp5_ASAP7_75t_L g759 ( 
.A1(n_677),
.A2(n_414),
.B(n_405),
.Y(n_759)
);

OAI21x1_ASAP7_75t_L g760 ( 
.A1(n_669),
.A2(n_390),
.B(n_388),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_676),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_717),
.B(n_3),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_693),
.A2(n_439),
.B1(n_390),
.B2(n_388),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_718),
.Y(n_764)
);

NOR2x1_ASAP7_75t_SL g765 ( 
.A(n_715),
.B(n_439),
.Y(n_765)
);

OAI21x1_ASAP7_75t_L g766 ( 
.A1(n_698),
.A2(n_390),
.B(n_388),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_692),
.Y(n_767)
);

AO21x2_ASAP7_75t_L g768 ( 
.A1(n_713),
.A2(n_695),
.B(n_703),
.Y(n_768)
);

AOI221xp5_ASAP7_75t_L g769 ( 
.A1(n_697),
.A2(n_439),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_684),
.Y(n_770)
);

OAI21x1_ASAP7_75t_L g771 ( 
.A1(n_690),
.A2(n_439),
.B(n_37),
.Y(n_771)
);

AO21x2_ASAP7_75t_L g772 ( 
.A1(n_713),
.A2(n_439),
.B(n_331),
.Y(n_772)
);

OAI21x1_ASAP7_75t_L g773 ( 
.A1(n_690),
.A2(n_38),
.B(n_36),
.Y(n_773)
);

OAI21xp5_ASAP7_75t_L g774 ( 
.A1(n_705),
.A2(n_4),
.B(n_5),
.Y(n_774)
);

OAI21x1_ASAP7_75t_L g775 ( 
.A1(n_721),
.A2(n_40),
.B(n_39),
.Y(n_775)
);

OAI21x1_ASAP7_75t_L g776 ( 
.A1(n_719),
.A2(n_42),
.B(n_41),
.Y(n_776)
);

OAI21xp5_ASAP7_75t_L g777 ( 
.A1(n_705),
.A2(n_4),
.B(n_6),
.Y(n_777)
);

A2O1A1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_720),
.A2(n_7),
.B(n_8),
.C(n_11),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_671),
.B(n_43),
.Y(n_779)
);

OAI22xp5_ASAP7_75t_L g780 ( 
.A1(n_704),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_780)
);

OAI21xp33_ASAP7_75t_L g781 ( 
.A1(n_667),
.A2(n_13),
.B(n_14),
.Y(n_781)
);

OA21x2_ASAP7_75t_L g782 ( 
.A1(n_671),
.A2(n_13),
.B(n_14),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_670),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_718),
.Y(n_784)
);

BUFx2_ASAP7_75t_L g785 ( 
.A(n_722),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_678),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_678),
.Y(n_787)
);

OAI21x1_ASAP7_75t_L g788 ( 
.A1(n_688),
.A2(n_45),
.B(n_44),
.Y(n_788)
);

OAI21x1_ASAP7_75t_L g789 ( 
.A1(n_688),
.A2(n_695),
.B(n_682),
.Y(n_789)
);

BUFx3_ASAP7_75t_L g790 ( 
.A(n_672),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_727),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_727),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_747),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_761),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_732),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_740),
.B(n_678),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_745),
.Y(n_797)
);

OAI21x1_ASAP7_75t_L g798 ( 
.A1(n_724),
.A2(n_702),
.B(n_671),
.Y(n_798)
);

AND2x2_ASAP7_75t_SL g799 ( 
.A(n_782),
.B(n_680),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_761),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_SL g801 ( 
.A1(n_774),
.A2(n_709),
.B1(n_700),
.B2(n_722),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_732),
.Y(n_802)
);

OAI22xp5_ASAP7_75t_L g803 ( 
.A1(n_731),
.A2(n_704),
.B1(n_709),
.B2(n_665),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_735),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_781),
.A2(n_777),
.B1(n_769),
.B2(n_780),
.Y(n_805)
);

AO21x2_ASAP7_75t_L g806 ( 
.A1(n_749),
.A2(n_702),
.B(n_670),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_738),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_756),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_737),
.B(n_670),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_725),
.A2(n_668),
.B1(n_679),
.B2(n_672),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_779),
.A2(n_679),
.B1(n_668),
.B2(n_708),
.Y(n_811)
);

INVx4_ASAP7_75t_L g812 ( 
.A(n_758),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_745),
.Y(n_813)
);

BUFx10_ASAP7_75t_L g814 ( 
.A(n_756),
.Y(n_814)
);

OR2x6_ASAP7_75t_L g815 ( 
.A(n_749),
.B(n_708),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_726),
.Y(n_816)
);

NOR2xp67_ASAP7_75t_L g817 ( 
.A(n_730),
.B(n_701),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_735),
.Y(n_818)
);

CKINVDCx11_ASAP7_75t_R g819 ( 
.A(n_738),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_786),
.B(n_711),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_SL g821 ( 
.A1(n_782),
.A2(n_779),
.B1(n_773),
.B2(n_754),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_737),
.B(n_701),
.Y(n_822)
);

BUFx12f_ASAP7_75t_L g823 ( 
.A(n_785),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_787),
.B(n_711),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_779),
.A2(n_685),
.B1(n_694),
.B2(n_18),
.Y(n_825)
);

INVx4_ASAP7_75t_SL g826 ( 
.A(n_790),
.Y(n_826)
);

INVx4_ASAP7_75t_L g827 ( 
.A(n_758),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_740),
.B(n_685),
.Y(n_828)
);

OR2x2_ASAP7_75t_L g829 ( 
.A(n_770),
.B(n_15),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_SL g830 ( 
.A1(n_782),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_750),
.B(n_46),
.Y(n_831)
);

AND3x2_ASAP7_75t_L g832 ( 
.A(n_784),
.B(n_755),
.C(n_778),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_756),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_SL g834 ( 
.A1(n_773),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_SL g835 ( 
.A1(n_778),
.A2(n_765),
.B1(n_771),
.B2(n_729),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_736),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_768),
.Y(n_837)
);

NOR2x1_ASAP7_75t_SL g838 ( 
.A(n_768),
.B(n_52),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_736),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_750),
.A2(n_743),
.B1(n_739),
.B2(n_762),
.Y(n_840)
);

NOR3xp33_ASAP7_75t_SL g841 ( 
.A(n_746),
.B(n_20),
.C(n_22),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_751),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_742),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_742),
.B(n_54),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_733),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_767),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_724),
.A2(n_122),
.B(n_198),
.Y(n_847)
);

BUFx2_ASAP7_75t_L g848 ( 
.A(n_756),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_760),
.A2(n_121),
.B(n_197),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_751),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_752),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_783),
.B(n_55),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_752),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_784),
.Y(n_854)
);

OAI21x1_ASAP7_75t_SL g855 ( 
.A1(n_759),
.A2(n_24),
.B(n_25),
.Y(n_855)
);

AOI221xp5_ASAP7_75t_L g856 ( 
.A1(n_753),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.C(n_29),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_768),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_793),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_795),
.Y(n_859)
);

OAI21x1_ASAP7_75t_L g860 ( 
.A1(n_847),
.A2(n_849),
.B(n_766),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_795),
.B(n_753),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_792),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_796),
.B(n_755),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_802),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_802),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_846),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_794),
.B(n_783),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_828),
.B(n_783),
.Y(n_868)
);

CKINVDCx16_ASAP7_75t_R g869 ( 
.A(n_823),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_800),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_826),
.B(n_783),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_819),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_854),
.Y(n_873)
);

OAI22xp33_ASAP7_75t_L g874 ( 
.A1(n_856),
.A2(n_741),
.B1(n_790),
.B2(n_764),
.Y(n_874)
);

OR2x2_ASAP7_75t_L g875 ( 
.A(n_816),
.B(n_734),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_845),
.Y(n_876)
);

OR2x6_ASAP7_75t_L g877 ( 
.A(n_815),
.B(n_775),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_798),
.Y(n_878)
);

INVxp33_ASAP7_75t_SL g879 ( 
.A(n_807),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_805),
.A2(n_763),
.B1(n_757),
.B2(n_741),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_801),
.B(n_728),
.Y(n_881)
);

A2O1A1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_841),
.A2(n_775),
.B(n_771),
.C(n_788),
.Y(n_882)
);

NAND2xp33_ASAP7_75t_SL g883 ( 
.A(n_841),
.B(n_741),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_805),
.A2(n_776),
.B1(n_728),
.B2(n_764),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_791),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_792),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_804),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_815),
.A2(n_760),
.B(n_772),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_820),
.B(n_728),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_850),
.B(n_734),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_792),
.Y(n_891)
);

NAND2x1p5_ASAP7_75t_L g892 ( 
.A(n_812),
.B(n_744),
.Y(n_892)
);

INVx5_ASAP7_75t_L g893 ( 
.A(n_815),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_797),
.Y(n_894)
);

OR2x2_ASAP7_75t_L g895 ( 
.A(n_853),
.B(n_766),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_818),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_836),
.B(n_744),
.Y(n_897)
);

NAND3xp33_ASAP7_75t_SL g898 ( 
.A(n_801),
.B(n_776),
.C(n_788),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_SL g899 ( 
.A1(n_855),
.A2(n_764),
.B1(n_744),
.B2(n_789),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_826),
.B(n_789),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_R g901 ( 
.A(n_797),
.B(n_56),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_826),
.B(n_748),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_825),
.A2(n_772),
.B1(n_748),
.B2(n_29),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_839),
.B(n_26),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_848),
.B(n_772),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_858),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_858),
.Y(n_907)
);

INVxp67_ASAP7_75t_L g908 ( 
.A(n_873),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_866),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_859),
.B(n_799),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_876),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_900),
.B(n_837),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_864),
.Y(n_913)
);

OAI31xp33_ASAP7_75t_SL g914 ( 
.A1(n_874),
.A2(n_830),
.A3(n_856),
.B(n_834),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_865),
.B(n_861),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_875),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_896),
.B(n_799),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_900),
.Y(n_918)
);

OAI221xp5_ASAP7_75t_L g919 ( 
.A1(n_882),
.A2(n_834),
.B1(n_830),
.B2(n_840),
.C(n_843),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_878),
.B(n_837),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_870),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_868),
.B(n_857),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_890),
.B(n_857),
.Y(n_923)
);

OR2x2_ASAP7_75t_L g924 ( 
.A(n_895),
.B(n_887),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_889),
.B(n_821),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_897),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_902),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_863),
.B(n_821),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_893),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_902),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_L g931 ( 
.A1(n_881),
.A2(n_844),
.B1(n_803),
.B2(n_832),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_905),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_905),
.Y(n_933)
);

INVxp67_ASAP7_75t_SL g934 ( 
.A(n_867),
.Y(n_934)
);

OR2x2_ASAP7_75t_L g935 ( 
.A(n_888),
.B(n_829),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_893),
.B(n_835),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_893),
.B(n_835),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_877),
.B(n_842),
.Y(n_938)
);

OAI21xp33_ASAP7_75t_SL g939 ( 
.A1(n_914),
.A2(n_884),
.B(n_877),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_934),
.B(n_899),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_925),
.B(n_869),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_919),
.A2(n_811),
.B1(n_880),
.B2(n_886),
.Y(n_942)
);

NAND3xp33_ASAP7_75t_L g943 ( 
.A(n_914),
.B(n_883),
.C(n_904),
.Y(n_943)
);

OAI21xp33_ASAP7_75t_L g944 ( 
.A1(n_919),
.A2(n_898),
.B(n_901),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_SL g945 ( 
.A(n_936),
.B(n_872),
.Y(n_945)
);

NAND3xp33_ASAP7_75t_L g946 ( 
.A(n_935),
.B(n_931),
.C(n_917),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_925),
.B(n_891),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_935),
.A2(n_849),
.B(n_847),
.Y(n_948)
);

NOR3xp33_ASAP7_75t_SL g949 ( 
.A(n_917),
.B(n_885),
.C(n_810),
.Y(n_949)
);

OAI221xp5_ASAP7_75t_L g950 ( 
.A1(n_915),
.A2(n_892),
.B1(n_817),
.B2(n_824),
.C(n_903),
.Y(n_950)
);

AOI22xp33_ASAP7_75t_SL g951 ( 
.A1(n_936),
.A2(n_838),
.B1(n_879),
.B2(n_832),
.Y(n_951)
);

NAND3xp33_ASAP7_75t_L g952 ( 
.A(n_926),
.B(n_852),
.C(n_812),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_926),
.B(n_862),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_922),
.B(n_862),
.Y(n_954)
);

AOI211xp5_ASAP7_75t_SL g955 ( 
.A1(n_937),
.A2(n_871),
.B(n_831),
.C(n_809),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_922),
.B(n_862),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_915),
.B(n_908),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_908),
.B(n_894),
.Y(n_958)
);

OA21x2_ASAP7_75t_L g959 ( 
.A1(n_920),
.A2(n_860),
.B(n_809),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_937),
.B(n_894),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_939),
.B(n_945),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_960),
.B(n_918),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_957),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_946),
.B(n_910),
.Y(n_964)
);

NAND2x1_ASAP7_75t_L g965 ( 
.A(n_959),
.B(n_929),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_960),
.B(n_918),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_941),
.B(n_918),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_947),
.B(n_927),
.Y(n_968)
);

OR2x2_ASAP7_75t_L g969 ( 
.A(n_940),
.B(n_924),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_954),
.B(n_927),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_956),
.B(n_927),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_959),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_953),
.Y(n_973)
);

INVxp67_ASAP7_75t_SL g974 ( 
.A(n_958),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_959),
.B(n_930),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_948),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_955),
.B(n_930),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_976),
.B(n_943),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_962),
.B(n_930),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_977),
.B(n_928),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_977),
.B(n_932),
.Y(n_981)
);

OR3x2_ASAP7_75t_L g982 ( 
.A(n_961),
.B(n_944),
.C(n_963),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_962),
.B(n_966),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_964),
.B(n_928),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_972),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_973),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_966),
.B(n_932),
.Y(n_987)
);

INVx2_ASAP7_75t_SL g988 ( 
.A(n_967),
.Y(n_988)
);

NOR2x1p5_ASAP7_75t_L g989 ( 
.A(n_974),
.B(n_952),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_967),
.B(n_968),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_990),
.B(n_968),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_982),
.A2(n_961),
.B1(n_951),
.B2(n_942),
.Y(n_992)
);

OA222x2_ASAP7_75t_L g993 ( 
.A1(n_982),
.A2(n_972),
.B1(n_969),
.B2(n_965),
.C1(n_949),
.C2(n_951),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_986),
.Y(n_994)
);

INVxp67_ASAP7_75t_L g995 ( 
.A(n_978),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_985),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_990),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_980),
.B(n_968),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_983),
.B(n_970),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_999),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_992),
.B(n_988),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_995),
.B(n_988),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_991),
.B(n_981),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_995),
.B(n_997),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_998),
.B(n_981),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_1004),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_1002),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_1001),
.A2(n_993),
.B(n_998),
.Y(n_1008)
);

OAI221xp5_ASAP7_75t_L g1009 ( 
.A1(n_1000),
.A2(n_994),
.B1(n_984),
.B2(n_996),
.C(n_949),
.Y(n_1009)
);

AOI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_1005),
.A2(n_989),
.B1(n_979),
.B2(n_950),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_1003),
.B(n_987),
.Y(n_1011)
);

OAI221xp5_ASAP7_75t_L g1012 ( 
.A1(n_1001),
.A2(n_985),
.B1(n_929),
.B2(n_975),
.C(n_913),
.Y(n_1012)
);

OAI21xp33_ASAP7_75t_L g1013 ( 
.A1(n_1001),
.A2(n_979),
.B(n_975),
.Y(n_1013)
);

INVxp67_ASAP7_75t_SL g1014 ( 
.A(n_1001),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_1001),
.B(n_979),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_1014),
.B(n_970),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1006),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_1007),
.B(n_797),
.Y(n_1018)
);

AOI211xp5_ASAP7_75t_L g1019 ( 
.A1(n_1008),
.A2(n_813),
.B(n_894),
.C(n_871),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_1015),
.B(n_971),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_1010),
.A2(n_933),
.B1(n_932),
.B2(n_971),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1011),
.Y(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_1009),
.A2(n_921),
.B(n_822),
.C(n_909),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_1013),
.A2(n_827),
.B(n_911),
.Y(n_1024)
);

AO22x1_ASAP7_75t_L g1025 ( 
.A1(n_1018),
.A2(n_813),
.B1(n_1012),
.B2(n_827),
.Y(n_1025)
);

NAND2x1_ASAP7_75t_L g1026 ( 
.A(n_1016),
.B(n_813),
.Y(n_1026)
);

AOI322xp5_ASAP7_75t_L g1027 ( 
.A1(n_1017),
.A2(n_910),
.A3(n_920),
.B1(n_933),
.B2(n_912),
.C1(n_923),
.C2(n_909),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_1019),
.A2(n_911),
.B(n_916),
.C(n_938),
.Y(n_1028)
);

AOI21xp33_ASAP7_75t_L g1029 ( 
.A1(n_1022),
.A2(n_27),
.B(n_30),
.Y(n_1029)
);

AOI221xp5_ASAP7_75t_L g1030 ( 
.A1(n_1023),
.A2(n_916),
.B1(n_820),
.B2(n_938),
.C(n_907),
.Y(n_1030)
);

OAI221xp5_ASAP7_75t_L g1031 ( 
.A1(n_1024),
.A2(n_916),
.B1(n_924),
.B2(n_933),
.C(n_907),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1020),
.B(n_1021),
.Y(n_1032)
);

NOR2x1_ASAP7_75t_L g1033 ( 
.A(n_1026),
.B(n_1032),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1029),
.B(n_923),
.Y(n_1034)
);

AOI21xp33_ASAP7_75t_SL g1035 ( 
.A1(n_1025),
.A2(n_30),
.B(n_57),
.Y(n_1035)
);

NOR3xp33_ASAP7_75t_L g1036 ( 
.A(n_1031),
.B(n_833),
.C(n_808),
.Y(n_1036)
);

OAI21xp33_ASAP7_75t_L g1037 ( 
.A1(n_1028),
.A2(n_1027),
.B(n_1030),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_1026),
.Y(n_1038)
);

NOR2x1_ASAP7_75t_L g1039 ( 
.A(n_1026),
.B(n_806),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_1038),
.B(n_938),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_SL g1041 ( 
.A1(n_1035),
.A2(n_822),
.B(n_906),
.Y(n_1041)
);

NAND3xp33_ASAP7_75t_SL g1042 ( 
.A(n_1037),
.B(n_906),
.C(n_851),
.Y(n_1042)
);

OAI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_1034),
.A2(n_833),
.B1(n_808),
.B2(n_906),
.Y(n_1043)
);

AOI221xp5_ASAP7_75t_L g1044 ( 
.A1(n_1036),
.A2(n_938),
.B1(n_912),
.B2(n_806),
.C(n_61),
.Y(n_1044)
);

OA22x2_ASAP7_75t_L g1045 ( 
.A1(n_1033),
.A2(n_912),
.B1(n_814),
.B2(n_60),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_1039),
.B(n_814),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1040),
.Y(n_1047)
);

NAND3xp33_ASAP7_75t_SL g1048 ( 
.A(n_1044),
.B(n_58),
.C(n_59),
.Y(n_1048)
);

NOR2x1p5_ASAP7_75t_L g1049 ( 
.A(n_1042),
.B(n_912),
.Y(n_1049)
);

NOR2x1_ASAP7_75t_L g1050 ( 
.A(n_1046),
.B(n_62),
.Y(n_1050)
);

NAND3xp33_ASAP7_75t_L g1051 ( 
.A(n_1043),
.B(n_64),
.C(n_65),
.Y(n_1051)
);

NAND3xp33_ASAP7_75t_L g1052 ( 
.A(n_1045),
.B(n_67),
.C(n_69),
.Y(n_1052)
);

NOR3x1_ASAP7_75t_L g1053 ( 
.A(n_1041),
.B(n_70),
.C(n_71),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_1047),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_1054)
);

NOR2x1_ASAP7_75t_L g1055 ( 
.A(n_1052),
.B(n_75),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1053),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1050),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1049),
.Y(n_1058)
);

INVxp67_ASAP7_75t_SL g1059 ( 
.A(n_1051),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1048),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1047),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_1053),
.Y(n_1062)
);

INVx2_ASAP7_75t_SL g1063 ( 
.A(n_1057),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1062),
.B(n_76),
.Y(n_1064)
);

NOR3xp33_ASAP7_75t_L g1065 ( 
.A(n_1061),
.B(n_77),
.C(n_78),
.Y(n_1065)
);

OAI222xp33_ASAP7_75t_L g1066 ( 
.A1(n_1056),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.C1(n_82),
.C2(n_83),
.Y(n_1066)
);

NAND3xp33_ASAP7_75t_SL g1067 ( 
.A(n_1060),
.B(n_84),
.C(n_85),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1058),
.B(n_86),
.Y(n_1068)
);

NOR2x1_ASAP7_75t_L g1069 ( 
.A(n_1055),
.B(n_87),
.Y(n_1069)
);

OAI311xp33_ASAP7_75t_L g1070 ( 
.A1(n_1059),
.A2(n_88),
.A3(n_90),
.B1(n_91),
.C1(n_93),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_1063),
.Y(n_1071)
);

INVx1_ASAP7_75t_SL g1072 ( 
.A(n_1069),
.Y(n_1072)
);

HB1xp67_ASAP7_75t_L g1073 ( 
.A(n_1064),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1068),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_1065),
.A2(n_1054),
.B(n_97),
.C(n_98),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_R g1076 ( 
.A(n_1067),
.B(n_1054),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_1070),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1066),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_1063),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_1071),
.Y(n_1080)
);

AOI22xp33_ASAP7_75t_SL g1081 ( 
.A1(n_1079),
.A2(n_95),
.B1(n_100),
.B2(n_101),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1073),
.B(n_102),
.Y(n_1082)
);

AND3x4_ASAP7_75t_L g1083 ( 
.A(n_1077),
.B(n_103),
.C(n_107),
.Y(n_1083)
);

NOR3xp33_ASAP7_75t_L g1084 ( 
.A(n_1072),
.B(n_109),
.C(n_110),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_1078),
.B(n_114),
.Y(n_1085)
);

AOI221xp5_ASAP7_75t_L g1086 ( 
.A1(n_1076),
.A2(n_115),
.B1(n_116),
.B2(n_118),
.C(n_119),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1074),
.Y(n_1087)
);

OAI211xp5_ASAP7_75t_SL g1088 ( 
.A1(n_1075),
.A2(n_123),
.B(n_124),
.C(n_127),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1073),
.B(n_128),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1071),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_1071),
.Y(n_1091)
);

CKINVDCx20_ASAP7_75t_R g1092 ( 
.A(n_1071),
.Y(n_1092)
);

INVx1_ASAP7_75t_SL g1093 ( 
.A(n_1092),
.Y(n_1093)
);

OA22x2_ASAP7_75t_L g1094 ( 
.A1(n_1090),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_R g1095 ( 
.A(n_1091),
.B(n_132),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1091),
.B(n_134),
.Y(n_1096)
);

OR2x2_ASAP7_75t_L g1097 ( 
.A(n_1080),
.B(n_135),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1089),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1085),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1082),
.A2(n_137),
.B(n_140),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1083),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1093),
.A2(n_1087),
.B1(n_1086),
.B2(n_1081),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_1101),
.A2(n_1084),
.B1(n_1088),
.B2(n_146),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1097),
.Y(n_1104)
);

NOR2x1p5_ASAP7_75t_L g1105 ( 
.A(n_1096),
.B(n_143),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1098),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_1095),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_1106),
.Y(n_1108)
);

OAI222xp33_ASAP7_75t_L g1109 ( 
.A1(n_1102),
.A2(n_1099),
.B1(n_1094),
.B2(n_1100),
.C1(n_150),
.C2(n_151),
.Y(n_1109)
);

OR2x6_ASAP7_75t_L g1110 ( 
.A(n_1107),
.B(n_144),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_1108),
.A2(n_1104),
.B(n_1103),
.C(n_1105),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1111),
.Y(n_1112)
);

AND3x1_ASAP7_75t_L g1113 ( 
.A(n_1112),
.B(n_1109),
.C(n_1110),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_1112),
.A2(n_147),
.B(n_148),
.Y(n_1114)
);

OAI22xp33_ASAP7_75t_L g1115 ( 
.A1(n_1113),
.A2(n_152),
.B1(n_153),
.B2(n_156),
.Y(n_1115)
);

OAI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1114),
.A2(n_157),
.B1(n_161),
.B2(n_162),
.Y(n_1116)
);

OAI22xp33_ASAP7_75t_L g1117 ( 
.A1(n_1113),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1115),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1117),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_1119)
);

AOI221xp5_ASAP7_75t_L g1120 ( 
.A1(n_1116),
.A2(n_176),
.B1(n_178),
.B2(n_179),
.C(n_180),
.Y(n_1120)
);

AOI211xp5_ASAP7_75t_L g1121 ( 
.A1(n_1119),
.A2(n_1120),
.B(n_1118),
.C(n_183),
.Y(n_1121)
);


endmodule