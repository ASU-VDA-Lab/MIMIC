module real_jpeg_25188_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_288;
wire n_166;
wire n_176;
wire n_292;
wire n_215;
wire n_221;
wire n_249;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_293;
wire n_164;
wire n_275;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_0),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_0),
.B(n_51),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_0),
.B(n_25),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_0),
.B(n_36),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_0),
.B(n_17),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_0),
.B(n_31),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_0),
.B(n_45),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_0),
.B(n_43),
.Y(n_237)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_3),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_3),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_3),
.B(n_43),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_3),
.B(n_25),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_3),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_3),
.B(n_36),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_3),
.B(n_31),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_3),
.B(n_45),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_4),
.B(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_6),
.B(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_6),
.B(n_45),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_6),
.B(n_36),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_6),
.Y(n_113)
);

INVx8_ASAP7_75t_SL g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_8),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_8),
.B(n_69),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_8),
.B(n_43),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_8),
.B(n_25),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_8),
.B(n_45),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_8),
.B(n_62),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_8),
.B(n_36),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_8),
.B(n_31),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_9),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_9),
.B(n_45),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_9),
.B(n_36),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_9),
.B(n_43),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_9),
.B(n_25),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_9),
.B(n_51),
.Y(n_241)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_11),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_11),
.B(n_43),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_11),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_11),
.B(n_31),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_11),
.B(n_62),
.Y(n_134)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_13),
.B(n_51),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_13),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_13),
.B(n_25),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_13),
.B(n_31),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_13),
.B(n_17),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_13),
.B(n_36),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_43),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_15),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_15),
.B(n_36),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_15),
.B(n_31),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_15),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_16),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_16),
.B(n_51),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_16),
.B(n_31),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_16),
.B(n_36),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_16),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_16),
.B(n_45),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_16),
.B(n_43),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_16),
.B(n_25),
.Y(n_242)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_17),
.Y(n_114)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_17),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_153),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_123),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_93),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_53),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_33),
.B2(n_38),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_32),
.B(n_145),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_33),
.A2(n_38),
.B1(n_60),
.B2(n_64),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_33),
.B(n_56),
.C(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_34),
.B(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_35),
.B(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_47),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.C(n_44),
.Y(n_40)
);

FAx1_ASAP7_75t_SL g71 ( 
.A(n_41),
.B(n_42),
.CI(n_44),
.CON(n_71),
.SN(n_71)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx24_ASAP7_75t_SL g294 ( 
.A(n_47),
.Y(n_294)
);

FAx1_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_49),
.CI(n_50),
.CON(n_47),
.SN(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_51),
.Y(n_58)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_72),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_65),
.C(n_71),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_55),
.B(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_60),
.A2(n_64),
.B1(n_66),
.B2(n_105),
.Y(n_104)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_63),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_66),
.C(n_67),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_65),
.B(n_71),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_66),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_67),
.A2(n_68),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

BUFx24_ASAP7_75t_SL g299 ( 
.A(n_71),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_87),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_84),
.C(n_85),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_74),
.A2(n_75),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_78),
.C(n_81),
.Y(n_75)
);

FAx1_ASAP7_75t_SL g95 ( 
.A(n_76),
.B(n_78),
.CI(n_81),
.CON(n_95),
.SN(n_95)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_82),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_84),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_84),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_84),
.A2(n_85),
.B1(n_91),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_85),
.Y(n_108)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_86),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_92),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_89),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_106),
.C(n_110),
.Y(n_93)
);

FAx1_ASAP7_75t_SL g125 ( 
.A(n_94),
.B(n_106),
.CI(n_110),
.CON(n_125),
.SN(n_125)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.C(n_102),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_95),
.B(n_286),
.Y(n_285)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_95),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_96),
.B(n_102),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.C(n_100),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_97),
.A2(n_98),
.B1(n_100),
.B2(n_101),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_99),
.B(n_273),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_107),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_121),
.C(n_122),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_115),
.C(n_119),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_119),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_115),
.B(n_132),
.Y(n_131)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_122),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.C(n_129),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_293)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx24_ASAP7_75t_SL g298 ( 
.A(n_125),
.Y(n_298)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_129),
.B(n_293),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_140),
.C(n_142),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_130),
.B(n_288),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.C(n_136),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_131),
.B(n_279),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_133),
.A2(n_134),
.B(n_135),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_133),
.B(n_136),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.C(n_139),
.Y(n_136)
);

FAx1_ASAP7_75t_SL g252 ( 
.A(n_137),
.B(n_138),
.CI(n_139),
.CON(n_252),
.SN(n_252)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_140),
.B(n_142),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_149),
.C(n_151),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_143),
.B(n_275),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.C(n_148),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_144),
.B(n_263),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_147),
.B(n_148),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_149),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_291),
.C(n_292),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_281),
.C(n_282),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_266),
.C(n_267),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_245),
.C(n_246),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_223),
.C(n_224),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_205),
.C(n_206),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_185),
.C(n_186),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_173),
.C(n_178),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_169),
.B2(n_170),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_171),
.C(n_172),
.Y(n_185)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_164),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_168),
.Y(n_189)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.C(n_181),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_196),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_191),
.C(n_196),
.Y(n_205)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_192),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_193),
.B(n_195),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_204),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_197),
.Y(n_204)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_200),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_203),
.C(n_204),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_214),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_209),
.C(n_214),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_212),
.C(n_213),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_217),
.C(n_218),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_219),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_222),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_239),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_240),
.C(n_244),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_235),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_234),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_234),
.C(n_235),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_228),
.Y(n_233)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_233),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx24_ASAP7_75t_SL g297 ( 
.A(n_235),
.Y(n_297)
);

FAx1_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_237),
.CI(n_238),
.CON(n_235),
.SN(n_235)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_237),
.C(n_238),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_244),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_240),
.Y(n_259)
);

FAx1_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_242),
.CI(n_243),
.CON(n_240),
.SN(n_240)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_258),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_250),
.C(n_258),
.Y(n_266)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_254),
.C(n_257),
.Y(n_270)
);

BUFx24_ASAP7_75t_SL g295 ( 
.A(n_252),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_256),
.B2(n_257),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_262),
.C(n_264),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_264),
.B2(n_265),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_261),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_262),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_276),
.B2(n_280),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_277),
.C(n_278),
.Y(n_281)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_272),
.C(n_274),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_276),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_289),
.B2(n_290),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_283),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_284),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_287),
.C(n_289),
.Y(n_291)
);


endmodule