module fake_netlist_1_2484_n_16 (n_1, n_2, n_4, n_3, n_0, n_16);
input n_1;
input n_2;
input n_4;
input n_3;
input n_0;
output n_16;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
CKINVDCx5p33_ASAP7_75t_R g5 ( .A(n_3), .Y(n_5) );
BUFx3_ASAP7_75t_L g6 ( .A(n_4), .Y(n_6) );
AND2x2_ASAP7_75t_L g7 ( .A(n_6), .B(n_0), .Y(n_7) );
NOR3xp33_ASAP7_75t_SL g8 ( .A(n_5), .B(n_1), .C(n_2), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_7), .Y(n_9) );
NAND2x1p5_ASAP7_75t_L g10 ( .A(n_9), .B(n_8), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_10), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_11), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_13), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g15 ( .A(n_14), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
endmodule