module fake_jpeg_31638_n_541 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_541);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_541;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_419;
wire n_378;
wire n_133;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx11_ASAP7_75t_L g153 ( 
.A(n_56),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_9),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_57),
.B(n_73),
.Y(n_151)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_63),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

CKINVDCx9p33_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx2_ASAP7_75t_R g152 ( 
.A(n_65),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_69),
.Y(n_148)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_17),
.B(n_8),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_75),
.Y(n_160)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_76),
.Y(n_156)
);

BUFx16f_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_77),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_80),
.Y(n_155)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_82),
.Y(n_162)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_47),
.A2(n_16),
.B1(n_8),
.B2(n_10),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_86),
.A2(n_27),
.B1(n_36),
.B2(n_49),
.Y(n_140)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_88),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_17),
.B(n_7),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_91),
.B(n_48),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_94),
.Y(n_149)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_95),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_18),
.B(n_7),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_50),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_99),
.Y(n_165)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_100),
.Y(n_168)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_103),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_30),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_102),
.B(n_43),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_26),
.Y(n_104)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_30),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_77),
.B(n_18),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_106),
.B(n_110),
.Y(n_177)
);

AOI21xp33_ASAP7_75t_L g110 ( 
.A1(n_86),
.A2(n_51),
.B(n_26),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_102),
.B(n_28),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_112),
.B(n_132),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_122),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_89),
.A2(n_43),
.B1(n_30),
.B2(n_51),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_124),
.A2(n_125),
.B1(n_56),
.B2(n_63),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_99),
.A2(n_93),
.B1(n_66),
.B2(n_78),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_127),
.B(n_145),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_50),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_140),
.A2(n_44),
.B(n_32),
.Y(n_173)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_40),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_96),
.B(n_40),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_164),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_79),
.B(n_28),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_150),
.B(n_154),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_84),
.B(n_34),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_54),
.A2(n_43),
.B1(n_36),
.B2(n_27),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_157),
.A2(n_49),
.B1(n_37),
.B2(n_48),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_152),
.Y(n_174)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_109),
.Y(n_171)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_171),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_152),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_172),
.B(n_197),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_173),
.A2(n_221),
.B(n_6),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_174),
.B(n_179),
.Y(n_248)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_175),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_176),
.A2(n_182),
.B1(n_184),
.B2(n_191),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_118),
.B(n_69),
.C(n_95),
.Y(n_178)
);

FAx1_ASAP7_75t_SL g266 ( 
.A(n_178),
.B(n_200),
.CI(n_202),
.CON(n_266),
.SN(n_266)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_166),
.Y(n_179)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_180),
.Y(n_224)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_181),
.Y(n_247)
);

AO22x2_ASAP7_75t_SL g183 ( 
.A1(n_157),
.A2(n_87),
.B1(n_76),
.B2(n_75),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_L g236 ( 
.A1(n_183),
.A2(n_220),
.B1(n_222),
.B2(n_138),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_125),
.A2(n_85),
.B1(n_55),
.B2(n_67),
.Y(n_184)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_121),
.Y(n_187)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

AO22x1_ASAP7_75t_SL g188 ( 
.A1(n_115),
.A2(n_64),
.B1(n_62),
.B2(n_80),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_188),
.B(n_108),
.Y(n_243)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_131),
.Y(n_189)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_189),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_114),
.A2(n_37),
.B1(n_32),
.B2(n_44),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_190),
.A2(n_209),
.B1(n_166),
.B2(n_160),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_124),
.A2(n_80),
.B1(n_43),
.B2(n_34),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_192),
.Y(n_238)
);

AO22x2_ASAP7_75t_L g194 ( 
.A1(n_156),
.A2(n_43),
.B1(n_29),
.B2(n_21),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_194),
.B(n_206),
.Y(n_255)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_195),
.Y(n_252)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_130),
.Y(n_196)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_196),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_123),
.Y(n_197)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_149),
.Y(n_199)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

AND2x2_ASAP7_75t_SL g200 ( 
.A(n_107),
.B(n_0),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_130),
.Y(n_201)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_151),
.B(n_117),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_137),
.Y(n_203)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

BUFx4f_ASAP7_75t_SL g204 ( 
.A(n_129),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g254 ( 
.A(n_204),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_139),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_205),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_156),
.A2(n_60),
.B1(n_29),
.B2(n_21),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_111),
.Y(n_207)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_207),
.Y(n_241)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_113),
.Y(n_208)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_123),
.A2(n_29),
.B1(n_21),
.B2(n_11),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_142),
.Y(n_210)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_210),
.Y(n_253)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_158),
.Y(n_211)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_211),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_109),
.Y(n_212)
);

BUFx24_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_151),
.A2(n_11),
.B(n_16),
.C(n_15),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_L g230 ( 
.A1(n_213),
.A2(n_6),
.B(n_15),
.C(n_14),
.Y(n_230)
);

BUFx6f_ASAP7_75t_SL g214 ( 
.A(n_148),
.Y(n_214)
);

INVxp33_ASAP7_75t_L g244 ( 
.A(n_214),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_126),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_215),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_132),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_216),
.B(n_217),
.Y(n_251)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_134),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_148),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_218),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_L g220 ( 
.A1(n_159),
.A2(n_29),
.B1(n_21),
.B2(n_12),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_164),
.A2(n_29),
.B1(n_21),
.B2(n_12),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_116),
.A2(n_6),
.B1(n_15),
.B2(n_14),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_141),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_223),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_227),
.A2(n_230),
.B(n_194),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_198),
.B(n_129),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_233),
.B(n_261),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_234),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_236),
.A2(n_259),
.B1(n_220),
.B2(n_182),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_193),
.A2(n_163),
.B1(n_126),
.B2(n_144),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_237),
.A2(n_214),
.B1(n_163),
.B2(n_218),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_243),
.B(n_188),
.Y(n_287)
);

NOR2x1_ASAP7_75t_L g245 ( 
.A(n_169),
.B(n_162),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_245),
.B(n_202),
.Y(n_280)
);

CKINVDCx12_ASAP7_75t_R g258 ( 
.A(n_204),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_258),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_L g259 ( 
.A1(n_183),
.A2(n_184),
.B1(n_178),
.B2(n_191),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_205),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_200),
.B(n_108),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_263),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_200),
.B(n_160),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_215),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_264),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_240),
.A2(n_177),
.B1(n_183),
.B2(n_173),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_268),
.A2(n_272),
.B1(n_286),
.B2(n_288),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_269),
.A2(n_297),
.B1(n_267),
.B2(n_256),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_169),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_270),
.B(n_257),
.Y(n_307)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_239),
.Y(n_271)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_271),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_240),
.A2(n_243),
.B1(n_255),
.B2(n_259),
.Y(n_272)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_229),
.Y(n_273)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_273),
.Y(n_318)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_247),
.Y(n_274)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_274),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_169),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_277),
.B(n_281),
.Y(n_316)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_239),
.Y(n_278)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_278),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_227),
.A2(n_202),
.B(n_221),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_279),
.A2(n_282),
.B(n_253),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_280),
.A2(n_228),
.B(n_252),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_219),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_255),
.A2(n_174),
.B(n_179),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_283),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_186),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_284),
.B(n_287),
.Y(n_320)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_241),
.Y(n_285)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_285),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_236),
.A2(n_248),
.B1(n_266),
.B2(n_245),
.Y(n_286)
);

OAI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_230),
.A2(n_213),
.B1(n_188),
.B2(n_185),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_174),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_289),
.B(n_293),
.Y(n_326)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_225),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_290),
.A2(n_254),
.B1(n_225),
.B2(n_229),
.Y(n_324)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_241),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_291),
.B(n_299),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_265),
.B(n_199),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_248),
.B(n_181),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_295),
.B(n_296),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_251),
.A2(n_194),
.B1(n_147),
.B2(n_116),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_231),
.A2(n_232),
.B1(n_238),
.B2(n_194),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_298),
.B(n_254),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_235),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_231),
.B(n_195),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_300),
.B(n_302),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_232),
.B(n_170),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_238),
.B(n_210),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_257),
.C(n_256),
.Y(n_310)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_250),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_304),
.B(n_302),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_305),
.A2(n_311),
.B(n_279),
.Y(n_364)
);

MAJx2_ASAP7_75t_L g306 ( 
.A(n_281),
.B(n_250),
.C(n_253),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_306),
.B(n_307),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_308),
.A2(n_319),
.B1(n_329),
.B2(n_330),
.Y(n_340)
);

XNOR2x1_ASAP7_75t_L g309 ( 
.A(n_276),
.B(n_260),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_309),
.B(n_310),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_294),
.B(n_254),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_312),
.B(n_315),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_284),
.B(n_252),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_314),
.B(n_325),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_293),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_269),
.A2(n_138),
.B1(n_147),
.B2(n_171),
.Y(n_319)
);

OAI21xp33_ASAP7_75t_L g354 ( 
.A1(n_323),
.A2(n_254),
.B(n_224),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_324),
.A2(n_301),
.B1(n_273),
.B2(n_290),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_272),
.A2(n_212),
.B1(n_211),
.B2(n_247),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_297),
.A2(n_249),
.B1(n_226),
.B2(n_139),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_300),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_332),
.B(n_334),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_276),
.B(n_249),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_333),
.B(n_337),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_294),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_287),
.A2(n_228),
.B1(n_226),
.B2(n_246),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_335),
.A2(n_339),
.B1(n_296),
.B2(n_292),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_286),
.B(n_246),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_287),
.A2(n_224),
.B1(n_175),
.B2(n_135),
.Y(n_339)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_313),
.Y(n_343)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_343),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_317),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_344),
.B(n_351),
.Y(n_373)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_313),
.Y(n_346)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_346),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_335),
.B(n_287),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_347),
.Y(n_384)
);

OAI32xp33_ASAP7_75t_L g348 ( 
.A1(n_320),
.A2(n_268),
.A3(n_280),
.B1(n_277),
.B2(n_295),
.Y(n_348)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_348),
.Y(n_379)
);

OAI32xp33_ASAP7_75t_L g350 ( 
.A1(n_320),
.A2(n_289),
.A3(n_298),
.B1(n_299),
.B2(n_282),
.Y(n_350)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_350),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_317),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_352),
.A2(n_333),
.B1(n_326),
.B2(n_332),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_311),
.A2(n_275),
.B(n_292),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_353),
.A2(n_354),
.B(n_367),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_355),
.A2(n_366),
.B1(n_372),
.B2(n_330),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_312),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_356),
.B(n_365),
.Y(n_396)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_322),
.Y(n_358)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_358),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_307),
.B(n_270),
.C(n_303),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_359),
.B(n_334),
.C(n_314),
.Y(n_383)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_322),
.Y(n_360)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_360),
.Y(n_389)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_338),
.Y(n_361)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_361),
.Y(n_393)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_338),
.Y(n_362)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_362),
.Y(n_399)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_325),
.Y(n_363)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_363),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_364),
.B(n_323),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_326),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_328),
.A2(n_271),
.B1(n_291),
.B2(n_285),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_339),
.B(n_304),
.Y(n_367)
);

BUFx5_ASAP7_75t_L g368 ( 
.A(n_318),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_368),
.Y(n_381)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_321),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_369),
.Y(n_392)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_321),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_371),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_328),
.A2(n_327),
.B1(n_337),
.B2(n_315),
.Y(n_372)
);

OA21x2_ASAP7_75t_L g374 ( 
.A1(n_357),
.A2(n_327),
.B(n_305),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_374),
.B(n_402),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_363),
.B(n_331),
.Y(n_375)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_375),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_341),
.B(n_331),
.Y(n_377)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_377),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_383),
.B(n_350),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g386 ( 
.A(n_342),
.B(n_306),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_386),
.B(n_403),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_370),
.B(n_316),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_387),
.B(n_390),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_388),
.A2(n_391),
.B1(n_397),
.B2(n_346),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_349),
.B(n_316),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_352),
.A2(n_336),
.B1(n_308),
.B2(n_319),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_349),
.B(n_366),
.Y(n_394)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_394),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_395),
.A2(n_273),
.B1(n_274),
.B2(n_242),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_347),
.A2(n_310),
.B1(n_329),
.B2(n_309),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_372),
.B(n_278),
.Y(n_400)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_400),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_357),
.B(n_367),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_345),
.B(n_309),
.C(n_306),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_404),
.B(n_359),
.C(n_345),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_387),
.B(n_348),
.Y(n_405)
);

CKINVDCx14_ASAP7_75t_R g449 ( 
.A(n_405),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_373),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_406),
.Y(n_446)
);

INVx13_ASAP7_75t_L g409 ( 
.A(n_381),
.Y(n_409)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_409),
.Y(n_436)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_401),
.Y(n_410)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_410),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_396),
.B(n_360),
.Y(n_411)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_411),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_413),
.B(n_403),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_383),
.B(n_342),
.C(n_364),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_414),
.B(n_419),
.C(n_427),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_379),
.A2(n_340),
.B1(n_353),
.B2(n_367),
.Y(n_415)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_415),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_379),
.A2(n_382),
.B1(n_395),
.B2(n_340),
.Y(n_416)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_416),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_382),
.B(n_301),
.Y(n_418)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_418),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_380),
.A2(n_347),
.B(n_355),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_420),
.A2(n_374),
.B(n_389),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_390),
.B(n_343),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_421),
.A2(n_429),
.B1(n_433),
.B2(n_399),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_380),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_422),
.A2(n_430),
.B(n_399),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_423),
.A2(n_431),
.B1(n_432),
.B2(n_400),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_404),
.B(n_371),
.C(n_369),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_386),
.B(n_362),
.C(n_361),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_428),
.B(n_398),
.C(n_392),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_377),
.B(n_358),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_402),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_391),
.A2(n_368),
.B1(n_318),
.B2(n_290),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_401),
.B(n_180),
.Y(n_433)
);

XNOR2x1_ASAP7_75t_L g438 ( 
.A(n_426),
.B(n_397),
.Y(n_438)
);

XNOR2x1_ASAP7_75t_L g459 ( 
.A(n_438),
.B(n_455),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_440),
.B(n_454),
.C(n_413),
.Y(n_465)
);

AOI21x1_ASAP7_75t_SL g441 ( 
.A1(n_407),
.A2(n_374),
.B(n_384),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g458 ( 
.A(n_441),
.B(n_447),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_442),
.A2(n_444),
.B1(n_425),
.B2(n_424),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_423),
.A2(n_394),
.B1(n_384),
.B2(n_375),
.Y(n_443)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_443),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_425),
.A2(n_374),
.B1(n_388),
.B2(n_398),
.Y(n_444)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_445),
.Y(n_460)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_448),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_427),
.B(n_393),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_452),
.B(n_453),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_414),
.B(n_392),
.C(n_393),
.Y(n_454)
);

XNOR2x1_ASAP7_75t_L g455 ( 
.A(n_426),
.B(n_381),
.Y(n_455)
);

FAx1_ASAP7_75t_SL g456 ( 
.A(n_419),
.B(n_389),
.CI(n_385),
.CON(n_456),
.SN(n_456)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_456),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_454),
.B(n_417),
.Y(n_457)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_457),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_461),
.A2(n_475),
.B1(n_435),
.B2(n_378),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_452),
.B(n_428),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_463),
.B(n_465),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_449),
.A2(n_406),
.B1(n_431),
.B2(n_411),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_464),
.A2(n_467),
.B1(n_473),
.B2(n_422),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_437),
.A2(n_407),
.B1(n_424),
.B2(n_408),
.Y(n_467)
);

FAx1_ASAP7_75t_SL g470 ( 
.A(n_441),
.B(n_417),
.CI(n_430),
.CON(n_470),
.SN(n_470)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_470),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_448),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_471),
.B(n_472),
.Y(n_490)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_434),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_450),
.A2(n_439),
.B1(n_412),
.B2(n_408),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_412),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_474),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_442),
.A2(n_444),
.B1(n_443),
.B2(n_420),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_476),
.B(n_477),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_438),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_469),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_478),
.B(n_481),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_465),
.B(n_451),
.C(n_440),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_480),
.B(n_482),
.C(n_484),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_460),
.A2(n_432),
.B1(n_446),
.B2(n_436),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_462),
.B(n_451),
.C(n_463),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_466),
.A2(n_446),
.B1(n_436),
.B2(n_410),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_483),
.B(n_491),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_462),
.B(n_453),
.C(n_456),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_459),
.B(n_455),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_486),
.B(n_489),
.C(n_492),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_470),
.B(n_447),
.Y(n_488)
);

CKINVDCx14_ASAP7_75t_R g494 ( 
.A(n_488),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_475),
.B(n_385),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_461),
.B(n_378),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_487),
.A2(n_458),
.B(n_468),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_495),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_485),
.B(n_470),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_497),
.B(n_498),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_493),
.B(n_458),
.Y(n_498)
);

OAI21x1_ASAP7_75t_SL g499 ( 
.A1(n_488),
.A2(n_467),
.B(n_466),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_499),
.A2(n_242),
.B1(n_135),
.B2(n_133),
.Y(n_517)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_490),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_501),
.B(n_504),
.Y(n_513)
);

AO21x1_ASAP7_75t_L g502 ( 
.A1(n_489),
.A2(n_376),
.B(n_409),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_502),
.B(n_486),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_479),
.B(n_376),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_492),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_505),
.B(n_507),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_484),
.B(n_482),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_509),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_500),
.B(n_480),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_511),
.B(n_517),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_498),
.A2(n_477),
.B1(n_201),
.B2(n_196),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_515),
.B(n_516),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_500),
.B(n_242),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_507),
.A2(n_204),
.B(n_153),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_518),
.A2(n_519),
.B(n_502),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_494),
.A2(n_133),
.B1(n_244),
.B2(n_120),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_496),
.B(n_119),
.Y(n_520)
);

CKINVDCx14_ASAP7_75t_R g521 ( 
.A(n_520),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_522),
.B(n_509),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_512),
.A2(n_496),
.B(n_506),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_SL g529 ( 
.A1(n_524),
.A2(n_513),
.B(n_508),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_514),
.B(n_508),
.C(n_503),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_525),
.B(n_510),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_528),
.B(n_530),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_529),
.A2(n_531),
.B(n_526),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_527),
.A2(n_517),
.B(n_519),
.Y(n_531)
);

AOI21xp33_ASAP7_75t_L g532 ( 
.A1(n_530),
.A2(n_527),
.B(n_523),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_SL g536 ( 
.A1(n_532),
.A2(n_533),
.B(n_136),
.Y(n_536)
);

OAI311xp33_ASAP7_75t_L g535 ( 
.A1(n_534),
.A2(n_521),
.A3(n_244),
.B1(n_136),
.C1(n_3),
.Y(n_535)
);

AOI322xp5_ASAP7_75t_L g537 ( 
.A1(n_535),
.A2(n_536),
.A3(n_7),
.B1(n_15),
.B2(n_14),
.C1(n_3),
.C2(n_16),
.Y(n_537)
);

OAI21xp33_ASAP7_75t_SL g538 ( 
.A1(n_537),
.A2(n_16),
.B(n_1),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_538),
.A2(n_0),
.B(n_1),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_539),
.B(n_0),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_540),
.A2(n_0),
.B(n_2),
.Y(n_541)
);


endmodule