module fake_jpeg_3497_n_485 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_485);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_485;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_49),
.Y(n_143)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_51),
.Y(n_130)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_18),
.B(n_20),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_53),
.B(n_71),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_55),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_24),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_62),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g140 ( 
.A(n_58),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_70),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_41),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_24),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_78),
.Y(n_102)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_40),
.B(n_0),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_82),
.Y(n_121)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_84),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_40),
.B(n_0),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_28),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_28),
.B(n_14),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_86),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_35),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_22),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_94),
.Y(n_114)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_35),
.B(n_16),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_96),
.B(n_14),
.Y(n_145)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_26),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_80),
.A2(n_27),
.B1(n_48),
.B2(n_19),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_101),
.A2(n_79),
.B1(n_74),
.B2(n_73),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_75),
.A2(n_29),
.B1(n_45),
.B2(n_43),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_104),
.A2(n_113),
.B1(n_128),
.B2(n_132),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_77),
.A2(n_29),
.B1(n_45),
.B2(n_43),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_58),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_82),
.A2(n_26),
.B1(n_38),
.B2(n_36),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_118),
.A2(n_124),
.B1(n_125),
.B2(n_59),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_25),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_142),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_54),
.A2(n_19),
.B1(n_38),
.B2(n_36),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_50),
.A2(n_23),
.B1(n_25),
.B2(n_48),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_51),
.A2(n_29),
.B1(n_23),
.B2(n_30),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_55),
.A2(n_22),
.B1(n_1),
.B2(n_2),
.Y(n_132)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_52),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_137),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_60),
.B(n_16),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_61),
.B(n_16),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_150),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_145),
.B(n_0),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_64),
.B(n_13),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_83),
.A2(n_13),
.B1(n_2),
.B2(n_3),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_5),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_87),
.B(n_12),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_153),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_90),
.B(n_12),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_155),
.B(n_156),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_95),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_157),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_107),
.B(n_91),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_158),
.B(n_177),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_161),
.B(n_184),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_162),
.B(n_181),
.Y(n_221)
);

AO22x1_ASAP7_75t_SL g163 ( 
.A1(n_118),
.A2(n_57),
.B1(n_88),
.B2(n_89),
.Y(n_163)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_163),
.Y(n_215)
);

OA22x2_ASAP7_75t_L g232 ( 
.A1(n_164),
.A2(n_183),
.B1(n_120),
.B2(n_117),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_165),
.Y(n_234)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_168),
.Y(n_250)
);

FAx1_ASAP7_75t_SL g169 ( 
.A(n_121),
.B(n_72),
.CI(n_69),
.CON(n_169),
.SN(n_169)
);

BUFx24_ASAP7_75t_SL g237 ( 
.A(n_169),
.Y(n_237)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_170),
.Y(n_220)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_171),
.Y(n_233)
);

O2A1O1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_125),
.A2(n_67),
.B(n_65),
.C(n_63),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_172),
.A2(n_163),
.B(n_131),
.C(n_127),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_109),
.A2(n_68),
.B1(n_3),
.B2(n_4),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_173),
.A2(n_202),
.B1(n_151),
.B2(n_183),
.Y(n_218)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_174),
.Y(n_225)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_116),
.Y(n_175)
);

INVxp67_ASAP7_75t_SL g252 ( 
.A(n_175),
.Y(n_252)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_99),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_102),
.B(n_2),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_178),
.B(n_185),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g180 ( 
.A(n_123),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_180),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_114),
.Y(n_181)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_116),
.Y(n_182)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_182),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_149),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_98),
.B(n_5),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_110),
.Y(n_186)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_186),
.Y(n_238)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_139),
.Y(n_187)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_187),
.Y(n_243)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_139),
.Y(n_188)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_188),
.Y(n_246)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_110),
.Y(n_189)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_189),
.Y(n_254)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_190),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g191 ( 
.A(n_130),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_191),
.B(n_192),
.Y(n_239)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_149),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_195),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_145),
.B(n_6),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_194),
.B(n_203),
.Y(n_231)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_106),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_103),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_196),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_121),
.A2(n_153),
.B1(n_109),
.B2(n_148),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_197),
.Y(n_229)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_111),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_206),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_129),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_199),
.B(n_201),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_117),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_200),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_100),
.B(n_6),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_124),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_100),
.B(n_7),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_111),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_204),
.B(n_205),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_129),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_105),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_148),
.A2(n_9),
.B(n_11),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_207),
.A2(n_106),
.B(n_108),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_105),
.B(n_11),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_11),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_130),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_209),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_119),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_213),
.B(n_147),
.C(n_11),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_214),
.B(n_179),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_217),
.A2(n_172),
.B1(n_180),
.B2(n_198),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_218),
.A2(n_236),
.B1(n_184),
.B2(n_202),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_161),
.A2(n_119),
.B1(n_131),
.B2(n_120),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_228),
.A2(n_240),
.B1(n_174),
.B2(n_196),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_232),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_167),
.B(n_134),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_241),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_169),
.A2(n_146),
.B1(n_108),
.B2(n_134),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_169),
.A2(n_136),
.B1(n_127),
.B2(n_146),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_160),
.B(n_136),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_244),
.A2(n_166),
.B(n_140),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_159),
.B(n_141),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_251),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_163),
.B(n_141),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_207),
.B(n_173),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_218),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_171),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_179),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_216),
.B(n_193),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_258),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_259),
.B(n_266),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_227),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_260),
.B(n_262),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_212),
.B(n_175),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_261),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_227),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_263),
.A2(n_279),
.B1(n_294),
.B2(n_295),
.Y(n_301)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_264),
.Y(n_304)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_267),
.Y(n_312)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_268),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_210),
.B(n_206),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_269),
.B(n_273),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_270),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_271),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_239),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_272),
.B(n_276),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_210),
.B(n_247),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_225),
.Y(n_274)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_274),
.Y(n_335)
);

NOR2x1_ASAP7_75t_L g275 ( 
.A(n_213),
.B(n_187),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_275),
.A2(n_290),
.B(n_296),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_227),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_236),
.A2(n_166),
.B1(n_186),
.B2(n_189),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_277),
.A2(n_284),
.B(n_293),
.Y(n_313)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_225),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_278),
.B(n_282),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_215),
.A2(n_165),
.B1(n_200),
.B2(n_168),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_280),
.A2(n_281),
.B1(n_219),
.B2(n_223),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_215),
.A2(n_170),
.B1(n_133),
.B2(n_182),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_241),
.B(n_191),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_235),
.B(n_214),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_297),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_229),
.A2(n_140),
.B1(n_133),
.B2(n_195),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_226),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_285),
.A2(n_287),
.B1(n_288),
.B2(n_291),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_230),
.B(n_191),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_286),
.Y(n_325)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_225),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_243),
.Y(n_288)
);

NOR2x1_ASAP7_75t_L g290 ( 
.A(n_224),
.B(n_180),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_243),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_226),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_292),
.Y(n_331)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_226),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_249),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_240),
.A2(n_126),
.B1(n_147),
.B2(n_137),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_221),
.B(n_126),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_253),
.B(n_12),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_298),
.B(n_238),
.Y(n_329)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_250),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_299),
.A2(n_223),
.B1(n_219),
.B2(n_220),
.Y(n_303)
);

OAI32xp33_ASAP7_75t_L g300 ( 
.A1(n_266),
.A2(n_229),
.A3(n_224),
.B1(n_237),
.B2(n_251),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_300),
.Y(n_339)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_303),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_271),
.A2(n_244),
.B(n_217),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_307),
.A2(n_314),
.B(n_317),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_308),
.A2(n_318),
.B1(n_285),
.B2(n_295),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_289),
.A2(n_224),
.B1(n_228),
.B2(n_245),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_309),
.A2(n_311),
.B1(n_315),
.B2(n_328),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_289),
.A2(n_256),
.B1(n_232),
.B2(n_231),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_290),
.A2(n_265),
.B(n_264),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_265),
.A2(n_232),
.B1(n_231),
.B2(n_221),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_290),
.A2(n_248),
.B(n_252),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_273),
.A2(n_248),
.B(n_242),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_263),
.A2(n_232),
.B1(n_220),
.B2(n_233),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_323),
.A2(n_326),
.B1(n_260),
.B2(n_262),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_275),
.B(n_255),
.C(n_211),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_324),
.B(n_332),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_277),
.A2(n_250),
.B1(n_234),
.B2(n_255),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_279),
.A2(n_234),
.B1(n_238),
.B2(n_254),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_329),
.B(n_268),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_257),
.B(n_211),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_330),
.B(n_292),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_275),
.B(n_222),
.C(n_254),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_298),
.A2(n_222),
.B1(n_242),
.B2(n_257),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_333),
.A2(n_293),
.B1(n_280),
.B2(n_267),
.Y(n_354)
);

A2O1A1Ixp33_ASAP7_75t_L g340 ( 
.A1(n_302),
.A2(n_283),
.B(n_259),
.C(n_282),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_340),
.B(n_367),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_341),
.Y(n_388)
);

OAI22x1_ASAP7_75t_L g342 ( 
.A1(n_319),
.A2(n_284),
.B1(n_296),
.B2(n_281),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g389 ( 
.A1(n_342),
.A2(n_345),
.B1(n_363),
.B2(n_365),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_294),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_343),
.B(n_346),
.C(n_306),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_316),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_344),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_322),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_306),
.B(n_297),
.Y(n_346)
);

BUFx5_ASAP7_75t_L g349 ( 
.A(n_325),
.Y(n_349)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_349),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_351),
.A2(n_354),
.B1(n_304),
.B2(n_333),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_352),
.B(n_358),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_276),
.Y(n_353)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_353),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_323),
.A2(n_301),
.B1(n_311),
.B2(n_307),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_355),
.A2(n_351),
.B1(n_301),
.B2(n_309),
.Y(n_377)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_312),
.Y(n_356)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_356),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_327),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_357),
.B(n_360),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_334),
.A2(n_269),
.B1(n_288),
.B2(n_291),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_359),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_325),
.B(n_274),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_312),
.Y(n_361)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_361),
.Y(n_375)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_321),
.Y(n_362)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_362),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_318),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_321),
.Y(n_364)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_364),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_320),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_335),
.Y(n_366)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_366),
.Y(n_384)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_335),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_303),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_368),
.B(n_369),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_331),
.B(n_278),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_370),
.B(n_374),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_343),
.B(n_324),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_377),
.A2(n_391),
.B1(n_395),
.B2(n_393),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_353),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_378),
.B(n_396),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_346),
.B(n_332),
.C(n_310),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_379),
.B(n_387),
.C(n_390),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_338),
.B(n_314),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_385),
.B(n_367),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_338),
.B(n_310),
.C(n_305),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_352),
.B(n_304),
.C(n_329),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_355),
.A2(n_315),
.B1(n_334),
.B2(n_319),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_392),
.A2(n_348),
.B1(n_363),
.B2(n_368),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_339),
.A2(n_319),
.B1(n_313),
.B2(n_328),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_345),
.B(n_337),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_380),
.A2(n_365),
.B1(n_339),
.B2(n_344),
.Y(n_398)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_398),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_370),
.B(n_340),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_409),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_401),
.A2(n_403),
.B1(n_404),
.B2(n_392),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_387),
.A2(n_347),
.B(n_337),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_376),
.Y(n_405)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_405),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_383),
.B(n_369),
.Y(n_406)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_406),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_383),
.B(n_371),
.Y(n_407)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_407),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_393),
.A2(n_347),
.B(n_359),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_408),
.A2(n_416),
.B(n_382),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_379),
.B(n_374),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_385),
.B(n_300),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_410),
.B(n_411),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_390),
.B(n_317),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_394),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_412),
.B(n_417),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_389),
.Y(n_413)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_413),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_394),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_414),
.A2(n_413),
.B1(n_395),
.B2(n_342),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_373),
.B(n_350),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_415),
.B(n_418),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_386),
.A2(n_350),
.B(n_313),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_388),
.A2(n_336),
.B(n_349),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_386),
.Y(n_419)
);

BUFx12_ASAP7_75t_L g427 ( 
.A(n_419),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_L g450 ( 
.A1(n_421),
.A2(n_431),
.B1(n_429),
.B2(n_423),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_401),
.A2(n_388),
.B1(n_376),
.B2(n_384),
.Y(n_422)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_422),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_402),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_424),
.B(n_430),
.Y(n_451)
);

AO21x2_ASAP7_75t_L g428 ( 
.A1(n_408),
.A2(n_377),
.B(n_391),
.Y(n_428)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_428),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_416),
.A2(n_326),
.B(n_381),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_409),
.B(n_373),
.C(n_366),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_433),
.B(n_399),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_435),
.B(n_414),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_420),
.B(n_415),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_439),
.B(n_440),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_436),
.B(n_400),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_442),
.B(n_447),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_443),
.B(n_445),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_433),
.B(n_418),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_444),
.B(n_446),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_432),
.B(n_397),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_426),
.B(n_397),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_426),
.B(n_399),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_425),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_448),
.A2(n_449),
.B1(n_450),
.B2(n_430),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_435),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_451),
.A2(n_437),
.B(n_431),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_453),
.B(n_454),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_446),
.B(n_434),
.C(n_437),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_458),
.A2(n_463),
.B1(n_428),
.B2(n_462),
.Y(n_470)
);

BUFx24_ASAP7_75t_SL g459 ( 
.A(n_450),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_459),
.B(n_419),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_434),
.C(n_429),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_460),
.B(n_462),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_411),
.C(n_410),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_461),
.B(n_463),
.C(n_441),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_438),
.B(n_428),
.C(n_427),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_442),
.B(n_428),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_465),
.B(n_470),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_456),
.B(n_427),
.C(n_375),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_466),
.B(n_468),
.Y(n_474)
);

NOR3xp33_ASAP7_75t_L g469 ( 
.A(n_452),
.B(n_427),
.C(n_372),
.Y(n_469)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_469),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_455),
.B(n_460),
.C(n_454),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_471),
.B(n_364),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_464),
.B(n_457),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_473),
.B(n_475),
.Y(n_478)
);

AOI22xp33_ASAP7_75t_L g477 ( 
.A1(n_476),
.A2(n_464),
.B1(n_467),
.B2(n_361),
.Y(n_477)
);

O2A1O1Ixp33_ASAP7_75t_SL g480 ( 
.A1(n_477),
.A2(n_474),
.B(n_472),
.C(n_287),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_472),
.A2(n_356),
.B(n_362),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_479),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_480),
.Y(n_482)
);

AO21x1_ASAP7_75t_L g483 ( 
.A1(n_482),
.A2(n_481),
.B(n_478),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_483),
.B(n_299),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_484),
.B(n_308),
.Y(n_485)
);


endmodule