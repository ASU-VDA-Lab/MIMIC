module fake_jpeg_9289_n_274 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_274);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_4),
.B(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_43),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_34),
.B(n_26),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_50),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_21),
.C(n_26),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_53),
.B(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_21),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_20),
.B1(n_23),
.B2(n_34),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_59),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_23),
.B1(n_32),
.B2(n_22),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_10),
.B1(n_16),
.B2(n_2),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_22),
.B1(n_29),
.B2(n_17),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_32),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_31),
.Y(n_61)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_31),
.Y(n_64)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_10),
.Y(n_65)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_67),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_29),
.B1(n_18),
.B2(n_33),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_68),
.A2(n_57),
.B1(n_60),
.B2(n_49),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_29),
.B1(n_33),
.B2(n_27),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_69),
.A2(n_73),
.B1(n_83),
.B2(n_66),
.Y(n_100)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_72),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_71),
.B(n_80),
.Y(n_96)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_66),
.A2(n_18),
.B1(n_19),
.B2(n_25),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_78),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_66),
.A2(n_25),
.B1(n_19),
.B2(n_27),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_76),
.A2(n_85),
.B1(n_41),
.B2(n_12),
.Y(n_106)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_45),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_62),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_88),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_45),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_89),
.B(n_50),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_91),
.B(n_95),
.Y(n_117)
);

AO22x1_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_62),
.B1(n_49),
.B2(n_60),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_37),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_80),
.B(n_47),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_59),
.C(n_48),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_102),
.C(n_108),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_87),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_101),
.Y(n_119)
);

BUFx8_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_85),
.B1(n_90),
.B2(n_88),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_87),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_82),
.C(n_89),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_110),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_105),
.A2(n_74),
.B1(n_37),
.B2(n_86),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_106),
.A2(n_113),
.B1(n_74),
.B2(n_12),
.Y(n_134)
);

NOR2x1p5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_35),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_42),
.B(n_44),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_35),
.C(n_37),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_SL g109 ( 
.A(n_77),
.B(n_41),
.C(n_44),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_109),
.A2(n_107),
.B(n_108),
.Y(n_128)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_90),
.B(n_11),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_111),
.B(n_12),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_73),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_114),
.Y(n_130)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_122),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_125),
.B1(n_103),
.B2(n_74),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_120),
.A2(n_124),
.B(n_128),
.Y(n_148)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_107),
.A2(n_84),
.B1(n_78),
.B2(n_79),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_132),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_101),
.Y(n_127)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_84),
.Y(n_129)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_131),
.B(n_9),
.Y(n_143)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

INVx6_ASAP7_75t_SL g151 ( 
.A(n_133),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_SL g147 ( 
.A(n_134),
.B(n_92),
.C(n_7),
.Y(n_147)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_137),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_110),
.B1(n_113),
.B2(n_114),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_91),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_139),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_111),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_129),
.C(n_128),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_145),
.C(n_160),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_143),
.B(n_164),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_97),
.C(n_120),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_92),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_146),
.A2(n_149),
.B(n_156),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_147),
.A2(n_161),
.B1(n_116),
.B2(n_135),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_119),
.A2(n_95),
.B(n_112),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_121),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_152),
.B(n_154),
.Y(n_175)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_155),
.Y(n_188)
);

NOR4xp25_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_103),
.C(n_16),
.D(n_2),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_159),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_100),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_118),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_44),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_124),
.A2(n_99),
.B(n_44),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_138),
.B(n_11),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_55),
.C(n_54),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_165),
.B(n_142),
.C(n_145),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_186),
.C(n_151),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_141),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_168),
.B(n_172),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_169),
.A2(n_179),
.B1(n_147),
.B2(n_161),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_137),
.Y(n_170)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_157),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_181),
.Y(n_202)
);

AO22x1_ASAP7_75t_SL g174 ( 
.A1(n_146),
.A2(n_136),
.B1(n_126),
.B2(n_117),
.Y(n_174)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_122),
.C(n_115),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_178),
.C(n_52),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_139),
.C(n_132),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_162),
.A2(n_132),
.B1(n_131),
.B2(n_99),
.Y(n_179)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_140),
.A2(n_86),
.B1(n_55),
.B2(n_54),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_182),
.A2(n_183),
.B1(n_159),
.B2(n_158),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_140),
.A2(n_54),
.B1(n_52),
.B2(n_44),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_0),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_185),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_148),
.B(n_52),
.C(n_42),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_151),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_200),
.C(n_201),
.Y(n_212)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_174),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_199),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_171),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_194),
.B(n_196),
.Y(n_219)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_168),
.B(n_164),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_177),
.B(n_149),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_178),
.Y(n_215)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_198),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_171),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_160),
.C(n_165),
.Y(n_201)
);

AND2x6_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_146),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_206),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_188),
.A2(n_152),
.B1(n_155),
.B2(n_163),
.Y(n_204)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

NOR3xp33_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_156),
.C(n_143),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_167),
.C(n_181),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_210),
.C(n_217),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_208),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_192),
.A2(n_184),
.B1(n_172),
.B2(n_177),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_218),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_186),
.C(n_176),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_175),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_207),
.C(n_204),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_224),
.C(n_195),
.Y(n_237)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_223),
.B(n_182),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_180),
.C(n_184),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_216),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_226),
.Y(n_240)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_219),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_190),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_232),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_214),
.A2(n_191),
.B1(n_205),
.B2(n_203),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_230),
.A2(n_229),
.B1(n_236),
.B2(n_226),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_220),
.A2(n_205),
.B(n_193),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_235),
.Y(n_244)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_224),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_233),
.A2(n_236),
.B1(n_8),
.B2(n_16),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_185),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_218),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_215),
.C(n_179),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_212),
.C(n_217),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_239),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_212),
.C(n_221),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_243),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_183),
.C(n_187),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_245),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_229),
.A2(n_187),
.B1(n_8),
.B2(n_3),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_235),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_228),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_42),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_252),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_231),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_255),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_238),
.A2(n_230),
.B1(n_228),
.B2(n_0),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_254),
.A2(n_6),
.B1(n_13),
.B2(n_4),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_7),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_249),
.A2(n_240),
.B(n_7),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_251),
.C(n_254),
.Y(n_262)
);

OAI21x1_ASAP7_75t_L g258 ( 
.A1(n_248),
.A2(n_6),
.B(n_13),
.Y(n_258)
);

NAND3xp33_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_13),
.C(n_11),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_260),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_265),
.Y(n_269)
);

AO21x2_ASAP7_75t_L g267 ( 
.A1(n_264),
.A2(n_5),
.B(n_1),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_261),
.B(n_248),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_256),
.A2(n_250),
.B1(n_5),
.B2(n_9),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_266),
.B(n_261),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_267),
.B(n_268),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_269),
.A2(n_263),
.B(n_264),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_270),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_272),
.A2(n_271),
.B(n_1),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_0),
.C(n_42),
.Y(n_274)
);


endmodule