module fake_jpeg_19140_n_176 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_29),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_37),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx24_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_29),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_24),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_23),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_47),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_30),
.B1(n_21),
.B2(n_20),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_33),
.B(n_18),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_23),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_52),
.B(n_35),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_30),
.B1(n_21),
.B2(n_22),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_40),
.B1(n_38),
.B2(n_36),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_21),
.B1(n_18),
.B2(n_20),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_31),
.B1(n_38),
.B2(n_22),
.Y(n_67)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_40),
.B1(n_36),
.B2(n_31),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_60),
.A2(n_42),
.B1(n_55),
.B2(n_50),
.Y(n_88)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_67),
.B1(n_75),
.B2(n_49),
.Y(n_86)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_19),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_69),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_43),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_66),
.B(n_70),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_35),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_27),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_42),
.Y(n_78)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_44),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_45),
.A2(n_39),
.B1(n_38),
.B2(n_36),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_19),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_76),
.B(n_28),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_50),
.A2(n_36),
.B(n_34),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_77),
.A2(n_36),
.B(n_49),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_82),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_64),
.B1(n_62),
.B2(n_71),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_81),
.B(n_65),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_55),
.B(n_56),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_60),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_26),
.B(n_25),
.C(n_16),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_93),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_96),
.Y(n_102)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_74),
.B1(n_59),
.B2(n_60),
.Y(n_108)
);

A2O1A1O1Ixp25_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_15),
.B(n_24),
.C(n_23),
.D(n_27),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_94),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_24),
.Y(n_93)
);

BUFx24_ASAP7_75t_SL g94 ( 
.A(n_66),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_28),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_68),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_25),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_108),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_89),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_101),
.B(n_110),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_103),
.B(n_113),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_92),
.A2(n_68),
.B1(n_16),
.B2(n_26),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_115),
.Y(n_124)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_69),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_90),
.A2(n_68),
.B1(n_60),
.B2(n_74),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_112),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_70),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_73),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_114),
.B(n_74),
.Y(n_126)
);

A2O1A1O1Ixp25_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_83),
.B(n_78),
.C(n_80),
.D(n_91),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_116),
.A2(n_118),
.B(n_123),
.Y(n_134)
);

A2O1A1O1Ixp25_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_82),
.B(n_85),
.C(n_93),
.D(n_84),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_98),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_95),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_131),
.Y(n_135)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_103),
.B(n_79),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_127),
.A2(n_79),
.B(n_104),
.Y(n_133)
);

NOR3xp33_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_109),
.C(n_107),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_98),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_130),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_100),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_102),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_132),
.A2(n_119),
.B(n_122),
.Y(n_147)
);

AOI321xp33_ASAP7_75t_L g148 ( 
.A1(n_133),
.A2(n_125),
.A3(n_128),
.B1(n_13),
.B2(n_11),
.C(n_10),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_102),
.B1(n_106),
.B2(n_99),
.Y(n_136)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_121),
.A2(n_115),
.B(n_108),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_139),
.A2(n_118),
.B(n_116),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_115),
.C(n_85),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_143),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_77),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_142),
.B(n_140),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_88),
.C(n_60),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_151),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_124),
.B(n_121),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_145),
.A2(n_146),
.B(n_137),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_147),
.A2(n_135),
.B(n_139),
.Y(n_157)
);

AOI31xp67_ASAP7_75t_L g156 ( 
.A1(n_148),
.A2(n_137),
.A3(n_138),
.B(n_11),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_128),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_132),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_150),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_157),
.Y(n_161)
);

AOI31xp33_ASAP7_75t_L g162 ( 
.A1(n_154),
.A2(n_156),
.A3(n_149),
.B(n_3),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_141),
.Y(n_155)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_158),
.A2(n_143),
.B1(n_155),
.B2(n_151),
.Y(n_164)
);

XNOR2x1_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_146),
.Y(n_160)
);

O2A1O1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_160),
.A2(n_162),
.B(n_165),
.C(n_7),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_164),
.B(n_8),
.Y(n_169)
);

MAJx2_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_2),
.C(n_3),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_163),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_168),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_8),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_7),
.C(n_8),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_160),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_170),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_171),
.A2(n_165),
.B(n_166),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_172),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_174),
.Y(n_176)
);


endmodule