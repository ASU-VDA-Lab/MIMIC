module real_jpeg_24272_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_288;
wire n_166;
wire n_286;
wire n_176;
wire n_292;
wire n_249;
wire n_215;
wire n_221;
wire n_300;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_258;
wire n_205;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_216;
wire n_295;
wire n_202;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_213;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_2),
.A2(n_23),
.B1(n_36),
.B2(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_2),
.A2(n_31),
.B1(n_33),
.B2(n_60),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_2),
.A2(n_53),
.B1(n_55),
.B2(n_60),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_2),
.A2(n_60),
.B1(n_73),
.B2(n_74),
.Y(n_194)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_3),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_4),
.A2(n_15),
.B(n_301),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_4),
.B(n_302),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_7),
.A2(n_21),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_7),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_7),
.A2(n_35),
.B1(n_53),
.B2(n_55),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_7),
.A2(n_35),
.B1(n_73),
.B2(n_74),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_8),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_8),
.A2(n_25),
.B1(n_31),
.B2(n_33),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_8),
.A2(n_25),
.B1(n_53),
.B2(n_55),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_8),
.A2(n_25),
.B1(n_73),
.B2(n_74),
.Y(n_129)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_9),
.A2(n_23),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_43),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_10),
.A2(n_43),
.B1(n_53),
.B2(n_55),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_10),
.A2(n_31),
.B1(n_33),
.B2(n_43),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_10),
.A2(n_43),
.B1(n_73),
.B2(n_74),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_10),
.B(n_29),
.C(n_33),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_10),
.B(n_30),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_10),
.B(n_50),
.C(n_53),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_10),
.B(n_70),
.C(n_73),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_10),
.B(n_87),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_10),
.B(n_104),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_10),
.B(n_63),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_12),
.Y(n_302)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_13),
.Y(n_85)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_13),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_13),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_192)
);

AOI21xp33_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_294),
.B(n_298),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_76),
.B(n_293),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_37),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_18),
.B(n_37),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_18),
.B(n_295),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_18),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_26),
.B1(n_30),
.B2(n_34),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_20),
.A2(n_40),
.B(n_41),
.Y(n_39)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_26),
.A2(n_30),
.B1(n_42),
.B2(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_26),
.B(n_30),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

AO22x1_ASAP7_75t_SL g30 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_30)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g33 ( 
.A(n_31),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_31),
.A2(n_33),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

CKINVDCx6p67_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_33),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_34),
.B(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_36),
.B(n_190),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_38),
.B(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_38),
.B(n_291),
.Y(n_292)
);

FAx1_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_44),
.CI(n_56),
.CON(n_38),
.SN(n_38)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_40),
.A2(n_41),
.B(n_59),
.Y(n_113)
);

INVxp33_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_48),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_52),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_47),
.A2(n_52),
.B(n_170),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_48),
.A2(n_63),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_48),
.B(n_109),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

OA22x2_ASAP7_75t_SL g52 ( 
.A1(n_50),
.A2(n_51),
.B1(n_53),
.B2(n_55),
.Y(n_52)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_52),
.A2(n_118),
.B(n_119),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_52),
.A2(n_108),
.B(n_119),
.Y(n_136)
);

INVx5_ASAP7_75t_SL g55 ( 
.A(n_53),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_55),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_53),
.B(n_236),
.Y(n_235)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_61),
.C(n_64),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_SL g126 ( 
.A(n_57),
.B(n_127),
.C(n_135),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_57),
.A2(n_146),
.B1(n_148),
.B2(n_149),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_57),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_57),
.A2(n_135),
.B1(n_136),
.B2(n_149),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_57),
.A2(n_106),
.B1(n_149),
.B2(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_57),
.B(n_106),
.C(n_187),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_61),
.A2(n_64),
.B1(n_116),
.B2(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_61),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_64),
.A2(n_116),
.B1(n_117),
.B2(n_120),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_64),
.B(n_112),
.C(n_117),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_75),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_66),
.B(n_94),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_72),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_68),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_68),
.A2(n_94),
.B1(n_104),
.B2(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_72),
.A2(n_92),
.B(n_93),
.Y(n_91)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_72),
.A2(n_93),
.B(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_73),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_73),
.B(n_241),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_290),
.B(n_292),
.Y(n_76)
);

OAI211xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_137),
.B(n_151),
.C(n_289),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_121),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_79),
.B(n_121),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_99),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_80),
.B(n_101),
.C(n_110),
.Y(n_139)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_90),
.B(n_95),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_81),
.A2(n_95),
.B1(n_96),
.B2(n_124),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_81),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_81),
.A2(n_91),
.B1(n_124),
.B2(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_89),
.Y(n_81)
);

INVxp33_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_83),
.B(n_195),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_84),
.A2(n_89),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_84),
.B(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_84),
.Y(n_193)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_88),
.A2(n_129),
.B(n_164),
.Y(n_163)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_88),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_90),
.B(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_91),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_97),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_110),
.B2(n_111),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_101),
.A2(n_102),
.B(n_106),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_106),
.Y(n_101)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_106),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_106),
.B(n_207),
.C(n_209),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_106),
.A2(n_197),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_109),
.Y(n_170)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_112),
.A2(n_113),
.B1(n_145),
.B2(n_150),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_112),
.B(n_135),
.C(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_112),
.A2(n_113),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_112),
.A2(n_113),
.B1(n_169),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_113),
.B(n_161),
.C(n_169),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_113),
.B(n_141),
.C(n_145),
.Y(n_291)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_117),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_125),
.C(n_126),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_122),
.B(n_125),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_172),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_132),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_128),
.A2(n_132),
.B1(n_133),
.B2(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_128),
.Y(n_280)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_132),
.A2(n_133),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_132),
.A2(n_133),
.B1(n_220),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_133),
.B(n_214),
.C(n_220),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_133),
.B(n_192),
.C(n_251),
.Y(n_255)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_135),
.A2(n_136),
.B1(n_183),
.B2(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_135),
.A2(n_136),
.B1(n_167),
.B2(n_180),
.Y(n_257)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_136),
.B(n_167),
.C(n_258),
.Y(n_261)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND3xp33_ASAP7_75t_SL g151 ( 
.A(n_138),
.B(n_152),
.C(n_153),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_139),
.B(n_140),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_146),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_173),
.B(n_288),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_171),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_155),
.B(n_171),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_160),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_156),
.B(n_158),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_160),
.B(n_286),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_161),
.A2(n_162),
.B1(n_275),
.B2(n_276),
.Y(n_274)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_167),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_163),
.A2(n_167),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_163),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_165),
.A2(n_194),
.B(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_167),
.A2(n_180),
.B1(n_235),
.B2(n_237),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_167),
.B(n_237),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_169),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_283),
.B(n_287),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_210),
.B(n_269),
.C(n_282),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_199),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_176),
.B(n_199),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_186),
.B2(n_198),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_178)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_179),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_179),
.B(n_185),
.C(n_198),
.Y(n_270)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_182),
.Y(n_185)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_186),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_196),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_188),
.A2(n_189),
.B1(n_191),
.B2(n_192),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_191),
.A2(n_192),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_192),
.B(n_243),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_192),
.B(n_243),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_205),
.C(n_206),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_200),
.A2(n_201),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_206),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_207),
.A2(n_209),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_207),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_207),
.B(n_240),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_209),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_268),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_229),
.B(n_267),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_226),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_213),
.B(n_226),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_214),
.A2(n_215),
.B1(n_263),
.B2(n_265),
.Y(n_262)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_219),
.B(n_234),
.Y(n_245)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_220),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_224),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_221),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_260),
.B(n_266),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_254),
.B(n_259),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_246),
.B(n_253),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_238),
.B(n_245),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_235),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_242),
.B(n_244),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_247),
.B(n_248),
.Y(n_253)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_251),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_255),
.B(n_256),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_261),
.B(n_262),
.Y(n_266)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_263),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_271),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_281),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_278),
.B2(n_279),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_279),
.C(n_281),
.Y(n_284)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_285),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_296),
.B(n_300),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_299),
.Y(n_298)
);


endmodule