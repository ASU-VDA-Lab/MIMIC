module fake_jpeg_26261_n_300 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_300);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_11),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_28),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_23),
.B(n_11),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_29),
.B(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_33),
.Y(n_39)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_30),
.A2(n_23),
.B(n_25),
.C(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_40),
.B(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_30),
.B(n_12),
.Y(n_43)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_46),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_29),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_56),
.Y(n_67)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_55),
.Y(n_85)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_22),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_57),
.B(n_64),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_26),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_28),
.B(n_27),
.C(n_26),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_62),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_47),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_63),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_43),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_21),
.B1(n_15),
.B2(n_24),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_66),
.A2(n_13),
.B1(n_42),
.B2(n_34),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_69),
.A2(n_64),
.B(n_57),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_70),
.B(n_12),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_26),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_71),
.A2(n_13),
.B(n_50),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_65),
.A2(n_33),
.B1(n_45),
.B2(n_39),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_82),
.B1(n_61),
.B2(n_63),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_40),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_61),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_33),
.B1(n_45),
.B2(n_39),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_75),
.A2(n_18),
.B1(n_13),
.B2(n_15),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_45),
.B1(n_21),
.B2(n_39),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_80),
.B1(n_83),
.B2(n_86),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_48),
.A2(n_39),
.B1(n_21),
.B2(n_44),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_56),
.A2(n_21),
.B1(n_34),
.B2(n_15),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_21),
.B1(n_44),
.B2(n_41),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_76),
.Y(n_115)
);

INVx4_ASAP7_75t_SL g89 ( 
.A(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_100),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_53),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_91),
.B(n_93),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_81),
.Y(n_92)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_95),
.Y(n_132)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_71),
.A2(n_61),
.B1(n_48),
.B2(n_51),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_97),
.B1(n_105),
.B2(n_110),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_71),
.A2(n_52),
.B1(n_50),
.B2(n_63),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_98),
.B(n_104),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_103),
.B(n_106),
.Y(n_116)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_62),
.Y(n_101)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_62),
.Y(n_102)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_50),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_73),
.A2(n_63),
.B1(n_15),
.B2(n_16),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_25),
.B(n_22),
.C(n_17),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_108),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_58),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_35),
.Y(n_109)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_79),
.A2(n_15),
.B1(n_16),
.B2(n_25),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_111),
.A2(n_87),
.B1(n_16),
.B2(n_25),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_70),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_112),
.B(n_117),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_106),
.A2(n_73),
.B1(n_86),
.B2(n_82),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_114),
.A2(n_115),
.B1(n_119),
.B2(n_139),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_115),
.A2(n_119),
.B(n_137),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_69),
.C(n_83),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_69),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_79),
.C(n_78),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_125),
.C(n_126),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_108),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_121),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_78),
.C(n_84),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_84),
.C(n_87),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_13),
.B1(n_18),
.B2(n_81),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_104),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_130),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_72),
.C(n_47),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_26),
.C(n_31),
.Y(n_146)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_20),
.Y(n_173)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_31),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_95),
.A2(n_107),
.B1(n_88),
.B2(n_90),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_136),
.A2(n_138),
.B1(n_129),
.B2(n_140),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_88),
.A2(n_72),
.B(n_77),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_90),
.A2(n_80),
.B1(n_16),
.B2(n_18),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_93),
.A2(n_105),
.B1(n_110),
.B2(n_96),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_140),
.A2(n_49),
.B(n_35),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_134),
.A2(n_106),
.B(n_91),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_142),
.A2(n_145),
.B(n_169),
.Y(n_178)
);

NAND3xp33_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_98),
.C(n_13),
.Y(n_144)
);

AOI21xp33_ASAP7_75t_L g183 ( 
.A1(n_144),
.A2(n_163),
.B(n_127),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_111),
.B(n_89),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_149),
.C(n_113),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_150),
.B1(n_152),
.B2(n_155),
.Y(n_179)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_157),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_26),
.C(n_31),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_136),
.A2(n_89),
.B1(n_92),
.B2(n_100),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_156),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_129),
.A2(n_123),
.B1(n_118),
.B2(n_132),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_135),
.A2(n_89),
.B1(n_92),
.B2(n_12),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_153),
.A2(n_154),
.B1(n_165),
.B2(n_113),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_123),
.A2(n_92),
.B1(n_18),
.B2(n_81),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_60),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_160),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_27),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

AOI32xp33_ASAP7_75t_L g163 ( 
.A1(n_117),
.A2(n_28),
.A3(n_35),
.B1(n_81),
.B2(n_24),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_164),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_115),
.A2(n_58),
.B1(n_49),
.B2(n_19),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_22),
.Y(n_166)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_112),
.B(n_31),
.Y(n_167)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_31),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_124),
.Y(n_177)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_175),
.B(n_177),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_158),
.C(n_171),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_187),
.C(n_188),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_199),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_161),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_184),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_141),
.B(n_119),
.C(n_124),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_138),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_189),
.A2(n_147),
.B1(n_142),
.B2(n_173),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_170),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_190),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_32),
.C(n_20),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_193),
.C(n_194),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_14),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_143),
.B(n_14),
.Y(n_194)
);

XOR2x2_ASAP7_75t_L g195 ( 
.A(n_143),
.B(n_14),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_195),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_154),
.A2(n_11),
.B(n_10),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_165),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_162),
.Y(n_202)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_209),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_151),
.C(n_167),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_208),
.C(n_211),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_146),
.C(n_169),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_152),
.C(n_145),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_166),
.Y(n_212)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_212),
.Y(n_225)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_213),
.A2(n_217),
.B1(n_186),
.B2(n_180),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_150),
.Y(n_215)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_215),
.Y(n_230)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_185),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_219),
.A2(n_221),
.B1(n_222),
.B2(n_199),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_176),
.B(n_149),
.C(n_14),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_175),
.C(n_193),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_196),
.B(n_11),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_186),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_236),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_229),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_213),
.A2(n_189),
.B1(n_179),
.B2(n_198),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_228),
.A2(n_233),
.B1(n_234),
.B2(n_237),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_188),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_177),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_238),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_218),
.C(n_208),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_240),
.C(n_205),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_201),
.A2(n_179),
.B1(n_198),
.B2(n_197),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_207),
.A2(n_219),
.B1(n_201),
.B2(n_222),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_215),
.A2(n_180),
.B1(n_178),
.B2(n_194),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_211),
.B(n_178),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_192),
.C(n_19),
.Y(n_240)
);

AO21x1_ASAP7_75t_L g241 ( 
.A1(n_230),
.A2(n_202),
.B(n_212),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_241),
.A2(n_0),
.B(n_2),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_10),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_235),
.B(n_210),
.Y(n_245)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

OAI221xp5_ASAP7_75t_L g248 ( 
.A1(n_239),
.A2(n_214),
.B1(n_237),
.B2(n_225),
.C(n_224),
.Y(n_248)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_248),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_205),
.C(n_220),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_251),
.C(n_10),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_234),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_250),
.A2(n_253),
.B(n_9),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_19),
.C(n_17),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_228),
.A2(n_238),
.B1(n_240),
.B2(n_223),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_252),
.A2(n_254),
.B1(n_8),
.B2(n_1),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_223),
.A2(n_229),
.B(n_231),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_236),
.A2(n_19),
.B1(n_17),
.B2(n_2),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_255),
.B(n_251),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_247),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_254),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_10),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_259),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_243),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_241),
.A2(n_8),
.B(n_1),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_261),
.A2(n_4),
.B(n_5),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_262),
.A2(n_263),
.B1(n_4),
.B2(n_5),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_246),
.A2(n_8),
.B1(n_2),
.B2(n_3),
.Y(n_263)
);

O2A1O1Ixp33_ASAP7_75t_L g269 ( 
.A1(n_265),
.A2(n_247),
.B(n_5),
.C(n_6),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_0),
.C(n_3),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_4),
.C(n_5),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_267),
.Y(n_278)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_268),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_271),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_277),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_276),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_264),
.A2(n_244),
.B1(n_242),
.B2(n_6),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_275),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_257),
.A2(n_244),
.B1(n_242),
.B2(n_6),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_4),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_270),
.A2(n_265),
.B(n_259),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_280),
.Y(n_288)
);

OAI31xp67_ASAP7_75t_L g280 ( 
.A1(n_269),
.A2(n_256),
.A3(n_258),
.B(n_266),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_273),
.A2(n_255),
.B(n_5),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_271),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_285),
.B(n_273),
.Y(n_287)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_287),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_277),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_289),
.A2(n_291),
.B(n_283),
.Y(n_293)
);

AO21x1_ASAP7_75t_L g292 ( 
.A1(n_290),
.A2(n_281),
.B(n_283),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_4),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_293),
.Y(n_296)
);

AO21x1_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_288),
.B(n_278),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_295),
.A2(n_296),
.B1(n_6),
.B2(n_7),
.Y(n_297)
);

NAND2xp33_ASAP7_75t_SL g298 ( 
.A(n_297),
.B(n_7),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_7),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_7),
.Y(n_300)
);


endmodule