module fake_jpeg_4839_n_68 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_68);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_68;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_66;

BUFx3_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx13_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx2_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_18),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_12),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_19),
.B(n_20),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

OA22x2_ASAP7_75t_L g23 ( 
.A1(n_16),
.A2(n_18),
.B1(n_20),
.B2(n_19),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_15),
.C(n_10),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_19),
.B(n_15),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_13),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_23),
.B1(n_14),
.B2(n_10),
.Y(n_36)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_28),
.Y(n_32)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_14),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_21),
.Y(n_35)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_24),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_34),
.A2(n_31),
.B1(n_24),
.B2(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_37),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_27),
.B1(n_9),
.B2(n_13),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_34),
.A2(n_32),
.B(n_35),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_42),
.A2(n_26),
.B(n_22),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_33),
.C(n_29),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_42),
.C(n_41),
.Y(n_50)
);

NAND3xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_23),
.C(n_26),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_46),
.B(n_9),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_27),
.B1(n_28),
.B2(n_22),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_49),
.B1(n_40),
.B2(n_28),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_54),
.C(n_12),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_51),
.A2(n_45),
.B1(n_11),
.B2(n_8),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_8),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_53),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_8),
.Y(n_53)
);

INVxp33_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_58),
.C(n_0),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_12),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_61),
.B1(n_56),
.B2(n_5),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_63),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_6),
.B1(n_7),
.B2(n_4),
.Y(n_63)
);

AOI322xp5_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_6),
.C1(n_7),
.C2(n_60),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_65),
.C(n_2),
.Y(n_67)
);

BUFx24_ASAP7_75t_SL g68 ( 
.A(n_67),
.Y(n_68)
);


endmodule