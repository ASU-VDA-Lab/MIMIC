module real_jpeg_25508_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_1),
.A2(n_42),
.B1(n_43),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_1),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_1),
.A2(n_58),
.B1(n_161),
.B2(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_1),
.A2(n_64),
.B1(n_65),
.B2(n_161),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_161),
.Y(n_251)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_4),
.A2(n_10),
.B1(n_51),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_4),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_4),
.A2(n_42),
.B1(n_43),
.B2(n_171),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_4),
.A2(n_64),
.B1(n_65),
.B2(n_171),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_171),
.Y(n_260)
);

INVx8_ASAP7_75t_SL g47 ( 
.A(n_5),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_6),
.A2(n_114),
.B(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_6),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_6),
.B(n_41),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_L g235 ( 
.A1(n_6),
.A2(n_64),
.B1(n_65),
.B2(n_168),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_6),
.B(n_30),
.C(n_67),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_6),
.B(n_89),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_6),
.A2(n_27),
.B1(n_254),
.B2(n_260),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_7),
.A2(n_51),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_7),
.A2(n_57),
.B1(n_64),
.B2(n_65),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_57),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_7),
.A2(n_42),
.B1(n_43),
.B2(n_57),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_8),
.A2(n_37),
.B1(n_51),
.B2(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_8),
.A2(n_37),
.B1(n_64),
.B2(n_65),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_8),
.A2(n_37),
.B1(n_42),
.B2(n_43),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_9),
.A2(n_64),
.B1(n_65),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_9),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_9),
.A2(n_42),
.B1(n_43),
.B2(n_72),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_72),
.Y(n_152)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_11),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_12),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_12),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_12),
.A2(n_42),
.B1(n_43),
.B2(n_112),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_12),
.A2(n_64),
.B1(n_65),
.B2(n_112),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_112),
.Y(n_246)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_14),
.A2(n_42),
.B1(n_43),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_14),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_14),
.A2(n_64),
.B1(n_65),
.B2(n_91),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_14),
.A2(n_50),
.B1(n_91),
.B2(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_91),
.Y(n_190)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_15),
.Y(n_102)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_15),
.Y(n_155)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_15),
.Y(n_261)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_141),
.B1(n_142),
.B2(n_317),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_18),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_140),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_121),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_21),
.B(n_121),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_75),
.C(n_95),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_22),
.A2(n_23),
.B1(n_75),
.B2(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_60),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_38),
.B2(n_59),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_25),
.B(n_61),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_25),
.A2(n_59),
.B(n_60),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_25),
.A2(n_26),
.B1(n_61),
.B2(n_302),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_33),
.B(n_35),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_27),
.A2(n_151),
.B(n_153),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_27),
.A2(n_35),
.B(n_153),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_27),
.A2(n_100),
.B(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_27),
.A2(n_251),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_28),
.B(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_28),
.A2(n_31),
.B1(n_152),
.B2(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_28),
.A2(n_250),
.B1(n_252),
.B2(n_253),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_29),
.A2(n_30),
.B1(n_67),
.B2(n_69),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_29),
.B(n_265),
.Y(n_264)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_36),
.B(n_101),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_38),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_52),
.B(n_55),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_39),
.A2(n_111),
.B(n_116),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_39),
.B(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_39),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_39),
.A2(n_41),
.B1(n_170),
.B2(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_39),
.A2(n_41),
.B1(n_111),
.B2(n_178),
.Y(n_289)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_48),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_40),
.B(n_53),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_40),
.A2(n_125),
.B(n_127),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_40),
.A2(n_164),
.B1(n_165),
.B2(n_169),
.Y(n_163)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_42),
.A2(n_43),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_42),
.A2(n_46),
.B(n_167),
.C(n_186),
.Y(n_185)
);

HAxp5_ASAP7_75t_SL g212 ( 
.A(n_42),
.B(n_168),
.CON(n_212),
.SN(n_212)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

NAND3xp33_ASAP7_75t_L g186 ( 
.A(n_43),
.B(n_45),
.C(n_54),
.Y(n_186)
);

OAI32xp33_ASAP7_75t_L g211 ( 
.A1(n_43),
.A2(n_65),
.A3(n_88),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_46),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_51),
.Y(n_115)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_54),
.B(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_54),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_61),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_71),
.B(n_73),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_62),
.A2(n_71),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_62),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_62),
.A2(n_73),
.B(n_80),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_62),
.A2(n_109),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_62),
.A2(n_78),
.B(n_218),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_62),
.A2(n_109),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_62),
.A2(n_109),
.B1(n_217),
.B2(n_236),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_70),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_67),
.B2(n_69),
.Y(n_63)
);

AO22x1_ASAP7_75t_L g89 ( 
.A1(n_64),
.A2(n_65),
.B1(n_87),
.B2(n_88),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_64),
.B(n_87),
.Y(n_213)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_65),
.B(n_238),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_70),
.A2(n_79),
.B(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_70),
.A2(n_81),
.B(n_108),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_70),
.B(n_168),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_75),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_83),
.B(n_94),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_83),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_81),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_90),
.B1(n_92),
.B2(n_93),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_84),
.A2(n_93),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_L g181 ( 
.A1(n_84),
.A2(n_162),
.B(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_84),
.A2(n_93),
.B1(n_160),
.B2(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_84),
.A2(n_135),
.B(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_85),
.B(n_120),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_85),
.A2(n_133),
.B(n_134),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_85),
.A2(n_89),
.B1(n_203),
.B2(n_212),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_89),
.Y(n_85)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_89),
.B(n_120),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_89),
.B(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_93),
.B(n_119),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

FAx1_ASAP7_75t_SL g121 ( 
.A(n_94),
.B(n_122),
.CI(n_139),
.CON(n_121),
.SN(n_121)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_95),
.A2(n_96),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_110),
.C(n_117),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_97),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_105),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_98),
.A2(n_99),
.B1(n_105),
.B2(n_106),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_102),
.A2(n_103),
.B(n_190),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_102),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_102),
.B(n_168),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_104),
.B(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_110),
.A2(n_117),
.B1(n_118),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_110),
.Y(n_305)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx24_ASAP7_75t_SL g318 ( 
.A(n_121),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_129),
.B2(n_130),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_136),
.B2(n_137),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_310),
.B(n_316),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_297),
.B(n_309),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_204),
.B(n_280),
.C(n_296),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_191),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_146),
.B(n_191),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_174),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_156),
.B1(n_172),
.B2(n_173),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_148),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_148),
.B(n_173),
.C(n_174),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_149),
.B(n_150),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.C(n_163),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_157),
.A2(n_158),
.B1(n_159),
.B2(n_194),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_163),
.B(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_184),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_180),
.B2(n_181),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_177),
.B(n_180),
.C(n_184),
.Y(n_294)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_183),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_185),
.A2(n_187),
.B1(n_188),
.B2(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.C(n_197),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_192),
.B(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_195),
.B(n_197),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.C(n_201),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_223),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_198),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_275),
.B(n_279),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_230),
.B(n_274),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_219),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_209),
.B(n_219),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_215),
.C(n_216),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_210),
.B(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_214),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_215),
.B(n_216),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_224),
.B2(n_225),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_220),
.B(n_227),
.C(n_229),
.Y(n_276)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_226),
.Y(n_229)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_269),
.B(n_273),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_247),
.B(n_268),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_239),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_233),
.B(n_239),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_237),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_237),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_245),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_244),
.C(n_245),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_243),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_246),
.Y(n_252)
);

AOI21xp33_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_256),
.B(n_267),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_255),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_255),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_262),
.B(n_266),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_258),
.B(n_259),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_270),
.B(n_271),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_276),
.B(n_277),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_282),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_294),
.B2(n_295),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_286),
.C(n_295),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_293),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_290),
.C(n_293),
.Y(n_308)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_294),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_298),
.B(n_299),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_308),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_303),
.B1(n_306),
.B2(n_307),
.Y(n_300)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_301),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_307),
.C(n_308),
.Y(n_311)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_303),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_311),
.B(n_312),
.Y(n_316)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);


endmodule