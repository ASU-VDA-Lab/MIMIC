module fake_jpeg_2577_n_682 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_682);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_682;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_19),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_14),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_60),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_32),
.Y(n_61)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_61),
.Y(n_202)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_62),
.Y(n_174)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_63),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_41),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_64),
.B(n_80),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_66),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_67),
.Y(n_210)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_68),
.Y(n_148)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g169 ( 
.A(n_70),
.Y(n_169)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_71),
.Y(n_168)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_72),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_73),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_74),
.Y(n_175)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_75),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_76),
.Y(n_198)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_77),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_78),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_79),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_27),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_81),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_82),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_84),
.Y(n_192)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_23),
.B(n_16),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_86),
.B(n_95),
.Y(n_159)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_87),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_88),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_89),
.Y(n_201)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx8_ASAP7_75t_L g206 ( 
.A(n_90),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_91),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_92),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_23),
.B(n_16),
.Y(n_95)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx11_ASAP7_75t_L g173 ( 
.A(n_96),
.Y(n_173)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

INVx4_ASAP7_75t_SL g98 ( 
.A(n_54),
.Y(n_98)
);

INVx13_ASAP7_75t_L g209 ( 
.A(n_98),
.Y(n_209)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_99),
.Y(n_193)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_100),
.Y(n_221)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_101),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_102),
.Y(n_184)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_103),
.Y(n_204)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_104),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_105),
.Y(n_164)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_29),
.Y(n_106)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_106),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

BUFx8_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

BUFx16f_ASAP7_75t_L g109 ( 
.A(n_34),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_109),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_44),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g196 ( 
.A(n_110),
.Y(n_196)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_32),
.Y(n_111)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_38),
.Y(n_112)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_112),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g226 ( 
.A(n_113),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_37),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_118),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_29),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_116),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_22),
.B(n_16),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_117),
.B(n_123),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_37),
.Y(n_118)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_32),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_119),
.Y(n_190)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_43),
.Y(n_120)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_30),
.Y(n_121)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_38),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_130),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_22),
.B(n_40),
.Y(n_123)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_30),
.Y(n_124)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_124),
.Y(n_178)
);

BUFx24_ASAP7_75t_L g125 ( 
.A(n_30),
.Y(n_125)
);

CKINVDCx12_ASAP7_75t_R g134 ( 
.A(n_125),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_37),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_128),
.Y(n_162)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_43),
.Y(n_127)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_127),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_30),
.B(n_17),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_48),
.Y(n_129)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_129),
.Y(n_185)
);

INVxp67_ASAP7_75t_SL g130 ( 
.A(n_49),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_55),
.Y(n_131)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_131),
.Y(n_186)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_49),
.Y(n_132)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_132),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_57),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_136),
.B(n_170),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_116),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_137),
.B(n_138),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_95),
.B(n_57),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_74),
.A2(n_38),
.B1(n_42),
.B2(n_36),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_150),
.A2(n_163),
.B1(n_88),
.B2(n_113),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_123),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_152),
.B(n_155),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_62),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_60),
.A2(n_56),
.B1(n_55),
.B2(n_50),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_157),
.A2(n_165),
.B1(n_167),
.B2(n_172),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_85),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_160),
.B(n_228),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_78),
.A2(n_42),
.B1(n_36),
.B2(n_39),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_117),
.A2(n_50),
.B1(n_56),
.B2(n_55),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_87),
.A2(n_50),
.B1(n_56),
.B2(n_42),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_98),
.B(n_47),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_90),
.A2(n_39),
.B1(n_47),
.B2(n_46),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_130),
.B(n_128),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_177),
.B(n_181),
.Y(n_264)
);

HAxp5_ASAP7_75t_SL g180 ( 
.A(n_109),
.B(n_39),
.CON(n_180),
.SN(n_180)
);

AOI21xp33_ASAP7_75t_L g291 ( 
.A1(n_180),
.A2(n_227),
.B(n_6),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_61),
.B(n_53),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_102),
.B(n_46),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_183),
.B(n_187),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_102),
.B(n_40),
.Y(n_187)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_131),
.Y(n_197)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_197),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_89),
.B(n_53),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_199),
.B(n_217),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_106),
.A2(n_51),
.B(n_39),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_200),
.B(n_114),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_119),
.B(n_51),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_205),
.B(n_5),
.Y(n_285)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_129),
.Y(n_208)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_208),
.Y(n_261)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_67),
.Y(n_215)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_215),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_73),
.B(n_15),
.Y(n_217)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_79),
.Y(n_219)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_219),
.Y(n_283)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_81),
.Y(n_223)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_223),
.Y(n_308)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_83),
.Y(n_225)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

HAxp5_ASAP7_75t_SL g227 ( 
.A(n_125),
.B(n_15),
.CON(n_227),
.SN(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_91),
.Y(n_228)
);

BUFx4f_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_230),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_231),
.Y(n_329)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_184),
.Y(n_233)
);

INVx4_ASAP7_75t_SL g357 ( 
.A(n_233),
.Y(n_357)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_168),
.Y(n_236)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_236),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_15),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_237),
.B(n_255),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_201),
.Y(n_238)
);

INVx5_ASAP7_75t_L g339 ( 
.A(n_238),
.Y(n_339)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_156),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_239),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_205),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_240),
.B(n_244),
.Y(n_320)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_184),
.Y(n_241)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_241),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_242),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_133),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_209),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_245),
.B(n_272),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_246),
.A2(n_275),
.B1(n_279),
.B2(n_292),
.Y(n_317)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_207),
.Y(n_247)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_247),
.Y(n_346)
);

BUFx12f_ASAP7_75t_L g248 ( 
.A(n_209),
.Y(n_248)
);

INVx8_ASAP7_75t_L g368 ( 
.A(n_248),
.Y(n_368)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_192),
.Y(n_249)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_249),
.Y(n_327)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_194),
.Y(n_250)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_250),
.Y(n_335)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_194),
.Y(n_251)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_251),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_156),
.Y(n_253)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_253),
.Y(n_340)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_175),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_254),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_159),
.B(n_110),
.Y(n_255)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_210),
.Y(n_256)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_256),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_257),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_161),
.A2(n_0),
.B(n_1),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_258),
.A2(n_291),
.B(n_146),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_193),
.B(n_93),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_259),
.B(n_269),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_210),
.Y(n_260)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_260),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_157),
.A2(n_105),
.B1(n_92),
.B2(n_3),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_262),
.A2(n_218),
.B1(n_214),
.B2(n_206),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_188),
.Y(n_263)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_263),
.Y(n_350)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_194),
.Y(n_266)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_266),
.Y(n_351)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_204),
.Y(n_267)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_267),
.Y(n_353)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_216),
.Y(n_268)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_268),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_140),
.B(n_0),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_145),
.Y(n_270)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_270),
.Y(n_367)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_207),
.Y(n_271)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_271),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_189),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_158),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_273),
.A2(n_280),
.B1(n_141),
.B2(n_182),
.Y(n_313)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_224),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_274),
.B(n_284),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g275 ( 
.A(n_190),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_148),
.B(n_135),
.C(n_139),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_276),
.B(n_309),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_212),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_277),
.Y(n_337)
);

BUFx8_ASAP7_75t_L g279 ( 
.A(n_149),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_195),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_211),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_285),
.B(n_287),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_161),
.B(n_5),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_286),
.B(n_288),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_176),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_198),
.Y(n_288)
);

INVx6_ASAP7_75t_SL g289 ( 
.A(n_134),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_289),
.B(n_290),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_162),
.B(n_6),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_180),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_144),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_293),
.A2(n_297),
.B1(n_300),
.B2(n_306),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_142),
.B(n_7),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_294),
.B(n_295),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_213),
.B(n_8),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_143),
.B(n_222),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_296),
.B(n_298),
.Y(n_356)
);

AO22x2_ASAP7_75t_L g297 ( 
.A1(n_229),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_221),
.B(n_9),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_169),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_299),
.B(n_301),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_144),
.A2(n_13),
.B1(n_150),
.B2(n_176),
.Y(n_300)
);

NOR4xp25_ASAP7_75t_L g301 ( 
.A(n_166),
.B(n_13),
.C(n_178),
.D(n_149),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_169),
.B(n_154),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_302),
.B(n_303),
.Y(n_360)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_212),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_171),
.B(n_198),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_304),
.B(n_305),
.Y(n_365)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_147),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_171),
.A2(n_163),
.B1(n_220),
.B2(n_227),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_185),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_307),
.A2(n_310),
.B1(n_279),
.B2(n_248),
.Y(n_336)
);

AND2x2_ASAP7_75t_SL g309 ( 
.A(n_220),
.B(n_186),
.Y(n_309)
);

AND2x2_ASAP7_75t_SL g319 ( 
.A(n_309),
.B(n_226),
.Y(n_319)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_153),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_153),
.B(n_206),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_312),
.A2(n_214),
.B1(n_218),
.B2(n_174),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_313),
.B(n_324),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_315),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_264),
.B(n_282),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_316),
.B(n_322),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_319),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_276),
.B(n_174),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_323),
.A2(n_338),
.B1(n_343),
.B2(n_279),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_257),
.A2(n_191),
.B1(n_151),
.B2(n_164),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_232),
.B(n_141),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_328),
.B(n_330),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_278),
.B(n_286),
.Y(n_330)
);

AND2x2_ASAP7_75t_SL g332 ( 
.A(n_265),
.B(n_226),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g394 ( 
.A(n_332),
.Y(n_394)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_336),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_246),
.A2(n_179),
.B1(n_182),
.B2(n_191),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_306),
.A2(n_179),
.B1(n_151),
.B2(n_164),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_345),
.B(n_371),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_300),
.A2(n_146),
.B(n_173),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_354),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_L g358 ( 
.A1(n_311),
.A2(n_173),
.B1(n_164),
.B2(n_151),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_358),
.A2(n_361),
.B1(n_254),
.B2(n_263),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_262),
.A2(n_196),
.B1(n_226),
.B2(n_258),
.Y(n_361)
);

FAx1_ASAP7_75t_SL g362 ( 
.A(n_234),
.B(n_252),
.CI(n_309),
.CON(n_362),
.SN(n_362)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_362),
.B(n_230),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_230),
.A2(n_274),
.B1(n_288),
.B2(n_284),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_SL g396 ( 
.A1(n_366),
.A2(n_248),
.B1(n_266),
.B2(n_250),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_369),
.B(n_308),
.C(n_283),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_297),
.A2(n_196),
.B1(n_247),
.B2(n_271),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_297),
.B(n_196),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_374),
.B(n_293),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_331),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_375),
.B(n_407),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_376),
.A2(n_381),
.B1(n_400),
.B2(n_401),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_373),
.A2(n_235),
.B1(n_308),
.B2(n_283),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_377),
.A2(n_348),
.B1(n_340),
.B2(n_370),
.Y(n_456)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_314),
.Y(n_378)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_378),
.Y(n_431)
);

AND2x6_ASAP7_75t_L g380 ( 
.A(n_362),
.B(n_289),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_380),
.B(n_413),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_374),
.A2(n_292),
.B1(n_297),
.B2(n_303),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_382),
.B(n_404),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_383),
.B(n_384),
.C(n_332),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_369),
.B(n_307),
.C(n_231),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_368),
.Y(n_385)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_385),
.Y(n_438)
);

INVx13_ASAP7_75t_L g386 ( 
.A(n_368),
.Y(n_386)
);

CKINVDCx14_ASAP7_75t_R g454 ( 
.A(n_386),
.Y(n_454)
);

INVx8_ASAP7_75t_L g387 ( 
.A(n_363),
.Y(n_387)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_387),
.Y(n_442)
);

INVx8_ASAP7_75t_L g388 ( 
.A(n_363),
.Y(n_388)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_388),
.Y(n_464)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_314),
.Y(n_389)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_389),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_L g429 ( 
.A1(n_390),
.A2(n_337),
.B1(n_357),
.B2(n_315),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_372),
.B(n_233),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_391),
.Y(n_444)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_321),
.Y(n_395)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_395),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_SL g432 ( 
.A1(n_396),
.A2(n_406),
.B1(n_420),
.B2(n_357),
.Y(n_432)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_321),
.Y(n_399)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_399),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_318),
.A2(n_256),
.B1(n_239),
.B2(n_281),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_322),
.A2(n_253),
.B1(n_277),
.B2(n_260),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_372),
.B(n_241),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_402),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_316),
.B(n_243),
.Y(n_404)
);

INVx13_ASAP7_75t_L g406 ( 
.A(n_357),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_325),
.B(n_251),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_327),
.Y(n_408)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_408),
.Y(n_441)
);

CKINVDCx14_ASAP7_75t_R g409 ( 
.A(n_319),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_409),
.B(n_410),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_320),
.B(n_238),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_328),
.B(n_243),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_411),
.B(n_414),
.Y(n_448)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_342),
.Y(n_412)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_412),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_356),
.B(n_261),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_360),
.B(n_261),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_415),
.B(n_416),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_349),
.B(n_281),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_332),
.B(n_242),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_417),
.B(n_319),
.Y(n_426)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_327),
.Y(n_418)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_418),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_347),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_419),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_341),
.B(n_330),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_323),
.A2(n_371),
.B1(n_361),
.B2(n_324),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_421),
.A2(n_345),
.B1(n_313),
.B2(n_354),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_343),
.A2(n_338),
.B1(n_359),
.B2(n_334),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_423),
.A2(n_352),
.B(n_362),
.Y(n_437)
);

XNOR2x1_ASAP7_75t_SL g498 ( 
.A(n_426),
.B(n_434),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_427),
.A2(n_433),
.B1(n_439),
.B2(n_443),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_429),
.A2(n_457),
.B1(n_458),
.B2(n_376),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_432),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_393),
.A2(n_423),
.B1(n_413),
.B2(n_379),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_382),
.A2(n_317),
.B(n_365),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_436),
.B(n_384),
.C(n_383),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_437),
.B(n_445),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_393),
.A2(n_337),
.B1(n_367),
.B2(n_364),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_379),
.A2(n_353),
.B1(n_367),
.B2(n_364),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_392),
.A2(n_353),
.B(n_350),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_392),
.A2(n_394),
.B(n_422),
.Y(n_447)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_447),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_379),
.A2(n_342),
.B1(n_348),
.B2(n_340),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_452),
.B(n_455),
.Y(n_472)
);

OA21x2_ASAP7_75t_L g455 ( 
.A1(n_421),
.A2(n_370),
.B(n_350),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_SL g470 ( 
.A1(n_456),
.A2(n_390),
.B1(n_418),
.B2(n_395),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_381),
.A2(n_363),
.B1(n_333),
.B2(n_326),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_405),
.A2(n_333),
.B1(n_326),
.B2(n_346),
.Y(n_458)
);

AO22x1_ASAP7_75t_L g460 ( 
.A1(n_392),
.A2(n_346),
.B1(n_339),
.B2(n_329),
.Y(n_460)
);

OA21x2_ASAP7_75t_L g469 ( 
.A1(n_460),
.A2(n_462),
.B(n_447),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_405),
.A2(n_339),
.B1(n_351),
.B2(n_355),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_461),
.B(n_377),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_422),
.A2(n_398),
.B(n_417),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_440),
.B(n_419),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_466),
.B(n_490),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_433),
.A2(n_400),
.B1(n_403),
.B2(n_375),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_467),
.B(n_469),
.Y(n_523)
);

CKINVDCx12_ASAP7_75t_R g468 ( 
.A(n_454),
.Y(n_468)
);

CKINVDCx14_ASAP7_75t_R g517 ( 
.A(n_468),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_470),
.A2(n_473),
.B1(n_429),
.B2(n_425),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_SL g473 ( 
.A1(n_461),
.A2(n_403),
.B1(n_385),
.B2(n_401),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_439),
.Y(n_474)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_474),
.Y(n_507)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_428),
.Y(n_476)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_476),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_SL g525 ( 
.A1(n_478),
.A2(n_500),
.B1(n_455),
.B2(n_460),
.Y(n_525)
);

INVx5_ASAP7_75t_L g479 ( 
.A(n_442),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_479),
.B(n_501),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_440),
.B(n_397),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_480),
.B(n_485),
.Y(n_516)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_481),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_482),
.B(n_487),
.C(n_489),
.Y(n_529)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_431),
.Y(n_483)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_483),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_448),
.B(n_404),
.Y(n_484)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_484),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_444),
.B(n_463),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_448),
.B(n_411),
.Y(n_486)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_486),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_436),
.B(n_397),
.C(n_414),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_446),
.B(n_415),
.Y(n_488)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_488),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_426),
.B(n_416),
.C(n_380),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_446),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_453),
.B(n_399),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_491),
.B(n_492),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_453),
.B(n_408),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_430),
.B(n_351),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_493),
.B(n_424),
.Y(n_533)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_428),
.Y(n_494)
);

NAND2xp33_ASAP7_75t_SL g512 ( 
.A(n_494),
.B(n_497),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_437),
.B(n_412),
.C(n_344),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_495),
.B(n_445),
.Y(n_506)
);

INVx13_ASAP7_75t_L g496 ( 
.A(n_454),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_496),
.Y(n_526)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_435),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_443),
.B(n_378),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_499),
.B(n_502),
.Y(n_511)
);

INVx13_ASAP7_75t_L g500 ( 
.A(n_462),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_442),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_450),
.B(n_389),
.Y(n_502)
);

XNOR2x1_ASAP7_75t_L g503 ( 
.A(n_498),
.B(n_434),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_SL g548 ( 
.A(n_503),
.B(n_538),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_477),
.A2(n_425),
.B1(n_451),
.B2(n_427),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_504),
.A2(n_518),
.B1(n_515),
.B2(n_507),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_506),
.B(n_532),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_508),
.A2(n_522),
.B1(n_525),
.B2(n_469),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_500),
.A2(n_451),
.B(n_449),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_509),
.A2(n_471),
.B(n_472),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_466),
.B(n_430),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g560 ( 
.A(n_514),
.B(n_519),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_490),
.B(n_452),
.Y(n_515)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_515),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_487),
.B(n_449),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_491),
.B(n_450),
.Y(n_520)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_520),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_479),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_521),
.B(n_534),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_475),
.A2(n_460),
.B1(n_455),
.B2(n_457),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_492),
.B(n_486),
.Y(n_528)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_528),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_482),
.B(n_455),
.Y(n_532)
);

CKINVDCx14_ASAP7_75t_R g540 ( 
.A(n_533),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_488),
.B(n_495),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_489),
.B(n_435),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_535),
.B(n_538),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_501),
.B(n_438),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_536),
.B(n_464),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_498),
.B(n_441),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_465),
.B(n_441),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_539),
.B(n_477),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_516),
.B(n_484),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_SL g587 ( 
.A(n_543),
.B(n_550),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_527),
.B(n_474),
.Y(n_545)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_545),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_532),
.B(n_467),
.Y(n_546)
);

MAJx2_ASAP7_75t_L g590 ( 
.A(n_546),
.B(n_548),
.C(n_553),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_549),
.A2(n_558),
.B1(n_563),
.B2(n_523),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_517),
.B(n_438),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_SL g593 ( 
.A(n_551),
.B(n_510),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_529),
.B(n_535),
.C(n_506),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_552),
.B(n_541),
.C(n_553),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_529),
.B(n_469),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_520),
.B(n_512),
.Y(n_554)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_554),
.Y(n_591)
);

INVx1_ASAP7_75t_SL g555 ( 
.A(n_513),
.Y(n_555)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_555),
.Y(n_572)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_513),
.Y(n_557)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_557),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_518),
.A2(n_472),
.B1(n_475),
.B2(n_500),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_L g597 ( 
.A1(n_559),
.A2(n_522),
.B(n_478),
.Y(n_597)
);

NOR3xp33_ASAP7_75t_SL g562 ( 
.A(n_530),
.B(n_471),
.C(n_497),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_SL g595 ( 
.A(n_562),
.B(n_564),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_530),
.B(n_464),
.Y(n_564)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_539),
.B(n_469),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g592 ( 
.A(n_565),
.B(n_569),
.Y(n_592)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_511),
.Y(n_566)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_566),
.Y(n_580)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_567),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_537),
.B(n_494),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_568),
.B(n_540),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_537),
.B(n_499),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_511),
.Y(n_570)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_570),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_509),
.B(n_481),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g594 ( 
.A(n_571),
.B(n_551),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_560),
.B(n_505),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_573),
.B(n_575),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_SL g599 ( 
.A1(n_574),
.A2(n_597),
.B1(n_563),
.B2(n_542),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_554),
.Y(n_575)
);

BUFx5_ASAP7_75t_L g577 ( 
.A(n_562),
.Y(n_577)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_577),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_579),
.B(n_581),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_552),
.B(n_523),
.C(n_507),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_541),
.B(n_523),
.C(n_503),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_582),
.B(n_583),
.C(n_588),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_546),
.B(n_504),
.C(n_526),
.Y(n_583)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_585),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_547),
.B(n_526),
.C(n_531),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_569),
.B(n_528),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_589),
.B(n_597),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_SL g618 ( 
.A(n_593),
.B(n_594),
.Y(n_618)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_555),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_596),
.B(n_572),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_SL g598 ( 
.A1(n_574),
.A2(n_559),
.B(n_545),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_598),
.B(n_608),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_599),
.A2(n_577),
.B1(n_578),
.B2(n_458),
.Y(n_633)
);

XNOR2xp5_ASAP7_75t_L g600 ( 
.A(n_594),
.B(n_547),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g635 ( 
.A(n_600),
.B(n_611),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_591),
.A2(n_544),
.B1(n_556),
.B2(n_531),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_603),
.A2(n_596),
.B1(n_599),
.B2(n_601),
.Y(n_625)
);

CKINVDCx16_ASAP7_75t_R g605 ( 
.A(n_589),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_605),
.B(n_606),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_587),
.B(n_561),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_595),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_SL g609 ( 
.A1(n_576),
.A2(n_584),
.B1(n_580),
.B2(n_586),
.Y(n_609)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_609),
.Y(n_622)
);

XOR2xp5_ASAP7_75t_L g611 ( 
.A(n_581),
.B(n_571),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_SL g612 ( 
.A1(n_580),
.A2(n_558),
.B1(n_548),
.B2(n_565),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_612),
.B(n_578),
.Y(n_636)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_588),
.B(n_592),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_613),
.B(n_614),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g614 ( 
.A(n_592),
.B(n_510),
.Y(n_614)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_616),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_584),
.B(n_387),
.Y(n_617)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_617),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_572),
.B(n_524),
.Y(n_619)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_619),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_607),
.B(n_586),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_SL g641 ( 
.A(n_623),
.B(n_626),
.Y(n_641)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_625),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_615),
.B(n_583),
.Y(n_626)
);

AOI21x1_ASAP7_75t_L g629 ( 
.A1(n_604),
.A2(n_582),
.B(n_590),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_629),
.A2(n_600),
.B(n_618),
.Y(n_649)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_611),
.B(n_579),
.C(n_593),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_631),
.B(n_632),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_602),
.B(n_590),
.C(n_524),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_633),
.A2(n_603),
.B1(n_619),
.B2(n_614),
.Y(n_644)
);

BUFx24_ASAP7_75t_SL g634 ( 
.A(n_601),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_SL g650 ( 
.A(n_634),
.B(n_636),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_613),
.B(n_502),
.C(n_483),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_637),
.B(n_476),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_627),
.B(n_598),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_638),
.B(n_642),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_630),
.B(n_616),
.Y(n_640)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_640),
.B(n_644),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_621),
.Y(n_642)
);

CKINVDCx16_ASAP7_75t_R g645 ( 
.A(n_620),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_645),
.B(n_647),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_624),
.B(n_610),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_646),
.Y(n_660)
);

CKINVDCx16_ASAP7_75t_R g647 ( 
.A(n_637),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_622),
.B(n_610),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_648),
.B(n_652),
.Y(n_657)
);

OAI21xp5_ASAP7_75t_L g654 ( 
.A1(n_649),
.A2(n_636),
.B(n_612),
.Y(n_654)
);

XOR2xp5_ASAP7_75t_L g663 ( 
.A(n_651),
.B(n_459),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_632),
.B(n_635),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_654),
.B(n_659),
.Y(n_666)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_646),
.B(n_635),
.C(n_631),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_655),
.B(n_658),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_641),
.B(n_628),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_643),
.B(n_618),
.C(n_633),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_650),
.B(n_459),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_SL g668 ( 
.A(n_661),
.B(n_663),
.Y(n_668)
);

AOI221xp5_ASAP7_75t_L g664 ( 
.A1(n_660),
.A2(n_639),
.B1(n_644),
.B2(n_640),
.C(n_649),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_SL g672 ( 
.A1(n_664),
.A2(n_662),
.B(n_653),
.Y(n_672)
);

MAJIxp5_ASAP7_75t_L g665 ( 
.A(n_655),
.B(n_642),
.C(n_639),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_665),
.B(n_667),
.Y(n_671)
);

OAI22xp5_ASAP7_75t_SL g667 ( 
.A1(n_662),
.A2(n_424),
.B1(n_496),
.B2(n_468),
.Y(n_667)
);

MAJIxp5_ASAP7_75t_L g669 ( 
.A(n_657),
.B(n_431),
.C(n_456),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_669),
.B(n_659),
.Y(n_673)
);

XNOR2xp5_ASAP7_75t_L g675 ( 
.A(n_672),
.B(n_673),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_668),
.B(n_656),
.Y(n_674)
);

AOI322xp5_ASAP7_75t_L g676 ( 
.A1(n_674),
.A2(n_666),
.A3(n_670),
.B1(n_664),
.B2(n_496),
.C1(n_663),
.C2(n_386),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_676),
.B(n_335),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_SL g677 ( 
.A1(n_675),
.A2(n_671),
.B(n_344),
.Y(n_677)
);

OAI21xp33_ASAP7_75t_L g679 ( 
.A1(n_677),
.A2(n_678),
.B(n_406),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_679),
.B(n_335),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_680),
.B(n_388),
.Y(n_681)
);

MAJIxp5_ASAP7_75t_L g682 ( 
.A(n_681),
.B(n_329),
.C(n_406),
.Y(n_682)
);


endmodule