module fake_jpeg_16555_n_43 (n_3, n_2, n_1, n_0, n_4, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

INVx4_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx11_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

NAND3xp33_ASAP7_75t_L g14 ( 
.A(n_7),
.B(n_0),
.C(n_1),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_15),
.Y(n_22)
);

BUFx2_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_8),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_11),
.C(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_5),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_20),
.Y(n_24)
);

CKINVDCx12_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_7),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_28),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_17),
.C(n_13),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_6),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_30),
.B(n_31),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_24),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_27),
.C(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_13),
.Y(n_34)
);

NOR2xp67_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_35),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_9),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_33),
.C(n_34),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_39),
.A2(n_40),
.B1(n_38),
.B2(n_28),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_38),
.B(n_21),
.Y(n_43)
);


endmodule