module fake_jpeg_3314_n_204 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_204);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_23),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_9),
.Y(n_54)
);

BUFx4f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_4),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_28),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_17),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_39),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_12),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_20),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_80),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NOR2xp67_ASAP7_75t_SL g81 ( 
.A(n_76),
.B(n_58),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_73),
.A2(n_51),
.B1(n_62),
.B2(n_60),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_88),
.B1(n_55),
.B2(n_68),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_70),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_94),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_73),
.A2(n_51),
.B1(n_58),
.B2(n_63),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_64),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_55),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_74),
.B(n_54),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_93),
.B(n_68),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_65),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_95),
.A2(n_111),
.B1(n_57),
.B2(n_87),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_100),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_79),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_97),
.Y(n_126)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_72),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_102),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_50),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_106),
.Y(n_117)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_90),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_90),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_109),
.Y(n_127)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_110),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_81),
.A2(n_72),
.B1(n_57),
.B2(n_80),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_87),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_46),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

MAJx2_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_66),
.C(n_52),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_0),
.C(n_1),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_101),
.A2(n_80),
.B1(n_78),
.B2(n_56),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_115),
.A2(n_120),
.B1(n_131),
.B2(n_32),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_101),
.A2(n_86),
.B1(n_91),
.B2(n_66),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_119),
.A2(n_43),
.B(n_41),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_111),
.A2(n_56),
.B1(n_57),
.B2(n_69),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_91),
.B1(n_71),
.B2(n_67),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_122),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_49),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_132),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_37),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_102),
.A2(n_108),
.B1(n_110),
.B2(n_103),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_45),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_116),
.B(n_44),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_138),
.Y(n_164)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_126),
.A2(n_119),
.B1(n_123),
.B2(n_132),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_140),
.B1(n_22),
.B2(n_8),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_136),
.A2(n_149),
.B1(n_151),
.B2(n_10),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_139),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_117),
.B(n_2),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_114),
.A2(n_128),
.B1(n_122),
.B2(n_131),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_122),
.B(n_3),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_122),
.A2(n_36),
.B(n_35),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_147),
.A2(n_153),
.B(n_155),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_3),
.Y(n_148)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_5),
.Y(n_150)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_5),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_152),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_6),
.B(n_7),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_154),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_6),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_137),
.A2(n_30),
.B1(n_27),
.B2(n_24),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_157),
.A2(n_158),
.B1(n_163),
.B2(n_167),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_169),
.C(n_153),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_140),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_167)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_168),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_11),
.Y(n_169)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_176),
.Y(n_189)
);

AOI321xp33_ASAP7_75t_L g177 ( 
.A1(n_173),
.A2(n_133),
.A3(n_137),
.B1(n_142),
.B2(n_147),
.C(n_136),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_170),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_179),
.Y(n_190)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_181),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_149),
.C(n_14),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_182),
.Y(n_186)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_183),
.A2(n_165),
.B1(n_162),
.B2(n_156),
.Y(n_187)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_187),
.Y(n_193)
);

AO21x1_ASAP7_75t_L g188 ( 
.A1(n_177),
.A2(n_166),
.B(n_157),
.Y(n_188)
);

AOI31xp67_ASAP7_75t_L g194 ( 
.A1(n_188),
.A2(n_185),
.A3(n_184),
.B(n_189),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_185),
.A2(n_174),
.B1(n_166),
.B2(n_181),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_191),
.A2(n_194),
.B1(n_190),
.B2(n_15),
.Y(n_196)
);

NAND3xp33_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_180),
.C(n_159),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_195),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_169),
.C(n_175),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_196),
.A2(n_197),
.B1(n_13),
.B2(n_16),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_193),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_199),
.B(n_200),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_17),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_201),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_202),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_198),
.Y(n_204)
);


endmodule