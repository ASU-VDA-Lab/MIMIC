module fake_jpeg_17728_n_122 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_122);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_122;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx4_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_3),
.B(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_5),
.B(n_13),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_14),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_29),
.A2(n_26),
.B1(n_20),
.B2(n_4),
.Y(n_57)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_21),
.B(n_0),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_34),
.Y(n_56)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_21),
.B(n_2),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVxp33_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_16),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_26),
.B1(n_15),
.B2(n_22),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_18),
.Y(n_53)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_25),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_25),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_42),
.B(n_48),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_SL g43 ( 
.A1(n_37),
.A2(n_19),
.B(n_17),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_44),
.B1(n_58),
.B2(n_60),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_SL g44 ( 
.A1(n_32),
.A2(n_19),
.B(n_17),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_14),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_18),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_22),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_14),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_50),
.Y(n_75)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_53),
.B(n_59),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_57),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_36),
.A2(n_15),
.B1(n_26),
.B2(n_22),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_28),
.B(n_15),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_62),
.B(n_23),
.Y(n_74)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_31),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_74),
.Y(n_89)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_23),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_76),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_56),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_48),
.A2(n_23),
.B1(n_6),
.B2(n_8),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_77),
.B1(n_6),
.B2(n_12),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_23),
.Y(n_76)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_7),
.B(n_12),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_78),
.A2(n_13),
.B(n_55),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_55),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_79),
.A2(n_50),
.B1(n_49),
.B2(n_40),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_83),
.C(n_92),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_65),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_56),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_85),
.B(n_67),
.Y(n_101)
);

AOI322xp5_ASAP7_75t_SL g100 ( 
.A1(n_86),
.A2(n_63),
.A3(n_64),
.B1(n_67),
.B2(n_83),
.C1(n_81),
.C2(n_89),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_40),
.B1(n_54),
.B2(n_58),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_90),
.B1(n_93),
.B2(n_92),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_66),
.A2(n_58),
.B1(n_52),
.B2(n_62),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_58),
.C(n_47),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_70),
.A2(n_47),
.B1(n_76),
.B2(n_73),
.Y(n_93)
);

FAx1_ASAP7_75t_SL g94 ( 
.A(n_80),
.B(n_65),
.CI(n_67),
.CON(n_94),
.SN(n_94)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_94),
.B(n_96),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_95),
.A2(n_101),
.B1(n_103),
.B2(n_102),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_79),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_68),
.B1(n_77),
.B2(n_87),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_97),
.A2(n_82),
.B(n_84),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_75),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_99),
.Y(n_106)
);

NOR3xp33_ASAP7_75t_SL g99 ( 
.A(n_85),
.B(n_71),
.C(n_70),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_104),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_84),
.B(n_86),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_108),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_94),
.C(n_104),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_111),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_95),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_107),
.Y(n_114)
);

AOI322xp5_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_94),
.A3(n_99),
.B1(n_101),
.B2(n_103),
.C1(n_110),
.C2(n_106),
.Y(n_113)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

NOR2xp67_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_100),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_114),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_120),
.B(n_121),
.C(n_115),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_119),
.A2(n_116),
.B(n_113),
.Y(n_121)
);


endmodule