module fake_jpeg_13528_n_160 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_160);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_13),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_16),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVxp33_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_15),
.Y(n_64)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_29),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_45),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_2),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_19),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

BUFx24_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_74),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_54),
.Y(n_100)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_61),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_69),
.B1(n_77),
.B2(n_62),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_88),
.A2(n_66),
.B1(n_52),
.B2(n_4),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_77),
.B1(n_75),
.B2(n_71),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_90),
.A2(n_92),
.B1(n_99),
.B2(n_58),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_84),
.A2(n_62),
.B1(n_76),
.B2(n_50),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_64),
.Y(n_108)
);

AOI21xp33_ASAP7_75t_SL g97 ( 
.A1(n_78),
.A2(n_54),
.B(n_56),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_97),
.A2(n_56),
.B(n_66),
.C(n_52),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_55),
.B1(n_57),
.B2(n_70),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_100),
.B(n_67),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_89),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_107),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_72),
.B1(n_68),
.B2(n_60),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_110),
.B1(n_112),
.B2(n_113),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_11),
.Y(n_128)
);

HAxp5_ASAP7_75t_SL g133 ( 
.A(n_105),
.B(n_22),
.CON(n_133),
.SN(n_133)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_106),
.B(n_108),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_88),
.A2(n_73),
.B1(n_63),
.B2(n_66),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_1),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_118),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_97),
.A2(n_52),
.B1(n_3),
.B2(n_4),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_91),
.A2(n_93),
.B1(n_101),
.B2(n_94),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_91),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_115),
.A2(n_116),
.B1(n_9),
.B2(n_11),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_93),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_7),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_125),
.A2(n_130),
.B1(n_26),
.B2(n_27),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_128),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_49),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_125),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_46),
.C(n_25),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_137),
.C(n_139),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_124),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_136),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_24),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_140),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_30),
.C(n_35),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_133),
.A2(n_37),
.B(n_39),
.C(n_40),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_126),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_132),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_144),
.B(n_131),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_122),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_149),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_121),
.B(n_120),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_150),
.A2(n_143),
.B(n_141),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_151),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_154),
.B(n_145),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_152),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_148),
.C(n_146),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_157),
.B(n_147),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_158),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_147),
.Y(n_160)
);


endmodule