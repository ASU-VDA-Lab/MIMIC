module real_aes_6359_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_354;
wire n_265;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g169 ( .A1(n_0), .A2(n_170), .B(n_171), .C(n_175), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_1), .B(n_164), .Y(n_177) );
INVx1_ASAP7_75t_L g105 ( .A(n_2), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_3), .B(n_149), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_4), .A2(n_158), .B(n_467), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_5), .A2(n_138), .B(n_155), .C(n_511), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_6), .A2(n_158), .B(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_7), .B(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_8), .B(n_164), .Y(n_473) );
AO21x2_ASAP7_75t_L g251 ( .A1(n_9), .A2(n_130), .B(n_252), .Y(n_251) );
AOI222xp33_ASAP7_75t_L g442 ( .A1(n_10), .A2(n_443), .B1(n_712), .B2(n_715), .C1(n_719), .C2(n_720), .Y(n_442) );
AND2x6_ASAP7_75t_L g155 ( .A(n_11), .B(n_156), .Y(n_155) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_12), .A2(n_138), .B(n_155), .C(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g564 ( .A(n_13), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_14), .B(n_111), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_14), .B(n_41), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_15), .B(n_174), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_16), .A2(n_102), .B1(n_112), .B2(n_725), .Y(n_101) );
INVx1_ASAP7_75t_L g135 ( .A(n_17), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_18), .B(n_149), .Y(n_258) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_19), .A2(n_150), .B(n_522), .C(n_524), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_20), .B(n_164), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_21), .B(n_192), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_L g183 ( .A1(n_22), .A2(n_138), .B(n_184), .C(n_191), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_23), .A2(n_173), .B(n_226), .C(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_24), .B(n_174), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_25), .B(n_174), .Y(n_462) );
CKINVDCx16_ASAP7_75t_R g491 ( .A(n_26), .Y(n_491) );
INVx1_ASAP7_75t_L g461 ( .A(n_27), .Y(n_461) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_28), .A2(n_138), .B(n_191), .C(n_255), .Y(n_254) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_29), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_30), .Y(n_509) );
INVx1_ASAP7_75t_L g485 ( .A(n_31), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_32), .A2(n_158), .B(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g140 ( .A(n_33), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_34), .A2(n_153), .B(n_207), .C(n_208), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_35), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_36), .A2(n_173), .B(n_470), .C(n_472), .Y(n_469) );
INVxp67_ASAP7_75t_L g486 ( .A(n_37), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_38), .B(n_257), .Y(n_256) );
CKINVDCx14_ASAP7_75t_R g468 ( .A(n_39), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g459 ( .A1(n_40), .A2(n_138), .B(n_191), .C(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g111 ( .A(n_41), .Y(n_111) );
A2O1A1Ixp33_ASAP7_75t_L g561 ( .A1(n_42), .A2(n_175), .B(n_562), .C(n_563), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_43), .B(n_182), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_44), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_45), .B(n_149), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_46), .B(n_158), .Y(n_253) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_47), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_48), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_49), .A2(n_153), .B(n_207), .C(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g172 ( .A(n_50), .Y(n_172) );
INVx1_ASAP7_75t_L g236 ( .A(n_51), .Y(n_236) );
INVx1_ASAP7_75t_L g529 ( .A(n_52), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_53), .B(n_158), .Y(n_233) );
OAI22xp5_ASAP7_75t_SL g120 ( .A1(n_54), .A2(n_71), .B1(n_121), .B2(n_122), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_54), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_55), .Y(n_196) );
CKINVDCx14_ASAP7_75t_R g560 ( .A(n_56), .Y(n_560) );
INVx1_ASAP7_75t_L g156 ( .A(n_57), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_58), .B(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_59), .B(n_164), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_60), .A2(n_145), .B(n_190), .C(n_247), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_61), .A2(n_70), .B1(n_713), .B2(n_714), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_61), .Y(n_713) );
INVx1_ASAP7_75t_L g134 ( .A(n_62), .Y(n_134) );
INVx1_ASAP7_75t_SL g471 ( .A(n_63), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_64), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_65), .B(n_149), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_66), .B(n_164), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_67), .B(n_150), .Y(n_223) );
INVx1_ASAP7_75t_L g494 ( .A(n_68), .Y(n_494) );
CKINVDCx16_ASAP7_75t_R g167 ( .A(n_69), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_70), .Y(n_714) );
INVx1_ASAP7_75t_L g122 ( .A(n_71), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_72), .B(n_186), .Y(n_185) );
A2O1A1Ixp33_ASAP7_75t_L g137 ( .A1(n_73), .A2(n_138), .B(n_143), .C(n_153), .Y(n_137) );
CKINVDCx16_ASAP7_75t_R g245 ( .A(n_74), .Y(n_245) );
INVx1_ASAP7_75t_L g109 ( .A(n_75), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_76), .A2(n_158), .B(n_559), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_77), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_78), .A2(n_158), .B(n_519), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_79), .A2(n_182), .B(n_481), .Y(n_480) );
CKINVDCx16_ASAP7_75t_R g458 ( .A(n_80), .Y(n_458) );
INVx1_ASAP7_75t_L g520 ( .A(n_81), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_82), .B(n_188), .Y(n_187) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_83), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_84), .A2(n_158), .B(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g523 ( .A(n_85), .Y(n_523) );
INVx2_ASAP7_75t_L g132 ( .A(n_86), .Y(n_132) );
INVx1_ASAP7_75t_L g512 ( .A(n_87), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_88), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_89), .B(n_174), .Y(n_224) );
INVx2_ASAP7_75t_L g106 ( .A(n_90), .Y(n_106) );
OR2x2_ASAP7_75t_L g434 ( .A(n_90), .B(n_435), .Y(n_434) );
OR2x2_ASAP7_75t_L g447 ( .A(n_90), .B(n_436), .Y(n_447) );
A2O1A1Ixp33_ASAP7_75t_L g492 ( .A1(n_91), .A2(n_138), .B(n_153), .C(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_92), .B(n_158), .Y(n_205) );
INVx1_ASAP7_75t_L g209 ( .A(n_93), .Y(n_209) );
INVxp67_ASAP7_75t_L g248 ( .A(n_94), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_95), .B(n_130), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_96), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g144 ( .A(n_97), .Y(n_144) );
INVx1_ASAP7_75t_L g219 ( .A(n_98), .Y(n_219) );
INVx2_ASAP7_75t_L g532 ( .A(n_99), .Y(n_532) );
AND2x2_ASAP7_75t_L g238 ( .A(n_100), .B(n_194), .Y(n_238) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g726 ( .A(n_103), .Y(n_726) );
OR2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_110), .Y(n_103) );
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_105), .B(n_106), .C(n_107), .Y(n_104) );
AND2x2_ASAP7_75t_L g436 ( .A(n_105), .B(n_437), .Y(n_436) );
OR2x2_ASAP7_75t_L g711 ( .A(n_106), .B(n_436), .Y(n_711) );
NOR2x2_ASAP7_75t_L g722 ( .A(n_106), .B(n_435), .Y(n_722) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
OA21x2_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_118), .B(n_441), .Y(n_112) );
BUFx2_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_SL g724 ( .A(n_116), .Y(n_724) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI21xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_433), .B(n_438), .Y(n_118) );
XNOR2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_123), .Y(n_119) );
INVx1_ASAP7_75t_L g444 ( .A(n_123), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_123), .A2(n_449), .B1(n_716), .B2(n_717), .Y(n_715) );
OR3x1_ASAP7_75t_L g123 ( .A(n_124), .B(n_341), .C(n_390), .Y(n_123) );
NAND5xp2_ASAP7_75t_L g124 ( .A(n_125), .B(n_275), .C(n_304), .D(n_312), .E(n_327), .Y(n_124) );
O2A1O1Ixp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_198), .B(n_214), .C(n_259), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_127), .B(n_178), .Y(n_126) );
AND2x2_ASAP7_75t_L g270 ( .A(n_127), .B(n_267), .Y(n_270) );
AND2x2_ASAP7_75t_L g303 ( .A(n_127), .B(n_179), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_127), .B(n_202), .Y(n_396) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_163), .Y(n_127) );
INVx2_ASAP7_75t_L g201 ( .A(n_128), .Y(n_201) );
BUFx2_ASAP7_75t_L g370 ( .A(n_128), .Y(n_370) );
AO21x2_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_136), .B(n_161), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_129), .B(n_162), .Y(n_161) );
INVx3_ASAP7_75t_L g164 ( .A(n_129), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_129), .B(n_213), .Y(n_212) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_129), .A2(n_218), .B(n_228), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_129), .B(n_464), .Y(n_463) );
AO21x2_ASAP7_75t_L g489 ( .A1(n_129), .A2(n_490), .B(n_497), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_129), .B(n_515), .Y(n_514) );
INVx4_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_130), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_130), .A2(n_253), .B(n_254), .Y(n_252) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g230 ( .A(n_131), .Y(n_230) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
AND2x2_ASAP7_75t_SL g194 ( .A(n_132), .B(n_133), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_157), .Y(n_136) );
INVx5_ASAP7_75t_L g168 ( .A(n_138), .Y(n_168) );
AND2x6_ASAP7_75t_L g138 ( .A(n_139), .B(n_141), .Y(n_138) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_139), .Y(n_152) );
BUFx3_ASAP7_75t_L g176 ( .A(n_139), .Y(n_176) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g160 ( .A(n_140), .Y(n_160) );
INVx1_ASAP7_75t_L g227 ( .A(n_140), .Y(n_227) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_142), .Y(n_147) );
INVx3_ASAP7_75t_L g150 ( .A(n_142), .Y(n_150) );
AND2x2_ASAP7_75t_L g159 ( .A(n_142), .B(n_160), .Y(n_159) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_142), .Y(n_174) );
INVx1_ASAP7_75t_L g257 ( .A(n_142), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_145), .B(n_148), .C(n_151), .Y(n_143) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
OAI22xp33_ASAP7_75t_L g484 ( .A1(n_146), .A2(n_149), .B1(n_485), .B2(n_486), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_146), .B(n_523), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_146), .B(n_532), .Y(n_531) );
INVx4_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g186 ( .A(n_147), .Y(n_186) );
INVx2_ASAP7_75t_L g170 ( .A(n_149), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_149), .B(n_248), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_L g460 ( .A1(n_149), .A2(n_189), .B(n_461), .C(n_462), .Y(n_460) );
INVx5_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_150), .B(n_564), .Y(n_563) );
HB1xp67_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx3_ASAP7_75t_L g472 ( .A(n_152), .Y(n_472) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
O2A1O1Ixp33_ASAP7_75t_SL g166 ( .A1(n_154), .A2(n_167), .B(n_168), .C(n_169), .Y(n_166) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_154), .A2(n_168), .B(n_245), .C(n_246), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_L g467 ( .A1(n_154), .A2(n_168), .B(n_468), .C(n_469), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_SL g481 ( .A1(n_154), .A2(n_168), .B(n_482), .C(n_483), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_SL g519 ( .A1(n_154), .A2(n_168), .B(n_520), .C(n_521), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_SL g528 ( .A1(n_154), .A2(n_168), .B(n_529), .C(n_530), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_SL g559 ( .A1(n_154), .A2(n_168), .B(n_560), .C(n_561), .Y(n_559) );
INVx4_ASAP7_75t_SL g154 ( .A(n_155), .Y(n_154) );
AND2x4_ASAP7_75t_L g158 ( .A(n_155), .B(n_159), .Y(n_158) );
BUFx3_ASAP7_75t_L g191 ( .A(n_155), .Y(n_191) );
NAND2x1p5_ASAP7_75t_L g220 ( .A(n_155), .B(n_159), .Y(n_220) );
BUFx2_ASAP7_75t_L g182 ( .A(n_158), .Y(n_182) );
INVx1_ASAP7_75t_L g190 ( .A(n_160), .Y(n_190) );
AND2x2_ASAP7_75t_L g178 ( .A(n_163), .B(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g268 ( .A(n_163), .Y(n_268) );
AND2x2_ASAP7_75t_L g354 ( .A(n_163), .B(n_267), .Y(n_354) );
AND2x2_ASAP7_75t_L g409 ( .A(n_163), .B(n_201), .Y(n_409) );
OA21x2_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_165), .B(n_177), .Y(n_163) );
INVx2_ASAP7_75t_L g207 ( .A(n_168), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_172), .B(n_173), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_173), .B(n_471), .Y(n_470) );
INVx4_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g562 ( .A(n_174), .Y(n_562) );
INVx2_ASAP7_75t_L g496 ( .A(n_175), .Y(n_496) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_176), .Y(n_211) );
INVx1_ASAP7_75t_L g524 ( .A(n_176), .Y(n_524) );
INVx1_ASAP7_75t_L g326 ( .A(n_178), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_178), .B(n_202), .Y(n_373) );
INVx5_ASAP7_75t_L g267 ( .A(n_179), .Y(n_267) );
AND2x4_ASAP7_75t_L g288 ( .A(n_179), .B(n_268), .Y(n_288) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_179), .Y(n_310) );
AND2x2_ASAP7_75t_L g385 ( .A(n_179), .B(n_370), .Y(n_385) );
AND2x2_ASAP7_75t_L g388 ( .A(n_179), .B(n_203), .Y(n_388) );
OR2x6_ASAP7_75t_L g179 ( .A(n_180), .B(n_195), .Y(n_179) );
AOI21xp5_ASAP7_75t_SL g180 ( .A1(n_181), .A2(n_183), .B(n_192), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_187), .B(n_189), .Y(n_184) );
INVx2_ASAP7_75t_L g188 ( .A(n_186), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g208 ( .A1(n_188), .A2(n_209), .B(n_210), .C(n_211), .Y(n_208) );
O2A1O1Ixp33_ASAP7_75t_L g235 ( .A1(n_188), .A2(n_211), .B(n_236), .C(n_237), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_188), .A2(n_494), .B(n_495), .C(n_496), .Y(n_493) );
O2A1O1Ixp5_ASAP7_75t_L g511 ( .A1(n_188), .A2(n_496), .B(n_512), .C(n_513), .Y(n_511) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_190), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_193), .B(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx1_ASAP7_75t_L g197 ( .A(n_194), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_194), .A2(n_205), .B(n_206), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_194), .A2(n_233), .B(n_234), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g457 ( .A1(n_194), .A2(n_220), .B(n_458), .C(n_459), .Y(n_457) );
OA21x2_ASAP7_75t_L g557 ( .A1(n_194), .A2(n_558), .B(n_565), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_197), .A2(n_508), .B(n_514), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_198), .B(n_268), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_198), .B(n_399), .Y(n_398) );
INVx2_ASAP7_75t_SL g198 ( .A(n_199), .Y(n_198) );
OR2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_202), .Y(n_199) );
AND2x2_ASAP7_75t_L g293 ( .A(n_200), .B(n_268), .Y(n_293) );
AND2x2_ASAP7_75t_L g311 ( .A(n_200), .B(n_203), .Y(n_311) );
INVx1_ASAP7_75t_L g331 ( .A(n_200), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_200), .B(n_267), .Y(n_376) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_200), .Y(n_418) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_201), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_202), .B(n_266), .Y(n_265) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_202), .Y(n_320) );
O2A1O1Ixp33_ASAP7_75t_L g323 ( .A1(n_202), .A2(n_263), .B(n_324), .C(n_326), .Y(n_323) );
AND2x2_ASAP7_75t_L g330 ( .A(n_202), .B(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g339 ( .A(n_202), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g343 ( .A(n_202), .B(n_267), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_202), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g358 ( .A(n_202), .B(n_268), .Y(n_358) );
AND2x2_ASAP7_75t_L g408 ( .A(n_202), .B(n_409), .Y(n_408) );
INVx5_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
BUFx2_ASAP7_75t_L g272 ( .A(n_203), .Y(n_272) );
AND2x2_ASAP7_75t_L g313 ( .A(n_203), .B(n_266), .Y(n_313) );
AND2x2_ASAP7_75t_L g325 ( .A(n_203), .B(n_300), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_203), .B(n_354), .Y(n_372) );
OR2x6_ASAP7_75t_L g203 ( .A(n_204), .B(n_212), .Y(n_203) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_239), .Y(n_214) );
INVx1_ASAP7_75t_L g261 ( .A(n_215), .Y(n_261) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_231), .Y(n_215) );
OR2x2_ASAP7_75t_L g263 ( .A(n_216), .B(n_231), .Y(n_263) );
NAND3xp33_ASAP7_75t_L g269 ( .A(n_216), .B(n_270), .C(n_271), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_216), .B(n_241), .Y(n_280) );
OR2x2_ASAP7_75t_L g295 ( .A(n_216), .B(n_283), .Y(n_295) );
AND2x2_ASAP7_75t_L g301 ( .A(n_216), .B(n_250), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_216), .B(n_432), .Y(n_431) );
INVx5_ASAP7_75t_SL g216 ( .A(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_217), .B(n_241), .Y(n_298) );
AND2x2_ASAP7_75t_L g337 ( .A(n_217), .B(n_251), .Y(n_337) );
NAND2xp5_ASAP7_75t_SL g365 ( .A(n_217), .B(n_250), .Y(n_365) );
OR2x2_ASAP7_75t_L g368 ( .A(n_217), .B(n_250), .Y(n_368) );
OAI21xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_221), .Y(n_218) );
OAI21xp5_ASAP7_75t_L g490 ( .A1(n_220), .A2(n_491), .B(n_492), .Y(n_490) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_220), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_225), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_225), .A2(n_256), .B(n_258), .Y(n_255) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
INVx2_ASAP7_75t_L g479 ( .A(n_230), .Y(n_479) );
INVx5_ASAP7_75t_SL g283 ( .A(n_231), .Y(n_283) );
OR2x2_ASAP7_75t_L g289 ( .A(n_231), .B(n_240), .Y(n_289) );
AND2x2_ASAP7_75t_L g305 ( .A(n_231), .B(n_306), .Y(n_305) );
AOI321xp33_ASAP7_75t_L g312 ( .A1(n_231), .A2(n_313), .A3(n_314), .B1(n_315), .B2(n_321), .C(n_323), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_231), .B(n_239), .Y(n_322) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_231), .Y(n_335) );
OR2x2_ASAP7_75t_L g382 ( .A(n_231), .B(n_280), .Y(n_382) );
AND2x2_ASAP7_75t_L g404 ( .A(n_231), .B(n_301), .Y(n_404) );
AND2x2_ASAP7_75t_L g423 ( .A(n_231), .B(n_241), .Y(n_423) );
OR2x6_ASAP7_75t_L g231 ( .A(n_232), .B(n_238), .Y(n_231) );
INVx1_ASAP7_75t_SL g239 ( .A(n_240), .Y(n_239) );
OR2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_250), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_241), .B(n_250), .Y(n_264) );
AND2x2_ASAP7_75t_L g273 ( .A(n_241), .B(n_274), .Y(n_273) );
INVx3_ASAP7_75t_L g300 ( .A(n_241), .Y(n_300) );
AND2x2_ASAP7_75t_L g306 ( .A(n_241), .B(n_301), .Y(n_306) );
INVxp67_ASAP7_75t_L g336 ( .A(n_241), .Y(n_336) );
OR2x2_ASAP7_75t_L g378 ( .A(n_241), .B(n_283), .Y(n_378) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B(n_249), .Y(n_241) );
OA21x2_ASAP7_75t_L g465 ( .A1(n_242), .A2(n_466), .B(n_473), .Y(n_465) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_242), .A2(n_518), .B(n_525), .Y(n_517) );
OA21x2_ASAP7_75t_L g526 ( .A1(n_242), .A2(n_527), .B(n_533), .Y(n_526) );
OR2x2_ASAP7_75t_L g260 ( .A(n_250), .B(n_261), .Y(n_260) );
INVx1_ASAP7_75t_SL g274 ( .A(n_250), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_250), .B(n_263), .Y(n_307) );
AND2x2_ASAP7_75t_L g356 ( .A(n_250), .B(n_300), .Y(n_356) );
AND2x2_ASAP7_75t_L g394 ( .A(n_250), .B(n_283), .Y(n_394) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_251), .B(n_283), .Y(n_282) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_262), .B(n_265), .C(n_269), .Y(n_259) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_260), .A2(n_262), .B1(n_387), .B2(n_389), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_262), .A2(n_285), .B1(n_340), .B2(n_426), .Y(n_425) );
OR2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx1_ASAP7_75t_SL g414 ( .A(n_263), .Y(n_414) );
INVx1_ASAP7_75t_SL g314 ( .A(n_264), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_266), .B(n_286), .Y(n_316) );
AOI222xp33_ASAP7_75t_L g327 ( .A1(n_266), .A2(n_307), .B1(n_314), .B2(n_328), .C1(n_332), .C2(n_338), .Y(n_327) );
AND2x2_ASAP7_75t_L g417 ( .A(n_266), .B(n_418), .Y(n_417) );
AND2x4_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVx2_ASAP7_75t_L g292 ( .A(n_267), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_267), .B(n_287), .Y(n_362) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_267), .Y(n_399) );
AND2x2_ASAP7_75t_L g402 ( .A(n_267), .B(n_311), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_267), .B(n_418), .Y(n_428) );
INVx1_ASAP7_75t_L g319 ( .A(n_268), .Y(n_319) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_268), .Y(n_347) );
O2A1O1Ixp33_ASAP7_75t_L g410 ( .A1(n_270), .A2(n_411), .B(n_412), .C(n_415), .Y(n_410) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
NAND3xp33_ASAP7_75t_L g333 ( .A(n_272), .B(n_334), .C(n_337), .Y(n_333) );
OR2x2_ASAP7_75t_L g361 ( .A(n_272), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_272), .B(n_288), .Y(n_389) );
OR2x2_ASAP7_75t_L g294 ( .A(n_274), .B(n_295), .Y(n_294) );
AOI211xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_278), .B(n_284), .C(n_296), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_277), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g383 ( .A(n_278), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_279), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g297 ( .A(n_282), .B(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_283), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g351 ( .A(n_283), .B(n_301), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_283), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_283), .B(n_300), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_289), .B1(n_290), .B2(n_294), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_286), .B(n_358), .Y(n_357) );
BUFx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_288), .B(n_330), .Y(n_329) );
OAI221xp5_ASAP7_75t_SL g352 ( .A1(n_289), .A2(n_353), .B1(n_355), .B2(n_357), .C(n_359), .Y(n_352) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
AND2x2_ASAP7_75t_L g407 ( .A(n_292), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g420 ( .A(n_292), .B(n_409), .Y(n_420) );
INVx1_ASAP7_75t_L g340 ( .A(n_293), .Y(n_340) );
INVx1_ASAP7_75t_L g411 ( .A(n_294), .Y(n_411) );
AOI21xp5_ASAP7_75t_L g400 ( .A1(n_295), .A2(n_378), .B(n_401), .Y(n_400) );
AOI21xp33_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_299), .B(n_302), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OAI21xp5_ASAP7_75t_SL g304 ( .A1(n_305), .A2(n_307), .B(n_308), .Y(n_304) );
INVx1_ASAP7_75t_L g344 ( .A(n_305), .Y(n_344) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_306), .A2(n_392), .B1(n_395), .B2(n_397), .C(n_400), .Y(n_391) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_314), .A2(n_404), .B1(n_405), .B2(n_407), .Y(n_403) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx1_ASAP7_75t_L g380 ( .A(n_316), .Y(n_380) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NOR2xp67_ASAP7_75t_SL g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AND2x2_ASAP7_75t_L g384 ( .A(n_320), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g349 ( .A(n_325), .Y(n_349) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_330), .B(n_354), .Y(n_406) );
INVxp67_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_336), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g422 ( .A(n_337), .B(n_423), .Y(n_422) );
AND2x4_ASAP7_75t_L g429 ( .A(n_337), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OAI211xp5_ASAP7_75t_SL g341 ( .A1(n_342), .A2(n_344), .B(n_345), .C(n_379), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AOI211xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_348), .B(n_352), .C(n_371), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_SL g432 ( .A(n_356), .Y(n_432) );
AND2x2_ASAP7_75t_L g369 ( .A(n_358), .B(n_370), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_363), .B1(n_367), .B2(n_369), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
OR2x2_ASAP7_75t_L g377 ( .A(n_365), .B(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g430 ( .A(n_366), .Y(n_430) );
INVxp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AOI31xp33_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_373), .A3(n_374), .B(n_377), .Y(n_371) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AOI211xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_381), .B(n_383), .C(n_386), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
CKINVDCx16_ASAP7_75t_R g387 ( .A(n_388), .Y(n_387) );
NAND5xp2_ASAP7_75t_L g390 ( .A(n_391), .B(n_403), .C(n_410), .D(n_424), .E(n_427), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g427 ( .A1(n_402), .A2(n_428), .B1(n_429), .B2(n_431), .Y(n_427) );
INVx1_ASAP7_75t_SL g426 ( .A(n_404), .Y(n_426) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AOI21xp33_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_419), .B(n_421), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVxp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_434), .Y(n_440) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NAND3xp33_ASAP7_75t_L g441 ( .A(n_438), .B(n_442), .C(n_723), .Y(n_441) );
INVx1_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
OAI22xp5_ASAP7_75t_SL g443 ( .A1(n_444), .A2(n_445), .B1(n_448), .B2(n_711), .Y(n_443) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g716 ( .A(n_446), .Y(n_716) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OR3x1_ASAP7_75t_L g449 ( .A(n_450), .B(n_622), .C(n_669), .Y(n_449) );
NAND3xp33_ASAP7_75t_SL g450 ( .A(n_451), .B(n_568), .C(n_593), .Y(n_450) );
AOI221xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_506), .B1(n_534), .B2(n_537), .C(n_545), .Y(n_451) );
OAI21xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_474), .B(n_499), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_454), .B(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_454), .B(n_550), .Y(n_666) );
AND2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_465), .Y(n_454) );
AND2x2_ASAP7_75t_L g536 ( .A(n_455), .B(n_505), .Y(n_536) );
AND2x2_ASAP7_75t_L g586 ( .A(n_455), .B(n_504), .Y(n_586) );
AND2x2_ASAP7_75t_L g607 ( .A(n_455), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g612 ( .A(n_455), .B(n_579), .Y(n_612) );
OR2x2_ASAP7_75t_L g620 ( .A(n_455), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g692 ( .A(n_455), .B(n_488), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_455), .B(n_641), .Y(n_706) );
INVx3_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g551 ( .A(n_456), .B(n_465), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_456), .B(n_488), .Y(n_552) );
AND2x4_ASAP7_75t_L g574 ( .A(n_456), .B(n_505), .Y(n_574) );
AND2x2_ASAP7_75t_L g604 ( .A(n_456), .B(n_476), .Y(n_604) );
AND2x2_ASAP7_75t_L g613 ( .A(n_456), .B(n_603), .Y(n_613) );
AND2x2_ASAP7_75t_L g629 ( .A(n_456), .B(n_489), .Y(n_629) );
OR2x2_ASAP7_75t_L g638 ( .A(n_456), .B(n_621), .Y(n_638) );
AND2x2_ASAP7_75t_L g644 ( .A(n_456), .B(n_579), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_456), .B(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g658 ( .A(n_456), .B(n_501), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_456), .B(n_547), .Y(n_668) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_456), .B(n_608), .Y(n_697) );
OR2x6_ASAP7_75t_L g456 ( .A(n_457), .B(n_463), .Y(n_456) );
INVx2_ASAP7_75t_L g505 ( .A(n_465), .Y(n_505) );
AND2x2_ASAP7_75t_L g603 ( .A(n_465), .B(n_488), .Y(n_603) );
AND2x2_ASAP7_75t_L g608 ( .A(n_465), .B(n_489), .Y(n_608) );
INVx1_ASAP7_75t_L g664 ( .A(n_465), .Y(n_664) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g573 ( .A(n_475), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_488), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_476), .B(n_536), .Y(n_535) );
BUFx3_ASAP7_75t_L g550 ( .A(n_476), .Y(n_550) );
OR2x2_ASAP7_75t_L g621 ( .A(n_476), .B(n_488), .Y(n_621) );
OR2x2_ASAP7_75t_L g682 ( .A(n_476), .B(n_589), .Y(n_682) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_480), .B(n_487), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_478), .A2(n_502), .B(n_503), .Y(n_501) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g502 ( .A(n_480), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_487), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_488), .B(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g641 ( .A(n_488), .B(n_501), .Y(n_641) );
INVx2_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
BUFx2_ASAP7_75t_L g580 ( .A(n_489), .Y(n_580) );
INVx1_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_500), .A2(n_686), .B1(n_690), .B2(n_693), .C(n_694), .Y(n_685) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_504), .Y(n_500) );
INVx1_ASAP7_75t_SL g548 ( .A(n_501), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_501), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g680 ( .A(n_501), .B(n_536), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_504), .B(n_550), .Y(n_672) );
AND2x2_ASAP7_75t_L g579 ( .A(n_505), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_SL g583 ( .A(n_506), .Y(n_583) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_506), .B(n_589), .Y(n_619) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_516), .Y(n_506) );
AND2x2_ASAP7_75t_L g544 ( .A(n_507), .B(n_517), .Y(n_544) );
INVx4_ASAP7_75t_L g556 ( .A(n_507), .Y(n_556) );
BUFx3_ASAP7_75t_L g599 ( .A(n_507), .Y(n_599) );
AND3x2_ASAP7_75t_L g614 ( .A(n_507), .B(n_615), .C(n_616), .Y(n_614) );
AND2x2_ASAP7_75t_L g696 ( .A(n_516), .B(n_610), .Y(n_696) );
AND2x2_ASAP7_75t_L g704 ( .A(n_516), .B(n_589), .Y(n_704) );
INVx1_ASAP7_75t_SL g709 ( .A(n_516), .Y(n_709) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_526), .Y(n_516) );
INVx1_ASAP7_75t_SL g567 ( .A(n_517), .Y(n_567) );
AND2x2_ASAP7_75t_L g590 ( .A(n_517), .B(n_556), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_517), .B(n_540), .Y(n_592) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_517), .Y(n_632) );
OR2x2_ASAP7_75t_L g637 ( .A(n_517), .B(n_556), .Y(n_637) );
INVx2_ASAP7_75t_L g542 ( .A(n_526), .Y(n_542) );
AND2x2_ASAP7_75t_L g577 ( .A(n_526), .B(n_557), .Y(n_577) );
OR2x2_ASAP7_75t_L g597 ( .A(n_526), .B(n_557), .Y(n_597) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_526), .Y(n_617) );
INVx1_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
AOI21xp33_ASAP7_75t_L g667 ( .A1(n_535), .A2(n_576), .B(n_668), .Y(n_667) );
AOI322xp5_ASAP7_75t_L g703 ( .A1(n_537), .A2(n_547), .A3(n_574), .B1(n_704), .B2(n_705), .C1(n_707), .C2(n_710), .Y(n_703) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_543), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_539), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_540), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g566 ( .A(n_541), .B(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g634 ( .A(n_542), .B(n_556), .Y(n_634) );
AND2x2_ASAP7_75t_L g701 ( .A(n_542), .B(n_557), .Y(n_701) );
INVx1_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g642 ( .A(n_544), .B(n_596), .Y(n_642) );
AOI31xp33_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_549), .A3(n_552), .B(n_553), .Y(n_545) );
AND2x2_ASAP7_75t_L g601 ( .A(n_547), .B(n_579), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_547), .B(n_571), .Y(n_683) );
AND2x2_ASAP7_75t_L g702 ( .A(n_547), .B(n_607), .Y(n_702) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_550), .B(n_579), .Y(n_591) );
NAND2x1p5_ASAP7_75t_L g625 ( .A(n_550), .B(n_608), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g628 ( .A(n_550), .B(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_550), .B(n_692), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_551), .B(n_608), .Y(n_640) );
INVx1_ASAP7_75t_L g684 ( .A(n_551), .Y(n_684) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_566), .Y(n_554) );
INVxp67_ASAP7_75t_L g636 ( .A(n_555), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_556), .B(n_567), .Y(n_572) );
INVx1_ASAP7_75t_L g678 ( .A(n_556), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_556), .B(n_655), .Y(n_689) );
BUFx3_ASAP7_75t_L g589 ( .A(n_557), .Y(n_589) );
AND2x2_ASAP7_75t_L g615 ( .A(n_557), .B(n_567), .Y(n_615) );
INVx2_ASAP7_75t_L g655 ( .A(n_557), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_566), .B(n_688), .Y(n_687) );
AOI211xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_573), .B(n_575), .C(n_584), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AOI21xp33_ASAP7_75t_L g618 ( .A1(n_570), .A2(n_619), .B(n_620), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_571), .B(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_571), .B(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OR2x2_ASAP7_75t_L g651 ( .A(n_572), .B(n_597), .Y(n_651) );
INVx3_ASAP7_75t_L g582 ( .A(n_574), .Y(n_582) );
OAI22xp5_ASAP7_75t_SL g575 ( .A1(n_576), .A2(n_578), .B1(n_581), .B2(n_583), .Y(n_575) );
OAI21xp5_ASAP7_75t_SL g600 ( .A1(n_577), .A2(n_601), .B(n_602), .Y(n_600) );
AND2x2_ASAP7_75t_L g626 ( .A(n_577), .B(n_590), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_577), .B(n_678), .Y(n_677) );
INVxp67_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g581 ( .A(n_580), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g650 ( .A(n_580), .Y(n_650) );
OAI21xp5_ASAP7_75t_SL g594 ( .A1(n_581), .A2(n_595), .B(n_600), .Y(n_594) );
OAI22xp33_ASAP7_75t_SL g584 ( .A1(n_585), .A2(n_587), .B1(n_591), .B2(n_592), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_586), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx1_ASAP7_75t_L g610 ( .A(n_589), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_589), .B(n_632), .Y(n_631) );
NOR3xp33_ASAP7_75t_L g593 ( .A(n_594), .B(n_605), .C(n_618), .Y(n_593) );
OAI22xp5_ASAP7_75t_SL g660 ( .A1(n_595), .A2(n_661), .B1(n_665), .B2(n_666), .Y(n_660) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_596), .B(n_598), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g665 ( .A(n_597), .B(n_598), .Y(n_665) );
AND2x2_ASAP7_75t_L g673 ( .A(n_598), .B(n_654), .Y(n_673) );
CKINVDCx16_ASAP7_75t_R g598 ( .A(n_599), .Y(n_598) );
O2A1O1Ixp33_ASAP7_75t_SL g681 ( .A1(n_599), .A2(n_682), .B(n_683), .C(n_684), .Y(n_681) );
OR2x2_ASAP7_75t_L g708 ( .A(n_599), .B(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
OAI21xp33_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_609), .B(n_611), .Y(n_605) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
O2A1O1Ixp33_ASAP7_75t_L g643 ( .A1(n_607), .A2(n_644), .B(n_645), .C(n_648), .Y(n_643) );
OAI21xp33_ASAP7_75t_SL g611 ( .A1(n_612), .A2(n_613), .B(n_614), .Y(n_611) );
AND2x2_ASAP7_75t_L g676 ( .A(n_615), .B(n_634), .Y(n_676) );
INVxp67_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g654 ( .A(n_617), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g659 ( .A(n_619), .Y(n_659) );
NAND3xp33_ASAP7_75t_SL g622 ( .A(n_623), .B(n_643), .C(n_656), .Y(n_622) );
AOI211xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_626), .B(n_627), .C(n_635), .Y(n_623) );
INVx1_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_628), .B(n_630), .Y(n_627) );
INVx1_ASAP7_75t_L g693 ( .A(n_630), .Y(n_693) );
OR2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
INVx1_ASAP7_75t_L g653 ( .A(n_632), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_632), .B(n_701), .Y(n_700) );
INVxp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
A2O1A1Ixp33_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .B(n_638), .C(n_639), .Y(n_635) );
INVx2_ASAP7_75t_SL g647 ( .A(n_637), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_638), .A2(n_649), .B1(n_651), .B2(n_652), .Y(n_648) );
OAI21xp33_ASAP7_75t_SL g639 ( .A1(n_640), .A2(n_641), .B(n_642), .Y(n_639) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
AOI211xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_659), .B(n_660), .C(n_667), .Y(n_656) );
INVx1_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
INVxp33_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g710 ( .A(n_664), .Y(n_710) );
NAND4xp25_ASAP7_75t_L g669 ( .A(n_670), .B(n_685), .C(n_698), .D(n_703), .Y(n_669) );
AOI211xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_673), .B(n_674), .C(n_681), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_677), .B(n_679), .Y(n_674) );
AOI21xp33_ASAP7_75t_L g694 ( .A1(n_675), .A2(n_695), .B(n_697), .Y(n_694) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_682), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_702), .Y(n_698) );
INVxp67_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g718 ( .A(n_711), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_712), .Y(n_719) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
INVx3_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
endmodule