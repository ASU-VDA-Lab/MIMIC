module fake_aes_6882_n_29 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_29);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_29;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
AND3x2_ASAP7_75t_L g13 ( .A(n_3), .B(n_11), .C(n_6), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_5), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_9), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_2), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_1), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_10), .B(n_0), .Y(n_18) );
NAND3xp33_ASAP7_75t_L g19 ( .A(n_16), .B(n_4), .C(n_7), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_16), .Y(n_20) );
OAI21x1_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_14), .B(n_17), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
NOR3xp33_ASAP7_75t_L g27 ( .A(n_26), .B(n_19), .C(n_15), .Y(n_27) );
AO22x1_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_18), .B1(n_0), .B2(n_13), .Y(n_28) );
OAI21xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_8), .B(n_12), .Y(n_29) );
endmodule