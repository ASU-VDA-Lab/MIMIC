module fake_ibex_278_n_34 (n_4, n_2, n_7, n_5, n_11, n_6, n_8, n_10, n_0, n_9, n_3, n_1, n_34);

input n_4;
input n_2;
input n_7;
input n_5;
input n_11;
input n_6;
input n_8;
input n_10;
input n_0;
input n_9;
input n_3;
input n_1;

output n_34;

wire n_20;
wire n_17;
wire n_25;
wire n_18;
wire n_28;
wire n_22;
wire n_32;
wire n_33;
wire n_30;
wire n_29;
wire n_13;
wire n_26;
wire n_14;
wire n_12;
wire n_15;
wire n_24;
wire n_31;
wire n_23;
wire n_21;
wire n_27;
wire n_19;
wire n_16;

NAND2xp33_ASAP7_75t_SL g12 ( 
.A(n_4),
.B(n_10),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_11),
.B(n_8),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_0),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_1),
.B(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

OAI21x1_ASAP7_75t_L g22 ( 
.A1(n_13),
.A2(n_14),
.B(n_15),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

OAI21x1_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_20),
.B(n_21),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_12),
.A2(n_19),
.B(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_16),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_17),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_23),
.Y(n_31)
);

AOI211xp5_ASAP7_75t_SL g32 ( 
.A1(n_31),
.A2(n_25),
.B(n_29),
.C(n_27),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_33),
.A2(n_30),
.B(n_22),
.Y(n_34)
);


endmodule