module fake_jpeg_2918_n_613 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_613);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_613;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_14),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx5_ASAP7_75t_SL g164 ( 
.A(n_58),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_29),
.B(n_10),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_59),
.B(n_73),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_60),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_61),
.Y(n_188)
);

BUFx4f_ASAP7_75t_SL g62 ( 
.A(n_46),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_62),
.Y(n_160)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_64),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_65),
.Y(n_210)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_68),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_10),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_69),
.B(n_76),
.Y(n_140)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_29),
.B(n_42),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_21),
.B(n_9),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_75),
.B(n_102),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_20),
.B(n_18),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_77),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_78),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_79),
.Y(n_165)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_81),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_82),
.Y(n_185)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_83),
.Y(n_189)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_84),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_86),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_87),
.Y(n_186)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_88),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_89),
.Y(n_193)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_90),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_91),
.Y(n_202)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_22),
.Y(n_92)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_92),
.Y(n_221)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_95),
.Y(n_168)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g197 ( 
.A(n_96),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_97),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g204 ( 
.A(n_98),
.Y(n_204)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_26),
.Y(n_99)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_99),
.Y(n_190)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_100),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_31),
.B(n_9),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_103),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_38),
.B(n_9),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_104),
.B(n_116),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_24),
.A2(n_44),
.B1(n_52),
.B2(n_55),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_105),
.A2(n_30),
.B1(n_43),
.B2(n_39),
.Y(n_174)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_24),
.Y(n_106)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_106),
.Y(n_159)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_107),
.Y(n_209)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_26),
.Y(n_108)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_108),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_109),
.Y(n_196)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_110),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_24),
.Y(n_111)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_111),
.Y(n_161)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_112),
.Y(n_173)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_38),
.Y(n_113)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_26),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_26),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_115),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_20),
.B(n_11),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_34),
.Y(n_117)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_117),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_26),
.Y(n_118)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_118),
.Y(n_179)
);

INVx6_ASAP7_75t_SL g119 ( 
.A(n_47),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_119),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_49),
.Y(n_120)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_120),
.Y(n_181)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_121),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_49),
.Y(n_122)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_122),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_42),
.B(n_11),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_123),
.B(n_13),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_49),
.Y(n_124)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_124),
.Y(n_195)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_49),
.Y(n_125)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_125),
.Y(n_201)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_49),
.Y(n_126)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_126),
.Y(n_214)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_53),
.Y(n_127)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_127),
.Y(n_216)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_53),
.Y(n_128)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_128),
.Y(n_218)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_136),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_77),
.A2(n_29),
.B1(n_51),
.B2(n_33),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g240 ( 
.A1(n_143),
.A2(n_158),
.B1(n_171),
.B2(n_175),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_73),
.B(n_45),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_144),
.B(n_154),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_97),
.B(n_55),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_145),
.B(n_147),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_59),
.B(n_25),
.Y(n_147)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_67),
.Y(n_153)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_153),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_85),
.B(n_25),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_111),
.Y(n_155)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_155),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_107),
.B(n_41),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_157),
.B(n_162),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_117),
.A2(n_41),
.B1(n_51),
.B2(n_33),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_118),
.B(n_40),
.Y(n_162)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_112),
.Y(n_166)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_166),
.Y(n_257)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_101),
.Y(n_169)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_169),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_77),
.A2(n_30),
.B1(n_40),
.B2(n_43),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_174),
.A2(n_8),
.B1(n_164),
.B2(n_210),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_63),
.A2(n_39),
.B1(n_27),
.B2(n_32),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_84),
.Y(n_178)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_178),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_64),
.B(n_27),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_192),
.B(n_200),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_62),
.B(n_13),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_203),
.B(n_220),
.Y(n_250)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_120),
.Y(n_205)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_205),
.Y(n_283)
);

AND2x4_ASAP7_75t_SL g207 ( 
.A(n_58),
.B(n_47),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_L g223 ( 
.A1(n_207),
.A2(n_211),
.B(n_32),
.Y(n_223)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_122),
.Y(n_208)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_208),
.Y(n_289)
);

NAND2x1p5_ASAP7_75t_L g211 ( 
.A(n_124),
.B(n_32),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_82),
.A2(n_32),
.B1(n_47),
.B2(n_34),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_212),
.A2(n_60),
.B1(n_54),
.B2(n_19),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_87),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_213),
.B(n_217),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_78),
.B(n_32),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_89),
.B(n_12),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_222),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g342 ( 
.A(n_223),
.Y(n_342)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_130),
.Y(n_224)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_224),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_217),
.A2(n_91),
.B1(n_98),
.B2(n_81),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_225),
.A2(n_232),
.B1(n_243),
.B2(n_265),
.Y(n_340)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_148),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_227),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_228),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_144),
.A2(n_109),
.B1(n_114),
.B2(n_99),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_229),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_149),
.A2(n_109),
.B1(n_88),
.B2(n_92),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_230),
.A2(n_231),
.B1(n_233),
.B2(n_235),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_149),
.A2(n_96),
.B1(n_86),
.B2(n_79),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_L g232 ( 
.A1(n_143),
.A2(n_171),
.B1(n_175),
.B2(n_173),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_154),
.A2(n_71),
.B1(n_65),
.B2(n_61),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_131),
.Y(n_234)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_234),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_133),
.B(n_134),
.C(n_140),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_236),
.B(n_246),
.C(n_251),
.Y(n_322)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_163),
.Y(n_238)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_238),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_156),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_239),
.Y(n_305)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_160),
.Y(n_241)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_241),
.Y(n_347)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_138),
.Y(n_242)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_242),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_212),
.A2(n_54),
.B1(n_19),
.B2(n_2),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_141),
.Y(n_244)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_244),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_216),
.A2(n_54),
.B1(n_19),
.B2(n_12),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_245),
.A2(n_253),
.B1(n_259),
.B2(n_262),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_180),
.B(n_18),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_179),
.Y(n_247)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_247),
.Y(n_324)
);

AND2x2_ASAP7_75t_SL g249 ( 
.A(n_218),
.B(n_192),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_249),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_129),
.B(n_18),
.C(n_17),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_159),
.A2(n_17),
.B1(n_16),
.B2(n_15),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_152),
.B(n_0),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_254),
.B(n_256),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_152),
.B(n_1),
.Y(n_256)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_206),
.Y(n_258)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_258),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_147),
.A2(n_17),
.B1(n_14),
.B2(n_13),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_221),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_260),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_211),
.B(n_1),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_261),
.B(n_273),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_161),
.A2(n_17),
.B1(n_11),
.B2(n_3),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_151),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_263),
.A2(n_266),
.B1(n_280),
.B2(n_287),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_177),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_264),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_185),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_189),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_266)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_181),
.Y(n_270)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_270),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_139),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_271),
.A2(n_278),
.B1(n_146),
.B2(n_190),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_201),
.B(n_5),
.Y(n_273)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_188),
.Y(n_274)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_274),
.Y(n_337)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_194),
.Y(n_275)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_275),
.Y(n_345)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_160),
.Y(n_276)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_276),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_207),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_277),
.B(n_291),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_132),
.A2(n_6),
.B1(n_8),
.B2(n_209),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_191),
.A2(n_198),
.B1(n_210),
.B2(n_188),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_160),
.Y(n_281)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_281),
.Y(n_308)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_197),
.Y(n_282)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_282),
.Y(n_313)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_195),
.Y(n_284)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_284),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_187),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_285),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_135),
.B(n_6),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_286),
.B(n_204),
.C(n_137),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_214),
.B(n_176),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_288),
.B(n_296),
.Y(n_321)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_197),
.Y(n_290)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_290),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_170),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_164),
.B(n_8),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_292),
.B(n_167),
.Y(n_325)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_219),
.Y(n_293)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_293),
.Y(n_331)
);

OAI22xp33_ASAP7_75t_L g294 ( 
.A1(n_185),
.A2(n_193),
.B1(n_186),
.B2(n_184),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_294),
.A2(n_150),
.B1(n_165),
.B2(n_184),
.Y(n_349)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_197),
.Y(n_295)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_295),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_215),
.B(n_193),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_142),
.Y(n_297)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_297),
.Y(n_350)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_182),
.Y(n_298)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_298),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_146),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_299),
.B(n_237),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_223),
.A2(n_168),
.B(n_196),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_307),
.A2(n_298),
.B(n_281),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_261),
.A2(n_183),
.B(n_199),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_312),
.A2(n_339),
.B(n_301),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_288),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_318),
.B(n_335),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_323),
.A2(n_349),
.B1(n_336),
.B2(n_301),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_325),
.B(n_357),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_L g328 ( 
.A1(n_272),
.A2(n_294),
.B1(n_296),
.B2(n_232),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_328),
.A2(n_343),
.B1(n_286),
.B2(n_274),
.Y(n_377)
);

A2O1A1Ixp33_ASAP7_75t_L g332 ( 
.A1(n_226),
.A2(n_172),
.B(n_186),
.C(n_202),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_332),
.B(n_240),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_255),
.B(n_172),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_333),
.B(n_352),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_239),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_260),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_338),
.B(n_258),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_250),
.B(n_137),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_341),
.B(n_222),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_L g343 ( 
.A1(n_252),
.A2(n_202),
.B1(n_150),
.B2(n_165),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_348),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_236),
.B(n_204),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_353),
.B(n_243),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_246),
.B(n_204),
.C(n_249),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_355),
.B(n_286),
.C(n_273),
.Y(n_367)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_224),
.Y(n_356)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_356),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_269),
.B(n_256),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_359),
.B(n_367),
.C(n_381),
.Y(n_414)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_360),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_303),
.B(n_254),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_361),
.B(n_366),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_340),
.A2(n_287),
.B1(n_250),
.B2(n_249),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_362),
.A2(n_388),
.B1(n_396),
.B2(n_326),
.Y(n_405)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_319),
.Y(n_364)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_364),
.Y(n_419)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_319),
.Y(n_365)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_365),
.Y(n_420)
);

FAx1_ASAP7_75t_SL g366 ( 
.A(n_355),
.B(n_267),
.CI(n_225),
.CON(n_366),
.SN(n_366)
);

CKINVDCx6p67_ASAP7_75t_R g368 ( 
.A(n_335),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_368),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_344),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_369),
.B(n_350),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_303),
.B(n_248),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_370),
.B(n_331),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_371),
.A2(n_393),
.B1(n_326),
.B2(n_354),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_322),
.B(n_240),
.C(n_257),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_372),
.B(n_375),
.C(n_389),
.Y(n_412)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_356),
.Y(n_373)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_373),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_L g374 ( 
.A1(n_310),
.A2(n_268),
.B1(n_279),
.B2(n_289),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_374),
.A2(n_378),
.B1(n_392),
.B2(n_354),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_322),
.B(n_306),
.C(n_342),
.Y(n_375)
);

OR2x2_ASAP7_75t_L g376 ( 
.A(n_307),
.B(n_240),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_376),
.A2(n_313),
.B(n_330),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_377),
.B(n_399),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_340),
.A2(n_240),
.B1(n_265),
.B2(n_244),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_351),
.Y(n_379)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_379),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_341),
.B(n_251),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_382),
.B(n_383),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_318),
.B(n_283),
.Y(n_383)
);

NAND2xp33_ASAP7_75t_SL g436 ( 
.A(n_384),
.B(n_387),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_321),
.B(n_270),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_385),
.B(n_386),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_321),
.B(n_275),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_332),
.B(n_336),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_346),
.A2(n_317),
.B1(n_353),
.B2(n_311),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_317),
.B(n_242),
.C(n_234),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_312),
.B(n_247),
.C(n_284),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_390),
.B(n_398),
.C(n_331),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_309),
.B(n_293),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_391),
.B(n_395),
.Y(n_438)
);

AOI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_349),
.A2(n_241),
.B1(n_276),
.B2(n_227),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_309),
.B(n_282),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_323),
.A2(n_264),
.B1(n_290),
.B2(n_295),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_338),
.B(n_238),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_397),
.B(n_400),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_350),
.B(n_339),
.C(n_334),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_300),
.B(n_302),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_314),
.Y(n_401)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_401),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_378),
.A2(n_371),
.B1(n_376),
.B2(n_387),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_403),
.A2(n_415),
.B1(n_416),
.B2(n_360),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_404),
.A2(n_407),
.B(n_384),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_405),
.A2(n_434),
.B1(n_397),
.B2(n_365),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_395),
.B(n_351),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_406),
.B(n_409),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_376),
.A2(n_387),
.B(n_399),
.Y(n_407)
);

OAI22x1_ASAP7_75t_L g469 ( 
.A1(n_408),
.A2(n_305),
.B1(n_304),
.B2(n_373),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_400),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_411),
.B(n_417),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_382),
.A2(n_337),
.B1(n_314),
.B2(n_327),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_383),
.A2(n_337),
.B1(n_314),
.B2(n_327),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_368),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_421),
.B(n_389),
.Y(n_454)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_363),
.Y(n_427)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_427),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_375),
.B(n_330),
.C(n_313),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_428),
.B(n_437),
.C(n_398),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_429),
.B(n_302),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_368),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_430),
.B(n_431),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_369),
.B(n_334),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_L g442 ( 
.A1(n_432),
.A2(n_377),
.B1(n_390),
.B2(n_359),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_362),
.A2(n_327),
.B1(n_308),
.B2(n_300),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_363),
.Y(n_435)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_435),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_381),
.B(n_308),
.Y(n_437)
);

OAI21xp33_ASAP7_75t_L g482 ( 
.A1(n_440),
.A2(n_466),
.B(n_470),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_442),
.A2(n_445),
.B1(n_446),
.B2(n_448),
.Y(n_501)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_419),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_443),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_436),
.A2(n_358),
.B(n_388),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_444),
.A2(n_453),
.B(n_465),
.Y(n_499)
);

AOI22x1_ASAP7_75t_L g445 ( 
.A1(n_403),
.A2(n_396),
.B1(n_368),
.B2(n_391),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_405),
.A2(n_372),
.B1(n_358),
.B2(n_394),
.Y(n_448)
);

INVxp33_ASAP7_75t_L g497 ( 
.A(n_449),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_414),
.B(n_367),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_450),
.B(n_468),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_413),
.B(n_386),
.Y(n_452)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_452),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_436),
.A2(n_361),
.B(n_366),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_454),
.B(n_455),
.C(n_457),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_414),
.B(n_437),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_431),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_456),
.B(n_463),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g458 ( 
.A(n_407),
.Y(n_458)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_458),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_412),
.B(n_385),
.C(n_366),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_461),
.B(n_464),
.C(n_428),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_404),
.Y(n_462)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_462),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_439),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_412),
.B(n_370),
.C(n_402),
.Y(n_464)
);

FAx1_ASAP7_75t_SL g465 ( 
.A(n_424),
.B(n_380),
.CI(n_402),
.CON(n_465),
.SN(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_413),
.B(n_368),
.Y(n_466)
);

AOI22x1_ASAP7_75t_L g467 ( 
.A1(n_410),
.A2(n_432),
.B1(n_418),
.B2(n_438),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_467),
.A2(n_469),
.B1(n_473),
.B2(n_433),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_412),
.B(n_380),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_438),
.B(n_364),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_471),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_437),
.B(n_315),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_472),
.B(n_422),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_434),
.A2(n_401),
.B1(n_304),
.B2(n_305),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_446),
.A2(n_410),
.B1(n_409),
.B2(n_423),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_477),
.A2(n_479),
.B1(n_480),
.B2(n_487),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_478),
.B(n_470),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_462),
.A2(n_410),
.B1(n_466),
.B2(n_441),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_448),
.A2(n_410),
.B1(n_408),
.B2(n_423),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_440),
.A2(n_418),
.B(n_424),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_481),
.A2(n_490),
.B(n_493),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_455),
.B(n_428),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_483),
.B(n_484),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_450),
.B(n_421),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_457),
.B(n_421),
.C(n_406),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_486),
.B(n_494),
.C(n_459),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_458),
.A2(n_439),
.B1(n_411),
.B2(n_417),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_444),
.A2(n_433),
.B(n_430),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_SL g491 ( 
.A(n_461),
.B(n_435),
.Y(n_491)
);

MAJx2_ASAP7_75t_L g509 ( 
.A(n_491),
.B(n_492),
.C(n_496),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_454),
.B(n_425),
.C(n_427),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_SL g496 ( 
.A(n_453),
.B(n_422),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_468),
.B(n_429),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_500),
.B(n_502),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_464),
.B(n_425),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_472),
.B(n_420),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_503),
.B(n_504),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_452),
.B(n_420),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_474),
.Y(n_505)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_505),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_498),
.A2(n_467),
.B(n_451),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_506),
.A2(n_479),
.B(n_477),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_500),
.B(n_447),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_507),
.B(n_518),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_508),
.B(n_510),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_476),
.B(n_451),
.C(n_441),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_512),
.B(n_513),
.C(n_521),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_476),
.B(n_447),
.C(n_467),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_487),
.Y(n_514)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_514),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_486),
.B(n_419),
.Y(n_518)
);

OR2x2_ASAP7_75t_L g519 ( 
.A(n_481),
.B(n_465),
.Y(n_519)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_519),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_504),
.B(n_443),
.Y(n_520)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_520),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_488),
.B(n_445),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_488),
.B(n_445),
.C(n_460),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_522),
.B(n_524),
.C(n_525),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_483),
.B(n_469),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_484),
.B(n_460),
.C(n_433),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_502),
.B(n_465),
.Y(n_526)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_526),
.Y(n_546)
);

NAND2x1_ASAP7_75t_L g527 ( 
.A(n_490),
.B(n_416),
.Y(n_527)
);

XNOR2x1_ASAP7_75t_L g547 ( 
.A(n_527),
.B(n_530),
.Y(n_547)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_495),
.Y(n_528)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_528),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_478),
.B(n_415),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_529),
.B(n_503),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_SL g530 ( 
.A(n_491),
.B(n_315),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_511),
.A2(n_497),
.B1(n_501),
.B2(n_480),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_532),
.A2(n_533),
.B1(n_538),
.B2(n_542),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_511),
.A2(n_497),
.B1(n_482),
.B2(n_485),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g552 ( 
.A1(n_535),
.A2(n_527),
.B(n_516),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_519),
.A2(n_489),
.B1(n_475),
.B2(n_493),
.Y(n_538)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_520),
.Y(n_540)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_540),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_506),
.A2(n_495),
.B1(n_494),
.B2(n_492),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_516),
.A2(n_499),
.B1(n_496),
.B2(n_426),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_543),
.B(n_548),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_521),
.A2(n_524),
.B1(n_522),
.B2(n_513),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_550),
.A2(n_515),
.B1(n_517),
.B2(n_508),
.Y(n_558)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_552),
.B(n_563),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_537),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_SL g574 ( 
.A1(n_553),
.A2(n_545),
.B1(n_546),
.B2(n_540),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_531),
.B(n_544),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_SL g571 ( 
.A(n_554),
.B(n_555),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_531),
.B(n_512),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_534),
.B(n_510),
.C(n_515),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_556),
.B(n_549),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_536),
.B(n_528),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_557),
.B(n_566),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_558),
.B(n_562),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_541),
.B(n_529),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_560),
.B(n_548),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_SL g561 ( 
.A1(n_535),
.A2(n_527),
.B(n_525),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_SL g567 ( 
.A1(n_561),
.A2(n_543),
.B(n_533),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_549),
.B(n_517),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_536),
.B(n_523),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_539),
.A2(n_523),
.B1(n_530),
.B2(n_509),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_565),
.A2(n_542),
.B1(n_550),
.B2(n_547),
.Y(n_575)
);

FAx1_ASAP7_75t_SL g566 ( 
.A(n_534),
.B(n_509),
.CI(n_426),
.CON(n_566),
.SN(n_566)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_567),
.B(n_316),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_SL g583 ( 
.A(n_569),
.B(n_556),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_570),
.B(n_574),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_552),
.A2(n_547),
.B(n_532),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_572),
.A2(n_559),
.B1(n_565),
.B2(n_563),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_575),
.A2(n_576),
.B1(n_577),
.B2(n_559),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_557),
.B(n_401),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_564),
.A2(n_347),
.B1(n_320),
.B2(n_324),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_SL g578 ( 
.A(n_551),
.B(n_347),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_578),
.B(n_561),
.Y(n_584)
);

FAx1_ASAP7_75t_SL g579 ( 
.A(n_566),
.B(n_320),
.CI(n_316),
.CON(n_579),
.SN(n_579)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_579),
.B(n_345),
.Y(n_590)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_581),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g582 ( 
.A(n_568),
.B(n_551),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_582),
.B(n_573),
.C(n_580),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_583),
.B(n_585),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_584),
.B(n_590),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_571),
.B(n_562),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_SL g598 ( 
.A1(n_586),
.A2(n_591),
.B(n_567),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_568),
.B(n_558),
.C(n_566),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_588),
.B(n_589),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_573),
.B(n_553),
.C(n_324),
.Y(n_589)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_594),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_SL g596 ( 
.A(n_587),
.B(n_571),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_596),
.B(n_598),
.Y(n_602)
);

OAI21xp5_ASAP7_75t_SL g599 ( 
.A1(n_588),
.A2(n_580),
.B(n_570),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_599),
.B(n_584),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_593),
.B(n_582),
.C(n_589),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_L g605 ( 
.A1(n_600),
.A2(n_604),
.B(n_597),
.Y(n_605)
);

O2A1O1Ixp33_ASAP7_75t_SL g606 ( 
.A1(n_603),
.A2(n_595),
.B(n_597),
.C(n_578),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_592),
.B(n_591),
.C(n_576),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_605),
.B(n_600),
.C(n_601),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_606),
.A2(n_607),
.B(n_575),
.Y(n_609)
);

OAI21xp5_ASAP7_75t_SL g607 ( 
.A1(n_602),
.A2(n_572),
.B(n_579),
.Y(n_607)
);

NAND2xp33_ASAP7_75t_SL g610 ( 
.A(n_608),
.B(n_609),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_610),
.B(n_579),
.C(n_329),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_611),
.B(n_329),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_612),
.B(n_345),
.Y(n_613)
);


endmodule