module fake_jpeg_16940_n_369 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_369);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_369;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_40),
.B(n_42),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_19),
.Y(n_43)
);

NAND2x1_ASAP7_75t_SL g110 ( 
.A(n_43),
.B(n_3),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_7),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_45),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_7),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_7),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_23),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_16),
.B(n_18),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_52),
.Y(n_80)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_56),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_21),
.B(n_5),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_59),
.Y(n_90)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_5),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_31),
.Y(n_61)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

CKINVDCx9p33_ASAP7_75t_R g64 ( 
.A(n_33),
.Y(n_64)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_L g92 ( 
.A1(n_66),
.A2(n_8),
.B(n_13),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_68),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_37),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_70),
.B(n_72),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_36),
.B1(n_20),
.B2(n_14),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_71),
.A2(n_74),
.B1(n_108),
.B2(n_109),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_37),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_35),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_73),
.B(n_75),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_52),
.A2(n_14),
.B1(n_20),
.B2(n_29),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_33),
.C(n_34),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_83),
.B(n_85),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_35),
.Y(n_85)
);

OR2x2_ASAP7_75t_SL g86 ( 
.A(n_64),
.B(n_33),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_86),
.A2(n_100),
.B(n_95),
.C(n_114),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_63),
.A2(n_23),
.B1(n_21),
.B2(n_32),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_113),
.B1(n_104),
.B2(n_83),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_43),
.A2(n_34),
.B1(n_26),
.B2(n_24),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_91),
.A2(n_93),
.B1(n_13),
.B2(n_1),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_92),
.A2(n_110),
.B1(n_0),
.B2(n_1),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_43),
.A2(n_26),
.B1(n_24),
.B2(n_8),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_94),
.B(n_118),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_59),
.B(n_5),
.Y(n_96)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_48),
.B(n_42),
.C(n_54),
.Y(n_99)
);

FAx1_ASAP7_75t_SL g144 ( 
.A(n_99),
.B(n_75),
.CI(n_111),
.CON(n_144),
.SN(n_144)
);

AOI21xp33_ASAP7_75t_SL g100 ( 
.A1(n_61),
.A2(n_0),
.B(n_1),
.Y(n_100)
);

BUFx10_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_38),
.B(n_5),
.Y(n_106)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_58),
.B(n_4),
.Y(n_107)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_66),
.A2(n_4),
.B1(n_12),
.B2(n_11),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g109 ( 
.A1(n_62),
.A2(n_9),
.B1(n_12),
.B2(n_11),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_61),
.B(n_3),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_0),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_58),
.B(n_3),
.Y(n_112)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_39),
.A2(n_41),
.B1(n_68),
.B2(n_49),
.Y(n_113)
);

BUFx8_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g132 ( 
.A(n_114),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_47),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_67),
.B(n_9),
.Y(n_119)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_82),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_120),
.B(n_124),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_122),
.B(n_129),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_82),
.Y(n_124)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

INVxp67_ASAP7_75t_SL g195 ( 
.A(n_125),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_83),
.A2(n_53),
.B1(n_55),
.B2(n_12),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_126),
.A2(n_128),
.B1(n_131),
.B2(n_140),
.Y(n_180)
);

AO22x1_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_12),
.B1(n_13),
.B2(n_2),
.Y(n_128)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

AO22x2_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_134),
.B(n_146),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_138),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_139),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_70),
.A2(n_72),
.B1(n_74),
.B2(n_71),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_142),
.B(n_149),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_152),
.C(n_135),
.Y(n_175)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_113),
.A2(n_79),
.B1(n_95),
.B2(n_118),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_147),
.A2(n_165),
.B1(n_169),
.B2(n_155),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_108),
.A2(n_80),
.B1(n_73),
.B2(n_84),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_148),
.A2(n_123),
.B1(n_137),
.B2(n_130),
.Y(n_201)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_89),
.B(n_109),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_152),
.Y(n_182)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_103),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_151),
.B(n_159),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_99),
.B(n_90),
.Y(n_152)
);

AOI32xp33_ASAP7_75t_L g153 ( 
.A1(n_110),
.A2(n_76),
.A3(n_86),
.B1(n_77),
.B2(n_79),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_153),
.A2(n_131),
.B(n_145),
.C(n_143),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_104),
.A2(n_78),
.B1(n_69),
.B2(n_102),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_155),
.A2(n_160),
.B(n_135),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_81),
.A2(n_117),
.B1(n_98),
.B2(n_69),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_156),
.A2(n_158),
.B1(n_125),
.B2(n_166),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_117),
.A2(n_98),
.B1(n_102),
.B2(n_78),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_114),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_87),
.Y(n_162)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_97),
.Y(n_164)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_164),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_101),
.A2(n_97),
.B1(n_105),
.B2(n_116),
.Y(n_165)
);

INVx5_ASAP7_75t_SL g166 ( 
.A(n_114),
.Y(n_166)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_166),
.Y(n_212)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_167),
.Y(n_177)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_101),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_168),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_116),
.A2(n_70),
.B1(n_72),
.B2(n_74),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_160),
.A2(n_135),
.B(n_131),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_171),
.A2(n_173),
.B(n_181),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_191),
.C(n_208),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_157),
.B(n_154),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_176),
.B(n_203),
.Y(n_217)
);

O2A1O1Ixp33_ASAP7_75t_SL g181 ( 
.A1(n_150),
.A2(n_131),
.B(n_128),
.C(n_136),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_183),
.A2(n_188),
.B1(n_178),
.B2(n_170),
.Y(n_237)
);

AND2x4_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_128),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_184),
.B(n_191),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_122),
.A2(n_136),
.B1(n_140),
.B2(n_144),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_189),
.A2(n_190),
.B1(n_206),
.B2(n_184),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_169),
.A2(n_147),
.B1(n_126),
.B2(n_133),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_133),
.B(n_157),
.C(n_134),
.Y(n_191)
);

AO22x2_ASAP7_75t_L g192 ( 
.A1(n_133),
.A2(n_157),
.B1(n_165),
.B2(n_139),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_192),
.A2(n_198),
.B1(n_209),
.B2(n_182),
.Y(n_215)
);

AOI32xp33_ASAP7_75t_L g193 ( 
.A1(n_163),
.A2(n_143),
.A3(n_154),
.B1(n_132),
.B2(n_121),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_190),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_141),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_200),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_162),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_200),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_204),
.A2(n_205),
.B1(n_179),
.B2(n_178),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_151),
.A2(n_164),
.B1(n_132),
.B2(n_161),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_127),
.A2(n_150),
.B1(n_122),
.B2(n_136),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_127),
.B(n_144),
.C(n_152),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_142),
.B(n_133),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_209),
.B(n_211),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_160),
.A2(n_135),
.B(n_131),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_210),
.A2(n_171),
.B(n_181),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_149),
.B(n_83),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_213),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_215),
.A2(n_224),
.B(n_234),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_198),
.A2(n_182),
.B1(n_184),
.B2(n_206),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_216),
.A2(n_221),
.B1(n_223),
.B2(n_233),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_218),
.B(n_227),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_175),
.A2(n_192),
.B1(n_183),
.B2(n_208),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_193),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_222),
.B(n_225),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_192),
.A2(n_184),
.B1(n_198),
.B2(n_210),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_184),
.A2(n_192),
.B(n_173),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_203),
.B(n_192),
.Y(n_225)
);

INVxp33_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_239),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_228),
.A2(n_235),
.B(n_243),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_212),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_229),
.B(n_241),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_179),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_238),
.Y(n_264)
);

INVx8_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_172),
.A2(n_188),
.B1(n_181),
.B2(n_180),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_232),
.Y(n_267)
);

OAI21xp33_ASAP7_75t_L g235 ( 
.A1(n_189),
.A2(n_180),
.B(n_212),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_174),
.Y(n_236)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_236),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_237),
.A2(n_232),
.B1(n_238),
.B2(n_222),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_174),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_170),
.Y(n_240)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_240),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_186),
.B(n_177),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_195),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_231),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_197),
.A2(n_186),
.B(n_199),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_199),
.A2(n_207),
.B1(n_202),
.B2(n_177),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_244),
.A2(n_246),
.B1(n_233),
.B2(n_220),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_207),
.A2(n_204),
.B1(n_179),
.B2(n_166),
.Y(n_246)
);

AND2x2_ASAP7_75t_SL g247 ( 
.A(n_202),
.B(n_187),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_249),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_187),
.A2(n_210),
.B(n_171),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_248),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_187),
.B(n_185),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_252),
.A2(n_265),
.B(n_279),
.Y(n_303)
);

O2A1O1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_243),
.A2(n_235),
.B(n_237),
.C(n_224),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_253),
.A2(n_272),
.B(n_259),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_232),
.A2(n_215),
.B1(n_216),
.B2(n_218),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_256),
.A2(n_214),
.B1(n_219),
.B2(n_217),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_260),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_213),
.B(n_249),
.Y(n_262)
);

AND2x6_ASAP7_75t_L g265 ( 
.A(n_223),
.B(n_221),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_236),
.Y(n_266)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_266),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_268),
.A2(n_277),
.B1(n_255),
.B2(n_270),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_229),
.B(n_241),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_246),
.A2(n_228),
.B1(n_234),
.B2(n_218),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_240),
.Y(n_274)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_274),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_239),
.B(n_247),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_278),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_215),
.A2(n_216),
.B1(n_225),
.B2(n_228),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_220),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_244),
.Y(n_279)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_231),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_251),
.Y(n_293)
);

OAI32xp33_ASAP7_75t_L g281 ( 
.A1(n_273),
.A2(n_217),
.A3(n_245),
.B1(n_227),
.B2(n_219),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_281),
.B(n_288),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_267),
.A2(n_248),
.B1(n_214),
.B2(n_245),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_282),
.A2(n_290),
.B1(n_280),
.B2(n_288),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_214),
.Y(n_283)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_283),
.Y(n_313)
);

XNOR2x1_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_248),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_284),
.A2(n_286),
.B(n_291),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_285),
.A2(n_253),
.B1(n_268),
.B2(n_276),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_257),
.B(n_259),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_255),
.B(n_234),
.C(n_247),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_271),
.B(n_234),
.Y(n_289)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_293),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_258),
.B(n_275),
.Y(n_296)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_296),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_250),
.B(n_256),
.Y(n_297)
);

OA21x2_ASAP7_75t_SL g320 ( 
.A1(n_297),
.A2(n_261),
.B(n_251),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_258),
.B(n_264),
.Y(n_298)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_298),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_273),
.B(n_269),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_254),
.B(n_269),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_301),
.B(n_262),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_250),
.C(n_252),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_302),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_303),
.A2(n_305),
.B(n_290),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_278),
.B(n_276),
.C(n_265),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_304),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_253),
.B(n_265),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_306),
.B(n_297),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_291),
.A2(n_260),
.B(n_274),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_307),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_304),
.A2(n_263),
.B1(n_261),
.B2(n_266),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_308),
.A2(n_324),
.B1(n_295),
.B2(n_284),
.Y(n_334)
);

XOR2x2_ASAP7_75t_L g310 ( 
.A(n_284),
.B(n_263),
.Y(n_310)
);

NOR2xp67_ASAP7_75t_SL g328 ( 
.A(n_310),
.B(n_320),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_294),
.Y(n_314)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_314),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_254),
.Y(n_316)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_316),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_317),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_299),
.B(n_280),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_323),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_302),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_325),
.B(n_330),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_328),
.B(n_312),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_309),
.B(n_283),
.Y(n_330)
);

FAx1_ASAP7_75t_SL g331 ( 
.A(n_306),
.B(n_282),
.CI(n_285),
.CON(n_331),
.SN(n_331)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_331),
.B(n_337),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_334),
.A2(n_336),
.B1(n_338),
.B2(n_311),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_312),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_310),
.A2(n_311),
.B1(n_295),
.B2(n_322),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_313),
.B(n_297),
.C(n_289),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_324),
.A2(n_303),
.B1(n_296),
.B2(n_287),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_313),
.B(n_286),
.C(n_305),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_339),
.B(n_306),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_340),
.B(n_341),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_325),
.B(n_308),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_342),
.B(n_344),
.C(n_348),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_327),
.A2(n_310),
.B1(n_315),
.B2(n_300),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g356 ( 
.A(n_343),
.B(n_349),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_329),
.A2(n_326),
.B1(n_332),
.B2(n_333),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_345),
.B(n_350),
.Y(n_351)
);

A2O1A1Ixp33_ASAP7_75t_L g349 ( 
.A1(n_338),
.A2(n_281),
.B(n_318),
.C(n_321),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_339),
.A2(n_300),
.B1(n_319),
.B2(n_315),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_347),
.B(n_330),
.C(n_336),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_354),
.B(n_355),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_346),
.B(n_317),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_356),
.A2(n_307),
.B(n_343),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_358),
.A2(n_349),
.B(n_323),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_353),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_359),
.B(n_360),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_351),
.A2(n_308),
.B1(n_334),
.B2(n_319),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_361),
.B(n_352),
.Y(n_364)
);

AOI21xp33_ASAP7_75t_L g363 ( 
.A1(n_362),
.A2(n_357),
.B(n_358),
.Y(n_363)
);

NOR3xp33_ASAP7_75t_SL g365 ( 
.A(n_363),
.B(n_364),
.C(n_356),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_365),
.B(n_352),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_366),
.B(n_342),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_367),
.B(n_347),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g369 ( 
.A(n_368),
.B(n_331),
.Y(n_369)
);


endmodule