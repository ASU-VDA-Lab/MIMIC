module fake_jpeg_15693_n_46 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_46);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_46;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_7),
.B1(n_17),
.B2(n_16),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_31)
);

OAI32xp33_ASAP7_75t_L g27 ( 
.A1(n_20),
.A2(n_18),
.A3(n_14),
.B1(n_12),
.B2(n_9),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_28)
);

OAI21xp33_ASAP7_75t_L g29 ( 
.A1(n_20),
.A2(n_1),
.B(n_2),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_3),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_22),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_22),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_24),
.C(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_39),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_34),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_31),
.B1(n_4),
.B2(n_5),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_31),
.C(n_38),
.Y(n_42)
);

INVxp67_ASAP7_75t_SL g43 ( 
.A(n_42),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_41),
.Y(n_44)
);

OAI221xp5_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_35),
.B1(n_24),
.B2(n_6),
.C(n_3),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_45),
.B(n_6),
.Y(n_46)
);


endmodule