module fake_jpeg_29769_n_129 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_129);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx4f_ASAP7_75t_SL g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_25),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_39),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_54),
.Y(n_68)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

HAxp5_ASAP7_75t_SL g54 ( 
.A(n_45),
.B(n_0),
.CON(n_54),
.SN(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_60),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_44),
.B1(n_49),
.B2(n_48),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_59),
.A2(n_61),
.B1(n_50),
.B2(n_41),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_52),
.A2(n_42),
.B1(n_37),
.B2(n_46),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_69),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_36),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_40),
.C(n_43),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_70),
.B(n_37),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_68),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_85),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_38),
.B(n_1),
.C(n_2),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_6),
.Y(n_96)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_87),
.B1(n_4),
.B2(n_5),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_23),
.C(n_32),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_0),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_2),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_5),
.Y(n_92)
);

AO22x1_ASAP7_75t_SL g87 ( 
.A1(n_67),
.A2(n_21),
.B1(n_34),
.B2(n_33),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_3),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_7),
.B(n_10),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_92),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_95),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_96),
.B(n_11),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_80),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_81),
.Y(n_103)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_103),
.B(n_105),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_87),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_83),
.B1(n_72),
.B2(n_7),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_106),
.A2(n_94),
.B1(n_13),
.B2(n_18),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_24),
.C(n_8),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_107),
.A2(n_12),
.B(n_20),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_91),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_110),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_109),
.A2(n_98),
.B(n_100),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_89),
.Y(n_112)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

XNOR2x2_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_106),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_107),
.C(n_102),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

OAI322xp33_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_114),
.A3(n_116),
.B1(n_111),
.B2(n_115),
.C1(n_120),
.C2(n_121),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_123),
.Y(n_124)
);

FAx1_ASAP7_75t_SL g125 ( 
.A(n_124),
.B(n_115),
.CI(n_104),
.CON(n_125),
.SN(n_125)
);

OA21x2_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_27),
.B(n_29),
.Y(n_126)
);

INVxp67_ASAP7_75t_SL g127 ( 
.A(n_126),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_125),
.Y(n_129)
);


endmodule