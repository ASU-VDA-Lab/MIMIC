module fake_netlist_6_379_n_1454 (n_52, n_1, n_91, n_326, n_256, n_209, n_63, n_223, n_278, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_56, n_119, n_235, n_147, n_191, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_53, n_44, n_232, n_16, n_163, n_46, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_323, n_152, n_92, n_321, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_325, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_231, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_215, n_178, n_247, n_225, n_308, n_309, n_317, n_149, n_90, n_24, n_54, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_315, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1454);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_323;
input n_152;
input n_92;
input n_321;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_325;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_231;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_317;
input n_149;
input n_90;
input n_24;
input n_54;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1454;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1415;
wire n_1370;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1393;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_976;
wire n_1445;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_527;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1372;
wire n_505;
wire n_1339;
wire n_537;
wire n_1427;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_1429;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1443;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_934;
wire n_482;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_1343;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1416;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1147;
wire n_763;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_1311;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_339;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_241),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_274),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_232),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_202),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_98),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_18),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_306),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_166),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_226),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_301),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_83),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_278),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_161),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_218),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_77),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_176),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_171),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_248),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_158),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_319),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_199),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_73),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_267),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_55),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_116),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_260),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_215),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_220),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_280),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_174),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_52),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_147),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_327),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_196),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_325),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_96),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_193),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_259),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_194),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_216),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g368 ( 
.A(n_326),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_155),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_22),
.Y(n_370)
);

CKINVDCx14_ASAP7_75t_R g371 ( 
.A(n_236),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_234),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_320),
.Y(n_373)
);

BUFx8_ASAP7_75t_SL g374 ( 
.A(n_277),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_146),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_198),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_89),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_109),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_115),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_46),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_239),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_114),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_53),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_318),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_170),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_208),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_137),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_101),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_186),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_184),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_210),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_217),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_279),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_42),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_64),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_125),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_177),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_134),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_293),
.Y(n_399)
);

BUFx10_ASAP7_75t_L g400 ( 
.A(n_15),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_313),
.Y(n_401)
);

INVxp33_ASAP7_75t_L g402 ( 
.A(n_151),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_16),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_74),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_117),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_281),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_3),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_123),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_97),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_192),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_130),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_143),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_70),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_308),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_321),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_225),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_57),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_246),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_175),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_284),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_139),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_133),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_152),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_52),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_10),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_49),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_190),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_162),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_312),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_14),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_261),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_187),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_264),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_163),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_72),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_66),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_296),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_122),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_168),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_42),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_272),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_240),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_237),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_120),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_247),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_31),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_140),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_28),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_221),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_16),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_179),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_93),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_213),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_78),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_4),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_86),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_266),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_164),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_250),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_26),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_297),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_230),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_124),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_63),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_26),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_80),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_289),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_6),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_157),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_282),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_36),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_49),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_22),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_269),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_169),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_54),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_180),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_316),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_324),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_14),
.Y(n_480)
);

BUFx10_ASAP7_75t_L g481 ( 
.A(n_107),
.Y(n_481)
);

BUFx10_ASAP7_75t_L g482 ( 
.A(n_95),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_19),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_276),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_10),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_214),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_189),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_54),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_12),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_283),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_273),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_233),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_67),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_127),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_106),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_191),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_265),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_224),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_211),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_18),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_309),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_118),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_131),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g504 ( 
.A(n_87),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_121),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_58),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_268),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_317),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_185),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_32),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_144),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_270),
.Y(n_512)
);

BUFx8_ASAP7_75t_SL g513 ( 
.A(n_30),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_262),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_229),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_128),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_15),
.Y(n_517)
);

INVx5_ASAP7_75t_L g518 ( 
.A(n_354),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_354),
.Y(n_519)
);

INVx5_ASAP7_75t_L g520 ( 
.A(n_354),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_378),
.B(n_0),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_402),
.B(n_0),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_378),
.B(n_1),
.Y(n_523)
);

BUFx8_ASAP7_75t_SL g524 ( 
.A(n_513),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_455),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_473),
.Y(n_526)
);

INVx5_ASAP7_75t_L g527 ( 
.A(n_354),
.Y(n_527)
);

CKINVDCx11_ASAP7_75t_R g528 ( 
.A(n_400),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_473),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_406),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_342),
.B(n_1),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_406),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_394),
.B(n_2),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_342),
.B(n_2),
.Y(n_534)
);

NAND3xp33_ASAP7_75t_L g535 ( 
.A(n_464),
.B(n_3),
.C(n_4),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_473),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_455),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_513),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_361),
.B(n_5),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_406),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_361),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_406),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_495),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_473),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_417),
.B(n_5),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g546 ( 
.A(n_358),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_371),
.B(n_6),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_400),
.Y(n_548)
);

INVxp33_ASAP7_75t_SL g549 ( 
.A(n_351),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_362),
.B(n_7),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_383),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_362),
.B(n_7),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_389),
.B(n_8),
.Y(n_553)
);

INVx5_ASAP7_75t_L g554 ( 
.A(n_495),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_383),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_389),
.B(n_8),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_408),
.B(n_9),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_402),
.B(n_9),
.Y(n_558)
);

BUFx8_ASAP7_75t_SL g559 ( 
.A(n_374),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_333),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_495),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_380),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_408),
.B(n_11),
.Y(n_563)
);

INVx5_ASAP7_75t_L g564 ( 
.A(n_495),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_504),
.B(n_11),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_481),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_347),
.B(n_12),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_441),
.B(n_13),
.Y(n_568)
);

INVx5_ASAP7_75t_L g569 ( 
.A(n_481),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_395),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_441),
.B(n_13),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_442),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_368),
.B(n_17),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_481),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_400),
.Y(n_575)
);

INVx4_ASAP7_75t_R g576 ( 
.A(n_470),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_442),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_514),
.B(n_332),
.Y(n_578)
);

AND2x6_ASAP7_75t_L g579 ( 
.A(n_514),
.B(n_71),
.Y(n_579)
);

BUFx12f_ASAP7_75t_L g580 ( 
.A(n_482),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_337),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_480),
.B(n_17),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_480),
.B(n_19),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_511),
.B(n_20),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_343),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_403),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_349),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_482),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_353),
.B(n_20),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_407),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_372),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_386),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_446),
.B(n_21),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_448),
.B(n_21),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_450),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_465),
.B(n_23),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_471),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_483),
.B(n_23),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_387),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_482),
.B(n_24),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_374),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_485),
.B(n_24),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_393),
.B(n_25),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_328),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_413),
.B(n_25),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_396),
.B(n_27),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_329),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_424),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_398),
.B(n_27),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_425),
.B(n_28),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_418),
.B(n_29),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_419),
.B(n_29),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_493),
.Y(n_613)
);

INVx5_ASAP7_75t_L g614 ( 
.A(n_330),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_420),
.B(n_30),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_506),
.B(n_510),
.Y(n_616)
);

INVx5_ASAP7_75t_L g617 ( 
.A(n_331),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_428),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_426),
.B(n_31),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_433),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_430),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_435),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_443),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_445),
.Y(n_624)
);

INVx5_ASAP7_75t_L g625 ( 
.A(n_334),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_451),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_454),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_456),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_462),
.B(n_474),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_484),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_486),
.B(n_32),
.Y(n_631)
);

CKINVDCx16_ASAP7_75t_R g632 ( 
.A(n_336),
.Y(n_632)
);

INVxp33_ASAP7_75t_L g633 ( 
.A(n_524),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_526),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_565),
.A2(n_336),
.B1(n_350),
.B2(n_338),
.Y(n_635)
);

OR2x6_ASAP7_75t_L g636 ( 
.A(n_601),
.B(n_494),
.Y(n_636)
);

OAI22xp33_ASAP7_75t_R g637 ( 
.A1(n_546),
.A2(n_558),
.B1(n_522),
.B2(n_584),
.Y(n_637)
);

AOI22x1_ASAP7_75t_L g638 ( 
.A1(n_556),
.A2(n_440),
.B1(n_460),
.B2(n_436),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_529),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_536),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_547),
.A2(n_338),
.B1(n_359),
.B2(n_350),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_544),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_SL g643 ( 
.A1(n_522),
.A2(n_370),
.B1(n_500),
.B2(n_416),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_607),
.B(n_496),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_558),
.A2(n_567),
.B1(n_584),
.B2(n_600),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_574),
.B(n_498),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_621),
.B(n_335),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_572),
.Y(n_648)
);

OAI22xp33_ASAP7_75t_R g649 ( 
.A1(n_546),
.A2(n_500),
.B1(n_370),
.B2(n_503),
.Y(n_649)
);

OAI22xp33_ASAP7_75t_L g650 ( 
.A1(n_574),
.A2(n_472),
.B1(n_476),
.B2(n_468),
.Y(n_650)
);

OAI22xp33_ASAP7_75t_L g651 ( 
.A1(n_535),
.A2(n_489),
.B1(n_517),
.B2(n_488),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_621),
.B(n_339),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_519),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_533),
.A2(n_545),
.B1(n_549),
.B2(n_608),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_605),
.A2(n_416),
.B1(n_432),
.B2(n_359),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_610),
.A2(n_449),
.B1(n_459),
.B2(n_432),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_519),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_519),
.Y(n_658)
);

CKINVDCx6p67_ASAP7_75t_R g659 ( 
.A(n_528),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_530),
.Y(n_660)
);

OAI22xp33_ASAP7_75t_SL g661 ( 
.A1(n_569),
.A2(n_512),
.B1(n_515),
.B2(n_508),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_619),
.A2(n_459),
.B1(n_492),
.B2(n_449),
.Y(n_662)
);

INVx1_ASAP7_75t_SL g663 ( 
.A(n_559),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_548),
.A2(n_502),
.B1(n_492),
.B2(n_352),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_530),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_569),
.B(n_516),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_530),
.Y(n_667)
);

OR2x6_ASAP7_75t_L g668 ( 
.A(n_575),
.B(n_502),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_532),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_SL g670 ( 
.A1(n_632),
.A2(n_344),
.B1(n_341),
.B2(n_340),
.Y(n_670)
);

AO22x2_ASAP7_75t_L g671 ( 
.A1(n_535),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_572),
.Y(n_672)
);

OAI22xp33_ASAP7_75t_SL g673 ( 
.A1(n_569),
.A2(n_346),
.B1(n_348),
.B2(n_345),
.Y(n_673)
);

AO22x2_ASAP7_75t_L g674 ( 
.A1(n_531),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_674)
);

OR2x6_ASAP7_75t_L g675 ( 
.A(n_580),
.B(n_36),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_538),
.A2(n_356),
.B1(n_357),
.B2(n_355),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_532),
.Y(n_677)
);

OAI22xp33_ASAP7_75t_L g678 ( 
.A1(n_631),
.A2(n_363),
.B1(n_364),
.B2(n_360),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_573),
.A2(n_366),
.B1(n_367),
.B2(n_365),
.Y(n_679)
);

AND2x2_ASAP7_75t_SL g680 ( 
.A(n_550),
.B(n_37),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_532),
.Y(n_681)
);

AO22x2_ASAP7_75t_L g682 ( 
.A1(n_531),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_614),
.Y(n_683)
);

OAI22xp33_ASAP7_75t_SL g684 ( 
.A1(n_569),
.A2(n_373),
.B1(n_375),
.B2(n_369),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_541),
.B(n_376),
.Y(n_685)
);

OAI22xp33_ASAP7_75t_SL g686 ( 
.A1(n_521),
.A2(n_379),
.B1(n_381),
.B2(n_377),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_566),
.B(n_382),
.Y(n_687)
);

NAND3x1_ASAP7_75t_L g688 ( 
.A(n_521),
.B(n_38),
.C(n_39),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_589),
.A2(n_438),
.B1(n_507),
.B2(n_505),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_540),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_588),
.A2(n_509),
.B1(n_501),
.B2(n_499),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_540),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_525),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_604),
.B(n_384),
.Y(n_694)
);

OAI22xp33_ASAP7_75t_SL g695 ( 
.A1(n_523),
.A2(n_497),
.B1(n_491),
.B2(n_490),
.Y(n_695)
);

INVx8_ASAP7_75t_L g696 ( 
.A(n_614),
.Y(n_696)
);

OAI22xp33_ASAP7_75t_SL g697 ( 
.A1(n_523),
.A2(n_487),
.B1(n_479),
.B2(n_478),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_604),
.B(n_385),
.Y(n_698)
);

OAI22xp33_ASAP7_75t_L g699 ( 
.A1(n_631),
.A2(n_477),
.B1(n_475),
.B2(n_469),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_534),
.B(n_539),
.Y(n_700)
);

AO22x2_ASAP7_75t_L g701 ( 
.A1(n_534),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_701)
);

AOI22x1_ASAP7_75t_SL g702 ( 
.A1(n_560),
.A2(n_467),
.B1(n_466),
.B2(n_463),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_614),
.B(n_461),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_540),
.Y(n_704)
);

INVx1_ASAP7_75t_SL g705 ( 
.A(n_537),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_609),
.A2(n_458),
.B1(n_457),
.B2(n_453),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_551),
.B(n_388),
.Y(n_707)
);

HB1xp67_ASAP7_75t_L g708 ( 
.A(n_551),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_609),
.A2(n_452),
.B1(n_447),
.B2(n_444),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_539),
.A2(n_412),
.B1(n_437),
.B2(n_434),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_624),
.B(n_390),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_542),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_552),
.A2(n_411),
.B1(n_431),
.B2(n_429),
.Y(n_713)
);

AO22x2_ASAP7_75t_L g714 ( 
.A1(n_552),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_578),
.B(n_391),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_578),
.B(n_392),
.Y(n_716)
);

OAI22xp33_ASAP7_75t_L g717 ( 
.A1(n_553),
.A2(n_439),
.B1(n_427),
.B2(n_423),
.Y(n_717)
);

OR2x2_ASAP7_75t_L g718 ( 
.A(n_629),
.B(n_44),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_542),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_L g720 ( 
.A1(n_553),
.A2(n_422),
.B1(n_421),
.B2(n_415),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_597),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_660),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_700),
.B(n_618),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_660),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_645),
.B(n_556),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_700),
.B(n_627),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_644),
.B(n_603),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_667),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_667),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_648),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_672),
.Y(n_731)
);

NAND2xp33_ASAP7_75t_R g732 ( 
.A(n_668),
.B(n_702),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_647),
.B(n_614),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_653),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_639),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_657),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_707),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_708),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_665),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_665),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_658),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_652),
.B(n_617),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_640),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_634),
.Y(n_744)
);

INVxp33_ASAP7_75t_SL g745 ( 
.A(n_670),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_715),
.B(n_590),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_711),
.B(n_617),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_642),
.Y(n_748)
);

OAI21xp5_ASAP7_75t_L g749 ( 
.A1(n_716),
.A2(n_629),
.B(n_606),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_669),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_721),
.B(n_595),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_677),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_681),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_690),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_692),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_704),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_712),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_705),
.B(n_603),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_706),
.B(n_617),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_702),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_719),
.Y(n_761)
);

INVx1_ASAP7_75t_SL g762 ( 
.A(n_687),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_665),
.Y(n_763)
);

NAND2xp33_ASAP7_75t_R g764 ( 
.A(n_668),
.B(n_644),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_693),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_685),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_718),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_646),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_638),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_636),
.B(n_606),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_683),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_635),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_680),
.B(n_611),
.Y(n_773)
);

AND2x6_ASAP7_75t_L g774 ( 
.A(n_710),
.B(n_557),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_638),
.Y(n_775)
);

XNOR2x2_ASAP7_75t_L g776 ( 
.A(n_674),
.B(n_582),
.Y(n_776)
);

CKINVDCx14_ASAP7_75t_R g777 ( 
.A(n_659),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_694),
.B(n_611),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_698),
.B(n_612),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_683),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_703),
.Y(n_781)
);

XOR2xp5_ASAP7_75t_L g782 ( 
.A(n_643),
.B(n_655),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_666),
.Y(n_783)
);

INVxp33_ASAP7_75t_L g784 ( 
.A(n_656),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_688),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_674),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_682),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_682),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_701),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_701),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_714),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_654),
.B(n_612),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_714),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_717),
.B(n_617),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_671),
.Y(n_795)
);

BUFx8_ASAP7_75t_L g796 ( 
.A(n_649),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_661),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_709),
.Y(n_798)
);

XOR2xp5_ASAP7_75t_L g799 ( 
.A(n_662),
.B(n_597),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_636),
.Y(n_800)
);

NOR3xp33_ASAP7_75t_L g801 ( 
.A(n_651),
.B(n_594),
.C(n_593),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_720),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_671),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_689),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_713),
.B(n_615),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_696),
.A2(n_520),
.B(n_518),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_679),
.Y(n_807)
);

XOR2x2_ASAP7_75t_L g808 ( 
.A(n_664),
.B(n_593),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_696),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_758),
.B(n_641),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_758),
.B(n_615),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_749),
.B(n_557),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_767),
.B(n_778),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_R g814 ( 
.A(n_777),
.B(n_663),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_801),
.A2(n_637),
.B1(n_649),
.B2(n_568),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_777),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_735),
.Y(n_817)
);

HB1xp67_ASAP7_75t_L g818 ( 
.A(n_738),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_778),
.B(n_568),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_768),
.B(n_678),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_779),
.B(n_562),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_735),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_750),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_781),
.B(n_699),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_779),
.B(n_570),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_769),
.B(n_625),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_775),
.B(n_625),
.Y(n_827)
);

OAI21x1_ASAP7_75t_L g828 ( 
.A1(n_747),
.A2(n_571),
.B(n_563),
.Y(n_828)
);

OAI21xp5_ASAP7_75t_L g829 ( 
.A1(n_802),
.A2(n_676),
.B(n_691),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_746),
.B(n_586),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_783),
.B(n_625),
.Y(n_831)
);

INVxp67_ASAP7_75t_L g832 ( 
.A(n_751),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_723),
.B(n_579),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_748),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_733),
.B(n_625),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_746),
.B(n_613),
.Y(n_836)
);

INVx1_ASAP7_75t_SL g837 ( 
.A(n_762),
.Y(n_837)
);

BUFx2_ASAP7_75t_L g838 ( 
.A(n_785),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_748),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_743),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_737),
.B(n_773),
.Y(n_841)
);

INVxp67_ASAP7_75t_SL g842 ( 
.A(n_739),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_739),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_773),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_737),
.B(n_616),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_750),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_743),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_744),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_723),
.B(n_616),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_726),
.B(n_725),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_744),
.Y(n_851)
);

INVxp67_ASAP7_75t_L g852 ( 
.A(n_751),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_726),
.B(n_582),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_807),
.B(n_650),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_742),
.B(n_686),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_804),
.B(n_695),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_725),
.B(n_583),
.Y(n_857)
);

HB1xp67_ASAP7_75t_L g858 ( 
.A(n_785),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_727),
.B(n_583),
.Y(n_859)
);

INVx1_ASAP7_75t_SL g860 ( 
.A(n_792),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_727),
.B(n_594),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_727),
.B(n_697),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_766),
.Y(n_863)
);

HB1xp67_ASAP7_75t_L g864 ( 
.A(n_805),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_797),
.B(n_579),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_722),
.Y(n_866)
);

AND2x4_ASAP7_75t_SL g867 ( 
.A(n_795),
.B(n_675),
.Y(n_867)
);

INVx2_ASAP7_75t_SL g868 ( 
.A(n_734),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_798),
.A2(n_571),
.B(n_563),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_805),
.B(n_572),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_724),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_L g872 ( 
.A1(n_759),
.A2(n_794),
.B(n_792),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_728),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_774),
.B(n_771),
.Y(n_874)
);

AND2x2_ASAP7_75t_SL g875 ( 
.A(n_795),
.B(n_803),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_784),
.B(n_684),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_803),
.B(n_596),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_770),
.B(n_673),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_774),
.B(n_577),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_786),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_793),
.B(n_787),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_774),
.B(n_577),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_729),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_788),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_736),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_770),
.B(n_579),
.Y(n_886)
);

BUFx4_ASAP7_75t_SL g887 ( 
.A(n_760),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_774),
.B(n_577),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_793),
.B(n_789),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_774),
.B(n_579),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_790),
.B(n_596),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_741),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_774),
.B(n_581),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_791),
.B(n_598),
.Y(n_894)
);

AND2x2_ASAP7_75t_SL g895 ( 
.A(n_776),
.B(n_598),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_770),
.B(n_602),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_739),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_784),
.B(n_602),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_730),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_765),
.B(n_675),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_731),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_752),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_771),
.B(n_581),
.Y(n_903)
);

OAI21xp5_ASAP7_75t_L g904 ( 
.A1(n_780),
.A2(n_399),
.B(n_397),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_753),
.Y(n_905)
);

NAND2x1p5_ASAP7_75t_L g906 ( 
.A(n_837),
.B(n_740),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_863),
.B(n_754),
.Y(n_907)
);

INVx2_ASAP7_75t_SL g908 ( 
.A(n_837),
.Y(n_908)
);

AND2x6_ASAP7_75t_L g909 ( 
.A(n_890),
.B(n_776),
.Y(n_909)
);

INVx2_ASAP7_75t_SL g910 ( 
.A(n_818),
.Y(n_910)
);

BUFx4f_ASAP7_75t_L g911 ( 
.A(n_875),
.Y(n_911)
);

OR2x2_ASAP7_75t_L g912 ( 
.A(n_898),
.B(n_860),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_817),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_817),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_812),
.B(n_780),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_812),
.B(n_857),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_846),
.Y(n_917)
);

BUFx4_ASAP7_75t_SL g918 ( 
.A(n_816),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_863),
.B(n_755),
.Y(n_919)
);

BUFx6f_ASAP7_75t_SL g920 ( 
.A(n_900),
.Y(n_920)
);

BUFx2_ASAP7_75t_L g921 ( 
.A(n_864),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_850),
.B(n_756),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_857),
.B(n_808),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_898),
.B(n_808),
.Y(n_924)
);

BUFx12f_ASAP7_75t_L g925 ( 
.A(n_900),
.Y(n_925)
);

AND2x2_ASAP7_75t_SL g926 ( 
.A(n_895),
.B(n_815),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_848),
.Y(n_927)
);

NAND2x1p5_ASAP7_75t_L g928 ( 
.A(n_841),
.B(n_740),
.Y(n_928)
);

NAND2x1p5_ASAP7_75t_L g929 ( 
.A(n_841),
.B(n_809),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_853),
.B(n_757),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_843),
.Y(n_931)
);

OR2x6_ASAP7_75t_L g932 ( 
.A(n_838),
.B(n_800),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_848),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_845),
.B(n_799),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_860),
.Y(n_935)
);

OR2x6_ASAP7_75t_L g936 ( 
.A(n_838),
.B(n_809),
.Y(n_936)
);

NAND2x1p5_ASAP7_75t_L g937 ( 
.A(n_886),
.B(n_761),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_845),
.B(n_799),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_853),
.B(n_763),
.Y(n_939)
);

INVx1_ASAP7_75t_SL g940 ( 
.A(n_813),
.Y(n_940)
);

CKINVDCx16_ASAP7_75t_R g941 ( 
.A(n_814),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_849),
.B(n_782),
.Y(n_942)
);

CKINVDCx14_ASAP7_75t_R g943 ( 
.A(n_900),
.Y(n_943)
);

BUFx2_ASAP7_75t_L g944 ( 
.A(n_844),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_843),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_817),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_850),
.B(n_886),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_886),
.B(n_739),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_859),
.B(n_739),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_810),
.B(n_782),
.Y(n_950)
);

OR2x6_ASAP7_75t_L g951 ( 
.A(n_810),
.B(n_633),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_859),
.B(n_401),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_849),
.B(n_772),
.Y(n_953)
);

INVx6_ASAP7_75t_L g954 ( 
.A(n_900),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_846),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_822),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_861),
.B(n_404),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_861),
.B(n_405),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_811),
.B(n_409),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_813),
.B(n_772),
.Y(n_960)
);

INVx6_ASAP7_75t_L g961 ( 
.A(n_830),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_886),
.B(n_760),
.Y(n_962)
);

NOR2x1_ASAP7_75t_R g963 ( 
.A(n_856),
.B(n_410),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_822),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_846),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_832),
.B(n_555),
.Y(n_966)
);

NAND2x1_ASAP7_75t_SL g967 ( 
.A(n_865),
.B(n_745),
.Y(n_967)
);

NAND2x1p5_ASAP7_75t_L g968 ( 
.A(n_848),
.B(n_851),
.Y(n_968)
);

OR2x6_ASAP7_75t_L g969 ( 
.A(n_862),
.B(n_764),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_822),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_854),
.B(n_745),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_843),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_852),
.B(n_555),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_830),
.Y(n_974)
);

AO21x2_ASAP7_75t_L g975 ( 
.A1(n_874),
.A2(n_806),
.B(n_637),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_811),
.B(n_414),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_836),
.B(n_75),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_836),
.B(n_76),
.Y(n_978)
);

NAND2x1p5_ASAP7_75t_L g979 ( 
.A(n_851),
.B(n_542),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_SL g980 ( 
.A(n_895),
.B(n_796),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_851),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_896),
.B(n_576),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_839),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_918),
.Y(n_984)
);

INVx1_ASAP7_75t_SL g985 ( 
.A(n_908),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_911),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_927),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_927),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_933),
.Y(n_989)
);

BUFx12f_ASAP7_75t_L g990 ( 
.A(n_925),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_983),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_912),
.B(n_895),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_983),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_911),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_933),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_931),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_L g997 ( 
.A1(n_926),
.A2(n_815),
.B1(n_869),
.B2(n_796),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_910),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_916),
.B(n_974),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_961),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_961),
.Y(n_1001)
);

BUFx2_ASAP7_75t_SL g1002 ( 
.A(n_920),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_944),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_913),
.Y(n_1004)
);

BUFx5_ASAP7_75t_L g1005 ( 
.A(n_947),
.Y(n_1005)
);

NAND2x1_ASAP7_75t_L g1006 ( 
.A(n_981),
.B(n_843),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_931),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_931),
.Y(n_1008)
);

BUFx4_ASAP7_75t_SL g1009 ( 
.A(n_932),
.Y(n_1009)
);

BUFx5_ASAP7_75t_L g1010 ( 
.A(n_947),
.Y(n_1010)
);

INVx4_ASAP7_75t_L g1011 ( 
.A(n_945),
.Y(n_1011)
);

BUFx3_ASAP7_75t_L g1012 ( 
.A(n_921),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_922),
.B(n_896),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_909),
.A2(n_869),
.B1(n_796),
.B2(n_829),
.Y(n_1014)
);

NAND2x1p5_ASAP7_75t_L g1015 ( 
.A(n_948),
.B(n_843),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_945),
.Y(n_1016)
);

BUFx12f_ASAP7_75t_L g1017 ( 
.A(n_962),
.Y(n_1017)
);

INVx4_ASAP7_75t_L g1018 ( 
.A(n_945),
.Y(n_1018)
);

INVx8_ASAP7_75t_L g1019 ( 
.A(n_948),
.Y(n_1019)
);

INVx5_ASAP7_75t_SL g1020 ( 
.A(n_932),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_960),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_954),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_939),
.B(n_820),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_953),
.B(n_819),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_935),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_913),
.Y(n_1026)
);

INVx1_ASAP7_75t_SL g1027 ( 
.A(n_934),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_954),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_981),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_972),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_930),
.B(n_877),
.Y(n_1031)
);

BUFx12f_ASAP7_75t_L g1032 ( 
.A(n_962),
.Y(n_1032)
);

CKINVDCx11_ASAP7_75t_R g1033 ( 
.A(n_941),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_914),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_914),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_946),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_924),
.B(n_819),
.Y(n_1037)
);

BUFx12f_ASAP7_75t_L g1038 ( 
.A(n_951),
.Y(n_1038)
);

INVx2_ASAP7_75t_SL g1039 ( 
.A(n_906),
.Y(n_1039)
);

AOI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_971),
.A2(n_876),
.B1(n_872),
.B2(n_824),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_967),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_929),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_946),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_922),
.B(n_881),
.Y(n_1044)
);

INVx3_ASAP7_75t_L g1045 ( 
.A(n_972),
.Y(n_1045)
);

INVx3_ASAP7_75t_L g1046 ( 
.A(n_972),
.Y(n_1046)
);

CKINVDCx14_ASAP7_75t_R g1047 ( 
.A(n_943),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_977),
.B(n_881),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_977),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_1003),
.Y(n_1050)
);

BUFx2_ASAP7_75t_SL g1051 ( 
.A(n_1003),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_1040),
.B(n_978),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_997),
.A2(n_923),
.B1(n_909),
.B2(n_980),
.Y(n_1053)
);

BUFx3_ASAP7_75t_L g1054 ( 
.A(n_1012),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_1012),
.Y(n_1055)
);

BUFx10_ASAP7_75t_L g1056 ( 
.A(n_984),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_991),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_993),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_L g1059 ( 
.A1(n_997),
.A2(n_909),
.B1(n_975),
.B2(n_969),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_984),
.Y(n_1060)
);

BUFx4f_ASAP7_75t_SL g1061 ( 
.A(n_990),
.Y(n_1061)
);

OAI21xp5_ASAP7_75t_SL g1062 ( 
.A1(n_1014),
.A2(n_938),
.B(n_942),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_987),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_SL g1064 ( 
.A1(n_1014),
.A2(n_950),
.B1(n_941),
.B2(n_951),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_987),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_1023),
.B(n_909),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1004),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_988),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_985),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1026),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_996),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1031),
.B(n_875),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1034),
.Y(n_1073)
);

OAI22xp33_ASAP7_75t_L g1074 ( 
.A1(n_992),
.A2(n_940),
.B1(n_969),
.B2(n_732),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_SL g1075 ( 
.A1(n_992),
.A2(n_982),
.B1(n_978),
.B2(n_920),
.Y(n_1075)
);

OR2x2_ASAP7_75t_L g1076 ( 
.A(n_1027),
.B(n_957),
.Y(n_1076)
);

INVx2_ASAP7_75t_SL g1077 ( 
.A(n_1009),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_988),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_1037),
.A2(n_1024),
.B1(n_999),
.B2(n_1041),
.Y(n_1079)
);

OAI21xp33_ASAP7_75t_SL g1080 ( 
.A1(n_1049),
.A2(n_967),
.B(n_855),
.Y(n_1080)
);

CKINVDCx20_ASAP7_75t_R g1081 ( 
.A(n_1033),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1035),
.Y(n_1082)
);

AOI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_1013),
.A2(n_825),
.B1(n_821),
.B2(n_870),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1036),
.Y(n_1084)
);

INVx4_ASAP7_75t_L g1085 ( 
.A(n_1019),
.Y(n_1085)
);

CKINVDCx11_ASAP7_75t_R g1086 ( 
.A(n_1033),
.Y(n_1086)
);

BUFx8_ASAP7_75t_L g1087 ( 
.A(n_990),
.Y(n_1087)
);

INVx1_ASAP7_75t_SL g1088 ( 
.A(n_998),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_1049),
.A2(n_875),
.B1(n_949),
.B2(n_858),
.Y(n_1089)
);

OAI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_1021),
.A2(n_936),
.B1(n_958),
.B2(n_952),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_1047),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1043),
.Y(n_1092)
);

BUFx12f_ASAP7_75t_L g1093 ( 
.A(n_1017),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_989),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_996),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1044),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_989),
.Y(n_1097)
);

BUFx8_ASAP7_75t_L g1098 ( 
.A(n_1017),
.Y(n_1098)
);

BUFx2_ASAP7_75t_SL g1099 ( 
.A(n_1000),
.Y(n_1099)
);

CKINVDCx11_ASAP7_75t_R g1100 ( 
.A(n_1038),
.Y(n_1100)
);

INVx6_ASAP7_75t_L g1101 ( 
.A(n_1032),
.Y(n_1101)
);

BUFx12f_ASAP7_75t_L g1102 ( 
.A(n_1032),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_SL g1103 ( 
.A1(n_1038),
.A2(n_867),
.B1(n_877),
.B2(n_891),
.Y(n_1103)
);

OR2x2_ASAP7_75t_L g1104 ( 
.A(n_1025),
.B(n_966),
.Y(n_1104)
);

CKINVDCx11_ASAP7_75t_R g1105 ( 
.A(n_1000),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_1013),
.A2(n_825),
.B1(n_821),
.B2(n_840),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_996),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1044),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_1013),
.B(n_966),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_995),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_995),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_SL g1112 ( 
.A1(n_1020),
.A2(n_867),
.B1(n_894),
.B2(n_891),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_SL g1113 ( 
.A1(n_1020),
.A2(n_867),
.B1(n_894),
.B2(n_904),
.Y(n_1113)
);

NAND2x1p5_ASAP7_75t_L g1114 ( 
.A(n_1011),
.B(n_956),
.Y(n_1114)
);

BUFx4f_ASAP7_75t_L g1115 ( 
.A(n_1048),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1044),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_1060),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1057),
.Y(n_1118)
);

INVx11_ASAP7_75t_L g1119 ( 
.A(n_1098),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_1069),
.B(n_1001),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_1090),
.B(n_986),
.Y(n_1121)
);

HB1xp67_ASAP7_75t_L g1122 ( 
.A(n_1058),
.Y(n_1122)
);

INVx4_ASAP7_75t_L g1123 ( 
.A(n_1105),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1053),
.A2(n_1048),
.B1(n_959),
.B2(n_976),
.Y(n_1124)
);

OAI21xp33_ASAP7_75t_L g1125 ( 
.A1(n_1079),
.A2(n_1062),
.B(n_1053),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1064),
.A2(n_1048),
.B1(n_994),
.B2(n_986),
.Y(n_1126)
);

OAI21xp33_ASAP7_75t_L g1127 ( 
.A1(n_1079),
.A2(n_904),
.B(n_973),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1067),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1070),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_1088),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1109),
.B(n_973),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1073),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1052),
.A2(n_1113),
.B1(n_1075),
.B2(n_1074),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_1085),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_SL g1135 ( 
.A1(n_1051),
.A2(n_1002),
.B1(n_1020),
.B2(n_1047),
.Y(n_1135)
);

OAI21xp5_ASAP7_75t_SL g1136 ( 
.A1(n_1075),
.A2(n_878),
.B(n_893),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_L g1137 ( 
.A1(n_1052),
.A2(n_994),
.B1(n_1010),
.B2(n_1005),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1076),
.B(n_1001),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_SL g1139 ( 
.A1(n_1113),
.A2(n_963),
.B(n_882),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_1085),
.B(n_1042),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1082),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1074),
.A2(n_1005),
.B1(n_1010),
.B2(n_936),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1066),
.B(n_1072),
.Y(n_1143)
);

AOI22xp33_ASAP7_75t_L g1144 ( 
.A1(n_1059),
.A2(n_1010),
.B1(n_1005),
.B2(n_919),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_1059),
.A2(n_1010),
.B1(n_1005),
.B2(n_919),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_L g1146 ( 
.A1(n_1090),
.A2(n_1005),
.B1(n_1010),
.B2(n_907),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_1084),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_1103),
.A2(n_1112),
.B1(n_1106),
.B2(n_1083),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1092),
.Y(n_1149)
);

OAI21xp33_ASAP7_75t_L g1150 ( 
.A1(n_1106),
.A2(n_873),
.B(n_871),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_L g1151 ( 
.A1(n_1112),
.A2(n_1005),
.B1(n_1010),
.B2(n_907),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_SL g1152 ( 
.A1(n_1103),
.A2(n_963),
.B(n_888),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1066),
.A2(n_1010),
.B1(n_1005),
.B2(n_899),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_SL g1154 ( 
.A1(n_1089),
.A2(n_879),
.B(n_915),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_SL g1155 ( 
.A1(n_1083),
.A2(n_1039),
.B(n_928),
.Y(n_1155)
);

AOI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_1096),
.A2(n_901),
.B1(n_899),
.B2(n_834),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1115),
.A2(n_1042),
.B1(n_968),
.B2(n_1019),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1115),
.A2(n_1019),
.B1(n_871),
.B2(n_883),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1108),
.A2(n_901),
.B1(n_899),
.B2(n_834),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1116),
.A2(n_901),
.B1(n_883),
.B2(n_873),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_1054),
.Y(n_1161)
);

AOI22xp33_ASAP7_75t_SL g1162 ( 
.A1(n_1089),
.A2(n_1019),
.B1(n_865),
.B2(n_1022),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1080),
.A2(n_840),
.B1(n_847),
.B2(n_866),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_1104),
.A2(n_847),
.B1(n_866),
.B2(n_868),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1063),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1072),
.A2(n_866),
.B1(n_868),
.B2(n_885),
.Y(n_1166)
);

OAI21xp33_ASAP7_75t_L g1167 ( 
.A1(n_1055),
.A2(n_892),
.B(n_885),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1050),
.A2(n_1022),
.B1(n_1028),
.B2(n_1015),
.Y(n_1168)
);

OAI222xp33_ASAP7_75t_L g1169 ( 
.A1(n_1081),
.A2(n_1029),
.B1(n_905),
.B2(n_892),
.C1(n_902),
.C2(n_937),
.Y(n_1169)
);

OAI21xp33_ASAP7_75t_L g1170 ( 
.A1(n_1091),
.A2(n_905),
.B(n_902),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_1071),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1099),
.A2(n_1028),
.B1(n_1015),
.B2(n_831),
.Y(n_1172)
);

AOI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1101),
.A2(n_833),
.B1(n_884),
.B2(n_880),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_SL g1174 ( 
.A1(n_1101),
.A2(n_865),
.B1(n_828),
.B2(n_833),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1093),
.A2(n_833),
.B1(n_839),
.B2(n_865),
.Y(n_1175)
);

AOI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1102),
.A2(n_833),
.B1(n_839),
.B2(n_828),
.Y(n_1176)
);

BUFx12f_ASAP7_75t_L g1177 ( 
.A(n_1086),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1101),
.A2(n_1029),
.B1(n_1006),
.B2(n_1011),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1100),
.A2(n_1098),
.B1(n_1077),
.B2(n_1065),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1068),
.B(n_889),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_SL g1181 ( 
.A1(n_1061),
.A2(n_889),
.B1(n_887),
.B2(n_581),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_SL g1182 ( 
.A1(n_1061),
.A2(n_585),
.B1(n_587),
.B2(n_591),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_1087),
.Y(n_1183)
);

BUFx12f_ASAP7_75t_L g1184 ( 
.A(n_1087),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_SL g1185 ( 
.A1(n_1114),
.A2(n_835),
.B(n_827),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1125),
.A2(n_1097),
.B1(n_1111),
.B2(n_1110),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1133),
.A2(n_1094),
.B1(n_1078),
.B2(n_1056),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1143),
.B(n_1071),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1129),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1130),
.B(n_1071),
.Y(n_1190)
);

AOI221xp5_ASAP7_75t_L g1191 ( 
.A1(n_1148),
.A2(n_628),
.B1(n_585),
.B2(n_587),
.C(n_591),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1138),
.B(n_1095),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1122),
.B(n_1095),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1127),
.A2(n_1056),
.B1(n_826),
.B2(n_1114),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1118),
.B(n_1095),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1126),
.A2(n_1046),
.B1(n_1045),
.B2(n_1030),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1124),
.A2(n_903),
.B1(n_592),
.B2(n_599),
.Y(n_1197)
);

OAI222xp33_ASAP7_75t_L g1198 ( 
.A1(n_1162),
.A2(n_970),
.B1(n_964),
.B2(n_956),
.C1(n_955),
.C2(n_917),
.Y(n_1198)
);

AOI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1170),
.A2(n_964),
.B1(n_970),
.B2(n_965),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1121),
.A2(n_628),
.B1(n_585),
.B2(n_587),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_SL g1201 ( 
.A1(n_1158),
.A2(n_1107),
.B1(n_1046),
.B2(n_1045),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1146),
.A2(n_1142),
.B1(n_1131),
.B2(n_1162),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1181),
.A2(n_1046),
.B1(n_1045),
.B2(n_1030),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1150),
.A2(n_628),
.B1(n_591),
.B2(n_592),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1144),
.A2(n_630),
.B1(n_592),
.B2(n_599),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1145),
.A2(n_630),
.B1(n_599),
.B2(n_620),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1167),
.A2(n_620),
.B1(n_622),
.B2(n_623),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1151),
.A2(n_620),
.B1(n_622),
.B2(n_623),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1122),
.B(n_1107),
.Y(n_1209)
);

AND2x2_ASAP7_75t_SL g1210 ( 
.A(n_1137),
.B(n_1011),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1181),
.A2(n_1030),
.B1(n_1018),
.B2(n_1107),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1147),
.B(n_622),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1128),
.B(n_996),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1147),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_SL g1215 ( 
.A1(n_1135),
.A2(n_1018),
.B1(n_1016),
.B2(n_1008),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_SL g1216 ( 
.A1(n_1123),
.A2(n_1018),
.B1(n_630),
.B2(n_623),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1175),
.A2(n_626),
.B1(n_823),
.B2(n_979),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1179),
.A2(n_626),
.B1(n_823),
.B2(n_1007),
.Y(n_1218)
);

OAI222xp33_ASAP7_75t_L g1219 ( 
.A1(n_1182),
.A2(n_1173),
.B1(n_1135),
.B2(n_1164),
.C1(n_1174),
.C2(n_1160),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1155),
.A2(n_1016),
.B1(n_1008),
.B2(n_1007),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1182),
.A2(n_626),
.B1(n_823),
.B2(n_1007),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1123),
.A2(n_823),
.B1(n_1008),
.B2(n_1007),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1132),
.Y(n_1223)
);

OAI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1139),
.A2(n_1016),
.B1(n_1008),
.B2(n_842),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1166),
.A2(n_1016),
.B1(n_897),
.B2(n_843),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1141),
.B(n_1149),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1152),
.A2(n_897),
.B1(n_543),
.B2(n_561),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1163),
.B(n_897),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1120),
.A2(n_897),
.B1(n_543),
.B2(n_561),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1165),
.B(n_44),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1153),
.A2(n_561),
.B1(n_543),
.B2(n_554),
.Y(n_1231)
);

AOI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1136),
.A2(n_564),
.B1(n_554),
.B2(n_527),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1180),
.B(n_45),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1172),
.A2(n_564),
.B1(n_554),
.B2(n_527),
.Y(n_1234)
);

AOI222xp33_ASAP7_75t_L g1235 ( 
.A1(n_1184),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.C1(n_48),
.C2(n_50),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1168),
.A2(n_564),
.B1(n_554),
.B2(n_527),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1140),
.B(n_47),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1174),
.A2(n_564),
.B1(n_527),
.B2(n_520),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1176),
.A2(n_520),
.B1(n_518),
.B2(n_51),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1177),
.A2(n_520),
.B1(n_518),
.B2(n_51),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1161),
.A2(n_518),
.B1(n_50),
.B2(n_53),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1140),
.B(n_48),
.Y(n_1242)
);

OAI221xp5_ASAP7_75t_L g1243 ( 
.A1(n_1185),
.A2(n_1154),
.B1(n_1156),
.B2(n_1159),
.C(n_1157),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_1178),
.B(n_55),
.Y(n_1244)
);

NAND3xp33_ASAP7_75t_L g1245 ( 
.A(n_1117),
.B(n_56),
.C(n_57),
.Y(n_1245)
);

AOI221xp5_ASAP7_75t_L g1246 ( 
.A1(n_1169),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.C(n_60),
.Y(n_1246)
);

OAI21xp33_ASAP7_75t_SL g1247 ( 
.A1(n_1134),
.A2(n_59),
.B(n_60),
.Y(n_1247)
);

AOI222xp33_ASAP7_75t_L g1248 ( 
.A1(n_1183),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.C1(n_64),
.C2(n_65),
.Y(n_1248)
);

OAI222xp33_ASAP7_75t_L g1249 ( 
.A1(n_1134),
.A2(n_61),
.B1(n_62),
.B2(n_65),
.C1(n_66),
.C2(n_67),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_SL g1250 ( 
.A1(n_1171),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1171),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1119),
.A2(n_68),
.B1(n_69),
.B2(n_79),
.Y(n_1252)
);

NAND3xp33_ASAP7_75t_L g1253 ( 
.A(n_1235),
.B(n_1171),
.C(n_82),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1226),
.B(n_1171),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_1194),
.B(n_81),
.Y(n_1255)
);

OA211x2_ASAP7_75t_L g1256 ( 
.A1(n_1191),
.A2(n_84),
.B(n_85),
.C(n_88),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1188),
.B(n_90),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1189),
.B(n_91),
.Y(n_1258)
);

NAND4xp25_ASAP7_75t_L g1259 ( 
.A(n_1248),
.B(n_92),
.C(n_94),
.D(n_99),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1189),
.B(n_100),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1223),
.B(n_102),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1226),
.B(n_103),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1192),
.B(n_104),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1195),
.B(n_105),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1246),
.A2(n_108),
.B1(n_110),
.B2(n_111),
.Y(n_1265)
);

NAND4xp25_ASAP7_75t_L g1266 ( 
.A(n_1245),
.B(n_112),
.C(n_113),
.D(n_119),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1195),
.B(n_323),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1214),
.B(n_126),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1214),
.B(n_129),
.Y(n_1269)
);

NAND3xp33_ASAP7_75t_L g1270 ( 
.A(n_1250),
.B(n_132),
.C(n_135),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1223),
.B(n_136),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1213),
.B(n_138),
.Y(n_1272)
);

NAND3xp33_ASAP7_75t_L g1273 ( 
.A(n_1241),
.B(n_141),
.C(n_142),
.Y(n_1273)
);

NAND4xp25_ASAP7_75t_L g1274 ( 
.A(n_1233),
.B(n_145),
.C(n_148),
.D(n_149),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1193),
.B(n_150),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1209),
.B(n_153),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1244),
.A2(n_1240),
.B1(n_1252),
.B2(n_1239),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1213),
.B(n_154),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1251),
.B(n_156),
.Y(n_1279)
);

OAI21xp5_ASAP7_75t_SL g1280 ( 
.A1(n_1219),
.A2(n_159),
.B(n_160),
.Y(n_1280)
);

OAI221xp5_ASAP7_75t_SL g1281 ( 
.A1(n_1247),
.A2(n_165),
.B1(n_167),
.B2(n_172),
.C(n_173),
.Y(n_1281)
);

OA21x2_ASAP7_75t_L g1282 ( 
.A1(n_1232),
.A2(n_1198),
.B(n_1227),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1190),
.B(n_178),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1187),
.B(n_181),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_SL g1285 ( 
.A1(n_1243),
.A2(n_182),
.B1(n_183),
.B2(n_188),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1244),
.B(n_195),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1230),
.B(n_1212),
.Y(n_1287)
);

OAI221xp5_ASAP7_75t_SL g1288 ( 
.A1(n_1247),
.A2(n_197),
.B1(n_200),
.B2(n_201),
.C(n_203),
.Y(n_1288)
);

NOR2xp67_ASAP7_75t_L g1289 ( 
.A(n_1237),
.B(n_204),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1251),
.B(n_205),
.Y(n_1290)
);

NAND3xp33_ASAP7_75t_L g1291 ( 
.A(n_1216),
.B(n_206),
.C(n_207),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1224),
.B(n_209),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1202),
.B(n_212),
.Y(n_1293)
);

AND2x2_ASAP7_75t_SL g1294 ( 
.A(n_1210),
.B(n_219),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1242),
.B(n_222),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1210),
.B(n_1220),
.Y(n_1296)
);

OA21x2_ASAP7_75t_L g1297 ( 
.A1(n_1238),
.A2(n_223),
.B(n_227),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1215),
.Y(n_1298)
);

NAND3xp33_ASAP7_75t_L g1299 ( 
.A(n_1186),
.B(n_228),
.C(n_231),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1197),
.A2(n_322),
.B1(n_238),
.B2(n_242),
.Y(n_1300)
);

NAND2xp33_ASAP7_75t_SL g1301 ( 
.A(n_1221),
.B(n_235),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1254),
.B(n_1201),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1296),
.B(n_1222),
.Y(n_1303)
);

AND2x4_ASAP7_75t_L g1304 ( 
.A(n_1279),
.B(n_1234),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1287),
.Y(n_1305)
);

INVxp67_ASAP7_75t_SL g1306 ( 
.A(n_1268),
.Y(n_1306)
);

AND4x1_ASAP7_75t_L g1307 ( 
.A(n_1253),
.B(n_1218),
.C(n_1200),
.D(n_1208),
.Y(n_1307)
);

NOR3xp33_ASAP7_75t_L g1308 ( 
.A(n_1280),
.B(n_1249),
.C(n_1196),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1269),
.B(n_1229),
.Y(n_1309)
);

OA211x2_ASAP7_75t_L g1310 ( 
.A1(n_1255),
.A2(n_1205),
.B(n_1206),
.C(n_1236),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1294),
.B(n_1211),
.Y(n_1311)
);

NAND3xp33_ASAP7_75t_L g1312 ( 
.A(n_1286),
.B(n_1207),
.C(n_1203),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_1298),
.B(n_1228),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1294),
.B(n_1228),
.Y(n_1314)
);

NAND4xp75_ASAP7_75t_L g1315 ( 
.A(n_1256),
.B(n_1199),
.C(n_1204),
.D(n_245),
.Y(n_1315)
);

NAND3xp33_ASAP7_75t_L g1316 ( 
.A(n_1286),
.B(n_1217),
.C(n_1231),
.Y(n_1316)
);

NAND3xp33_ASAP7_75t_L g1317 ( 
.A(n_1259),
.B(n_1199),
.C(n_1225),
.Y(n_1317)
);

NAND3xp33_ASAP7_75t_L g1318 ( 
.A(n_1285),
.B(n_243),
.C(n_244),
.Y(n_1318)
);

INVx2_ASAP7_75t_SL g1319 ( 
.A(n_1261),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1272),
.B(n_249),
.Y(n_1320)
);

NAND4xp75_ASAP7_75t_L g1321 ( 
.A(n_1255),
.B(n_251),
.C(n_252),
.D(n_253),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1262),
.B(n_254),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1261),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1279),
.B(n_255),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1258),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1278),
.B(n_256),
.Y(n_1326)
);

NAND3xp33_ASAP7_75t_L g1327 ( 
.A(n_1281),
.B(n_257),
.C(n_258),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1272),
.B(n_263),
.Y(n_1328)
);

NOR3xp33_ASAP7_75t_SL g1329 ( 
.A(n_1274),
.B(n_1266),
.C(n_1288),
.Y(n_1329)
);

NOR3xp33_ASAP7_75t_L g1330 ( 
.A(n_1273),
.B(n_271),
.C(n_275),
.Y(n_1330)
);

INVxp33_ASAP7_75t_SL g1331 ( 
.A(n_1311),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1319),
.B(n_1305),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1323),
.Y(n_1333)
);

NAND3xp33_ASAP7_75t_L g1334 ( 
.A(n_1329),
.B(n_1265),
.C(n_1292),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1325),
.Y(n_1335)
);

NOR3xp33_ASAP7_75t_L g1336 ( 
.A(n_1327),
.B(n_1270),
.C(n_1293),
.Y(n_1336)
);

NAND4xp75_ASAP7_75t_SL g1337 ( 
.A(n_1313),
.B(n_1282),
.C(n_1297),
.D(n_1292),
.Y(n_1337)
);

XOR2xp5_ASAP7_75t_L g1338 ( 
.A(n_1322),
.B(n_1264),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1306),
.B(n_1283),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1325),
.Y(n_1340)
);

INVx1_ASAP7_75t_SL g1341 ( 
.A(n_1302),
.Y(n_1341)
);

INVx4_ASAP7_75t_L g1342 ( 
.A(n_1324),
.Y(n_1342)
);

NOR3xp33_ASAP7_75t_L g1343 ( 
.A(n_1312),
.B(n_1289),
.C(n_1276),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1319),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1302),
.B(n_1267),
.Y(n_1345)
);

XOR2x2_ASAP7_75t_L g1346 ( 
.A(n_1308),
.B(n_1277),
.Y(n_1346)
);

NAND4xp75_ASAP7_75t_L g1347 ( 
.A(n_1329),
.B(n_1282),
.C(n_1295),
.D(n_1297),
.Y(n_1347)
);

INVx5_ASAP7_75t_L g1348 ( 
.A(n_1324),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_1320),
.Y(n_1349)
);

INVx4_ASAP7_75t_L g1350 ( 
.A(n_1324),
.Y(n_1350)
);

INVx2_ASAP7_75t_SL g1351 ( 
.A(n_1303),
.Y(n_1351)
);

INVx2_ASAP7_75t_SL g1352 ( 
.A(n_1333),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1335),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1340),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1333),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1342),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_SL g1357 ( 
.A(n_1331),
.B(n_1321),
.Y(n_1357)
);

XNOR2x1_ASAP7_75t_L g1358 ( 
.A(n_1346),
.B(n_1310),
.Y(n_1358)
);

XOR2xp5_ASAP7_75t_L g1359 ( 
.A(n_1346),
.B(n_1320),
.Y(n_1359)
);

XNOR2xp5_ASAP7_75t_L g1360 ( 
.A(n_1338),
.B(n_1314),
.Y(n_1360)
);

XNOR2x1_ASAP7_75t_L g1361 ( 
.A(n_1334),
.B(n_1315),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1351),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1332),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1351),
.Y(n_1364)
);

XNOR2xp5_ASAP7_75t_L g1365 ( 
.A(n_1331),
.B(n_1277),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1356),
.Y(n_1366)
);

CKINVDCx16_ASAP7_75t_R g1367 ( 
.A(n_1357),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1353),
.Y(n_1368)
);

INVx1_ASAP7_75t_SL g1369 ( 
.A(n_1358),
.Y(n_1369)
);

XNOR2x1_ASAP7_75t_L g1370 ( 
.A(n_1358),
.B(n_1341),
.Y(n_1370)
);

OA22x2_ASAP7_75t_L g1371 ( 
.A1(n_1365),
.A2(n_1342),
.B1(n_1350),
.B2(n_1349),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1356),
.B(n_1364),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1356),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1353),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1352),
.Y(n_1375)
);

OA22x2_ASAP7_75t_L g1376 ( 
.A1(n_1365),
.A2(n_1350),
.B1(n_1342),
.B2(n_1345),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1361),
.A2(n_1336),
.B1(n_1343),
.B2(n_1330),
.Y(n_1377)
);

XNOR2x1_ASAP7_75t_L g1378 ( 
.A(n_1359),
.B(n_1347),
.Y(n_1378)
);

OR2x6_ASAP7_75t_L g1379 ( 
.A(n_1364),
.B(n_1350),
.Y(n_1379)
);

OAI22xp33_ASAP7_75t_SL g1380 ( 
.A1(n_1359),
.A2(n_1348),
.B1(n_1339),
.B2(n_1344),
.Y(n_1380)
);

INVx1_ASAP7_75t_SL g1381 ( 
.A(n_1362),
.Y(n_1381)
);

OA22x2_ASAP7_75t_L g1382 ( 
.A1(n_1360),
.A2(n_1304),
.B1(n_1328),
.B2(n_1290),
.Y(n_1382)
);

XOR2x2_ASAP7_75t_L g1383 ( 
.A(n_1360),
.B(n_1337),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1378),
.A2(n_1361),
.B1(n_1348),
.B2(n_1313),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1368),
.Y(n_1385)
);

AOI322xp5_ASAP7_75t_L g1386 ( 
.A1(n_1369),
.A2(n_1377),
.A3(n_1367),
.B1(n_1381),
.B2(n_1383),
.C1(n_1370),
.C2(n_1380),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1381),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1372),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1368),
.Y(n_1389)
);

INVx2_ASAP7_75t_SL g1390 ( 
.A(n_1372),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1374),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1374),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1376),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1379),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_1394),
.Y(n_1395)
);

OAI322xp33_ASAP7_75t_L g1396 ( 
.A1(n_1384),
.A2(n_1367),
.A3(n_1371),
.B1(n_1382),
.B2(n_1373),
.C1(n_1366),
.C2(n_1380),
.Y(n_1396)
);

AOI22x1_ASAP7_75t_L g1397 ( 
.A1(n_1393),
.A2(n_1375),
.B1(n_1354),
.B2(n_1304),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1387),
.A2(n_1394),
.B1(n_1390),
.B2(n_1388),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1387),
.Y(n_1399)
);

AOI221xp5_ASAP7_75t_L g1400 ( 
.A1(n_1386),
.A2(n_1339),
.B1(n_1317),
.B2(n_1265),
.C(n_1355),
.Y(n_1400)
);

OAI322xp33_ASAP7_75t_L g1401 ( 
.A1(n_1390),
.A2(n_1352),
.A3(n_1363),
.B1(n_1309),
.B2(n_1326),
.C1(n_1316),
.C2(n_1284),
.Y(n_1401)
);

OA22x2_ASAP7_75t_SL g1402 ( 
.A1(n_1388),
.A2(n_1379),
.B1(n_1348),
.B2(n_1307),
.Y(n_1402)
);

INVxp67_ASAP7_75t_SL g1403 ( 
.A(n_1394),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1385),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1399),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1395),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1400),
.A2(n_1318),
.B(n_1326),
.C(n_1348),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1403),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1404),
.Y(n_1409)
);

O2A1O1Ixp5_ASAP7_75t_SL g1410 ( 
.A1(n_1395),
.A2(n_1392),
.B(n_1391),
.C(n_1389),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1398),
.Y(n_1411)
);

NOR4xp25_ASAP7_75t_L g1412 ( 
.A(n_1411),
.B(n_1396),
.C(n_1401),
.D(n_1402),
.Y(n_1412)
);

OAI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1408),
.A2(n_1397),
.B1(n_1299),
.B2(n_1291),
.Y(n_1413)
);

INVxp67_ASAP7_75t_SL g1414 ( 
.A(n_1406),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1405),
.Y(n_1415)
);

AO22x2_ASAP7_75t_L g1416 ( 
.A1(n_1409),
.A2(n_1304),
.B1(n_1271),
.B2(n_1275),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1407),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1407),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1410),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1408),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1414),
.Y(n_1421)
);

INVxp67_ASAP7_75t_L g1422 ( 
.A(n_1417),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1420),
.Y(n_1423)
);

AOI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1418),
.A2(n_1301),
.B1(n_1257),
.B2(n_1263),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1412),
.B(n_1260),
.Y(n_1425)
);

AOI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1419),
.A2(n_1301),
.B1(n_1282),
.B2(n_1297),
.Y(n_1426)
);

AOI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1413),
.A2(n_1300),
.B1(n_286),
.B2(n_287),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1421),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1423),
.Y(n_1429)
);

AOI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1425),
.A2(n_1416),
.B1(n_1415),
.B2(n_290),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1422),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1428),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1431),
.Y(n_1433)
);

INVxp67_ASAP7_75t_L g1434 ( 
.A(n_1429),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1430),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1428),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1428),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1432),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1435),
.A2(n_1427),
.B1(n_1426),
.B2(n_1416),
.Y(n_1439)
);

OAI22x1_ASAP7_75t_L g1440 ( 
.A1(n_1436),
.A2(n_1424),
.B1(n_288),
.B2(n_291),
.Y(n_1440)
);

OAI22x1_ASAP7_75t_L g1441 ( 
.A1(n_1437),
.A2(n_285),
.B1(n_292),
.B2(n_294),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1438),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1440),
.Y(n_1443)
);

INVxp67_ASAP7_75t_L g1444 ( 
.A(n_1441),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1439),
.Y(n_1445)
);

OAI22xp33_ASAP7_75t_SL g1446 ( 
.A1(n_1445),
.A2(n_1432),
.B1(n_1433),
.B2(n_1434),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1444),
.A2(n_295),
.B1(n_298),
.B2(n_299),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1443),
.A2(n_300),
.B1(n_302),
.B2(n_303),
.Y(n_1448)
);

INVxp67_ASAP7_75t_SL g1449 ( 
.A(n_1446),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1447),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1449),
.A2(n_1448),
.B1(n_1442),
.B2(n_307),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1451),
.Y(n_1452)
);

AOI221xp5_ASAP7_75t_L g1453 ( 
.A1(n_1452),
.A2(n_1450),
.B1(n_305),
.B2(n_310),
.C(n_311),
.Y(n_1453)
);

AOI211xp5_ASAP7_75t_L g1454 ( 
.A1(n_1453),
.A2(n_304),
.B(n_314),
.C(n_315),
.Y(n_1454)
);


endmodule