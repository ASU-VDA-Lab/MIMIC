module fake_jpeg_13403_n_340 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_0),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_1),
.B(n_2),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_17),
.B(n_23),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_38),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

NAND2xp33_ASAP7_75t_SL g43 ( 
.A(n_17),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_46),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_32),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_18),
.B(n_1),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_18),
.B(n_8),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_48),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_28),
.C(n_31),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_35),
.Y(n_75)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_53),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_29),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_63),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_31),
.B1(n_28),
.B2(n_16),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_59),
.A2(n_70),
.B1(n_28),
.B2(n_32),
.Y(n_87)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_37),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_60),
.Y(n_102)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_31),
.B1(n_28),
.B2(n_16),
.Y(n_70)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_51),
.A2(n_47),
.B1(n_22),
.B2(n_25),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_74),
.A2(n_93),
.B1(n_95),
.B2(n_100),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_41),
.C(n_64),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_35),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_76),
.B(n_77),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_35),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_36),
.B1(n_38),
.B2(n_40),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_81),
.A2(n_87),
.B1(n_101),
.B2(n_41),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_58),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_88),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_35),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_84),
.B(n_86),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_55),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_60),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_52),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_99),
.Y(n_115)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_51),
.A2(n_22),
.B1(n_25),
.B2(n_24),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_68),
.A2(n_24),
.B1(n_46),
.B2(n_27),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_38),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_54),
.A2(n_20),
.B1(n_40),
.B2(n_39),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_71),
.B1(n_54),
.B2(n_42),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_48),
.A2(n_35),
.B(n_30),
.C(n_27),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_69),
.A2(n_29),
.B1(n_20),
.B2(n_41),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_65),
.A2(n_41),
.B1(n_42),
.B2(n_39),
.Y(n_101)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_2),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_106),
.B(n_2),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_84),
.A2(n_103),
.B1(n_81),
.B2(n_76),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_108),
.A2(n_119),
.B1(n_128),
.B2(n_129),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_109),
.B(n_110),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_112),
.B(n_124),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_39),
.B1(n_42),
.B2(n_66),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_113),
.A2(n_114),
.B1(n_104),
.B2(n_79),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_82),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_118),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_103),
.A2(n_42),
.B1(n_71),
.B2(n_66),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_102),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_122),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_77),
.A2(n_30),
.B(n_57),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_78),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_80),
.B(n_15),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_125),
.B(n_126),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_15),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_87),
.A2(n_75),
.B1(n_99),
.B2(n_73),
.Y(n_128)
);

INVxp33_ASAP7_75t_SL g130 ( 
.A(n_88),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_130),
.B(n_90),
.Y(n_145)
);

INVxp33_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_131),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_19),
.B1(n_52),
.B2(n_57),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_135),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_91),
.A2(n_19),
.B1(n_30),
.B2(n_34),
.Y(n_135)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_143),
.A2(n_160),
.B1(n_165),
.B2(n_122),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_126),
.B(n_90),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_144),
.B(n_153),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_163),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_111),
.Y(n_146)
);

INVx13_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_111),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_127),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_79),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_155),
.Y(n_170)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_150),
.A2(n_130),
.B(n_121),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_112),
.B(n_85),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_151),
.B(n_156),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_85),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_152),
.A2(n_94),
.B(n_26),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_107),
.B(n_90),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_89),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_117),
.B(n_97),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_108),
.B(n_97),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_162),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_114),
.A2(n_83),
.B1(n_78),
.B2(n_94),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_117),
.B(n_83),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_SL g163 ( 
.A1(n_115),
.A2(n_133),
.B(n_123),
.Y(n_163)
);

OR2x2_ASAP7_75t_SL g164 ( 
.A(n_115),
.B(n_2),
.Y(n_164)
);

NOR3xp33_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_125),
.C(n_119),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_114),
.A2(n_94),
.B1(n_19),
.B2(n_34),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_108),
.B(n_3),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_3),
.Y(n_198)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_118),
.Y(n_168)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_168),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_169),
.A2(n_201),
.B(n_5),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_121),
.B1(n_128),
.B2(n_133),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_171),
.A2(n_174),
.B1(n_182),
.B2(n_34),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_145),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_172),
.B(n_199),
.Y(n_218)
);

AO22x1_ASAP7_75t_SL g176 ( 
.A1(n_163),
.A2(n_140),
.B1(n_152),
.B2(n_158),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_198),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_178),
.B(n_180),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_141),
.A2(n_113),
.B1(n_132),
.B2(n_129),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_183),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_152),
.A2(n_119),
.B1(n_135),
.B2(n_120),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_185),
.A2(n_165),
.B1(n_160),
.B2(n_141),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_186),
.A2(n_159),
.B(n_144),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_136),
.B(n_12),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_187),
.B(n_202),
.Y(n_228)
);

BUFx24_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_138),
.Y(n_192)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_138),
.Y(n_193)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_139),
.B(n_151),
.C(n_155),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_196),
.C(n_200),
.Y(n_204)
);

OA22x2_ASAP7_75t_L g195 ( 
.A1(n_146),
.A2(n_19),
.B1(n_26),
.B2(n_21),
.Y(n_195)
);

OA22x2_ASAP7_75t_L g203 ( 
.A1(n_195),
.A2(n_168),
.B1(n_150),
.B2(n_147),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_139),
.B(n_34),
.C(n_26),
.Y(n_196)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_154),
.Y(n_197)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_197),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_157),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_156),
.B(n_34),
.C(n_10),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_150),
.A2(n_3),
.B(n_4),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_157),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_223),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_205),
.A2(n_219),
.B1(n_229),
.B2(n_183),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_162),
.C(n_167),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_209),
.C(n_212),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_169),
.A2(n_143),
.B1(n_148),
.B2(n_168),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_208),
.A2(n_222),
.B1(n_197),
.B2(n_186),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_170),
.B(n_149),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_189),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_210),
.B(n_206),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_170),
.B(n_142),
.C(n_137),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_137),
.C(n_154),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_213),
.B(n_200),
.C(n_192),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_214),
.A2(n_221),
.B(n_224),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_185),
.A2(n_164),
.B1(n_136),
.B2(n_161),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_164),
.Y(n_220)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

OA22x2_ASAP7_75t_L g223 ( 
.A1(n_176),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_179),
.A2(n_10),
.B(n_14),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_179),
.A2(n_5),
.B(n_6),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_225),
.A2(n_201),
.B(n_221),
.Y(n_253)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_173),
.Y(n_227)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_227),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_174),
.A2(n_7),
.B1(n_9),
.B2(n_12),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_177),
.B(n_172),
.Y(n_231)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_230),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_233),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_179),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_234),
.B(n_241),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_237),
.A2(n_238),
.B1(n_252),
.B2(n_256),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_208),
.A2(n_177),
.B1(n_176),
.B2(n_184),
.Y(n_238)
);

A2O1A1O1Ixp25_ASAP7_75t_L g239 ( 
.A1(n_217),
.A2(n_231),
.B(n_218),
.C(n_220),
.D(n_212),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_239),
.A2(n_253),
.B(n_219),
.Y(n_262)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_227),
.Y(n_240)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_240),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_196),
.Y(n_241)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_242),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_204),
.B(n_184),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_245),
.C(n_254),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_209),
.B(n_190),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_211),
.Y(n_248)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_248),
.Y(n_268)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_215),
.Y(n_249)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_249),
.Y(n_275)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_206),
.Y(n_250)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_250),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_190),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_255),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_216),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_175),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_228),
.B(n_188),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_224),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_234),
.B(n_213),
.Y(n_260)
);

XNOR2x1_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_261),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_244),
.B(n_217),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_266),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_203),
.C(n_214),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_265),
.C(n_270),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_245),
.C(n_254),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_236),
.B(n_203),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_203),
.C(n_226),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_274),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_232),
.A2(n_225),
.B(n_226),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_243),
.B(n_205),
.C(n_175),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_251),
.C(n_255),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_223),
.Y(n_278)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_278),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_250),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_281),
.B(n_282),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_271),
.A2(n_238),
.B1(n_247),
.B2(n_237),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_232),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_288),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_286),
.B(n_290),
.Y(n_297)
);

INVxp33_ASAP7_75t_SL g287 ( 
.A(n_270),
.Y(n_287)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_287),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_246),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_268),
.Y(n_289)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_272),
.B(n_239),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_275),
.Y(n_291)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_291),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_258),
.A2(n_235),
.B1(n_248),
.B2(n_193),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_269),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_265),
.B(n_246),
.C(n_253),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_260),
.C(n_259),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_293),
.A2(n_262),
.B(n_279),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_296),
.A2(n_302),
.B(n_191),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_285),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_259),
.C(n_266),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_305),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_280),
.A2(n_264),
.B(n_294),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_283),
.B(n_287),
.C(n_288),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_280),
.B(n_277),
.C(n_271),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_307),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_284),
.B(n_261),
.C(n_274),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_276),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_286),
.C(n_284),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_310),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_299),
.A2(n_269),
.B(n_278),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_311),
.A2(n_314),
.B(n_316),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_263),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_295),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_297),
.A2(n_191),
.B(n_173),
.Y(n_317)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_317),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_195),
.C(n_198),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_300),
.C(n_308),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_306),
.A2(n_195),
.B(n_7),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_319),
.B(n_195),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_13),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_313),
.Y(n_323)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_323),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_324),
.A2(n_318),
.B1(n_303),
.B2(n_304),
.Y(n_331)
);

INVx6_ASAP7_75t_L g326 ( 
.A(n_310),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_327),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_321),
.A2(n_311),
.B(n_315),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_328),
.A2(n_329),
.B(n_331),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_309),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_333),
.B(n_320),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_335),
.B(n_336),
.Y(n_337)
);

AOI321xp33_ASAP7_75t_L g336 ( 
.A1(n_330),
.A2(n_322),
.A3(n_324),
.B1(n_326),
.B2(n_15),
.C(n_13),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_334),
.B1(n_332),
.B2(n_328),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_14),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_6),
.Y(n_340)
);


endmodule