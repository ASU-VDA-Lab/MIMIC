module real_jpeg_8499_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_164;
wire n_48;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_0),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_43),
.Y(n_104)
);

BUFx24_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_2),
.Y(n_101)
);

AOI21xp33_ASAP7_75t_L g102 ( 
.A1(n_2),
.A2(n_57),
.B(n_61),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_2),
.A2(n_55),
.B1(n_64),
.B2(n_101),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_2),
.B(n_121),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_2),
.A2(n_41),
.B(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_2),
.B(n_41),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_2),
.A2(n_30),
.B1(n_105),
.B2(n_172),
.Y(n_174)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_SL g72 ( 
.A(n_7),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_8),
.A2(n_35),
.B1(n_41),
.B2(n_44),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_8),
.A2(n_35),
.B1(n_60),
.B2(n_61),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_10),
.A2(n_55),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_10),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_10),
.A2(n_60),
.B1(n_61),
.B2(n_65),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_65),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_10),
.A2(n_41),
.B1(n_44),
.B2(n_65),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_11),
.A2(n_55),
.B1(n_64),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_11),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_11),
.A2(n_60),
.B1(n_61),
.B2(n_97),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_11),
.A2(n_41),
.B1(n_44),
.B2(n_97),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_97),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_12),
.A2(n_29),
.B1(n_41),
.B2(n_44),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_13),
.A2(n_55),
.B1(n_64),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_13),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_13),
.A2(n_60),
.B1(n_61),
.B2(n_67),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_67),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_13),
.A2(n_41),
.B1(n_44),
.B2(n_67),
.Y(n_193)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_15),
.A2(n_60),
.B1(n_61),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_15),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_76),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_15),
.A2(n_41),
.B1(n_44),
.B2(n_76),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_127),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_125),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_107),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_20),
.B(n_107),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_87),
.B1(n_88),
.B2(n_106),
.Y(n_20)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_21),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_80),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_51),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_24),
.B(n_36),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_30),
.B(n_33),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_25),
.A2(n_30),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_26),
.B(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_26),
.A2(n_27),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_26),
.B(n_39),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_26),
.B(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_27),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_163)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_30),
.A2(n_105),
.B1(n_154),
.B2(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_30),
.A2(n_83),
.B(n_156),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_30),
.A2(n_33),
.B(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_31),
.B(n_34),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_31),
.A2(n_32),
.B1(n_153),
.B2(n_155),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_32),
.B(n_84),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_32),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_40),
.B(n_45),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_38),
.B(n_41),
.C(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_37),
.A2(n_40),
.B1(n_49),
.B2(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_37),
.B(n_47),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_37),
.A2(n_49),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_37),
.B(n_101),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_37),
.A2(n_49),
.B1(n_162),
.B2(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_37),
.A2(n_49),
.B1(n_185),
.B2(n_193),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_37),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_38),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_41),
.Y(n_50)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_41),
.A2(n_44),
.B1(n_71),
.B2(n_72),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_41),
.B(n_71),
.Y(n_200)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_44),
.A2(n_73),
.B1(n_195),
.B2(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_48),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_48),
.A2(n_123),
.B(n_124),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_49),
.A2(n_193),
.B(n_217),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_50),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_68),
.B2(n_69),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_59),
.B1(n_63),
.B2(n_66),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_54),
.A2(n_59),
.B1(n_63),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_54),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B(n_58),
.C(n_59),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_56),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_55),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_55),
.A2(n_56),
.B(n_101),
.C(n_102),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_59),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

O2A1O1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_71),
.B(n_73),
.C(n_74),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_71),
.Y(n_73)
);

HAxp5_ASAP7_75t_SL g195 ( 
.A(n_61),
.B(n_101),
.CON(n_195),
.SN(n_195)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_75),
.B(n_77),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_70),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_70),
.A2(n_74),
.B1(n_140),
.B2(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_75),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_79),
.A2(n_91),
.B1(n_92),
.B2(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_79),
.A2(n_91),
.B1(n_116),
.B2(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_79),
.B(n_101),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_82),
.A2(n_104),
.B(n_105),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_84),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_94),
.C(n_98),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_90),
.B1(n_94),
.B2(n_95),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B(n_93),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_99),
.A2(n_100),
.B1(n_103),
.B2(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_101),
.B(n_105),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_103),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.C(n_112),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.C(n_122),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_115),
.B1(n_122),
.B2(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_122),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_123),
.B(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_146),
.B(n_228),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_144),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_129),
.B(n_144),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.C(n_135),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_130),
.B(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_133),
.A2(n_135),
.B1(n_136),
.B2(n_226),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_133),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_141),
.C(n_142),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_137),
.A2(n_138),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_141),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_222),
.B(n_227),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_205),
.B(n_221),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_188),
.B(n_204),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_179),
.B(n_187),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_168),
.B(n_178),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_157),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_152),
.B(n_157),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_163),
.B2(n_167),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_158),
.B(n_167),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_161),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_163),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_173),
.B(n_177),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_170),
.B(n_171),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_180),
.B(n_181),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_182),
.B(n_189),
.Y(n_204)
);

FAx1_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_184),
.CI(n_186),
.CON(n_182),
.SN(n_182)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_198),
.B2(n_203),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_194),
.B1(n_196),
.B2(n_197),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_192),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_194),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_197),
.C(n_203),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_198),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_201),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_206),
.B(n_207),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_213),
.B2(n_214),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_216),
.C(n_219),
.Y(n_223)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_219),
.B2(n_220),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_215),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_216),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_223),
.B(n_224),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);


endmodule