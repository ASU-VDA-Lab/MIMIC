module fake_netlist_5_1790_n_1537 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_1537);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1537;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_150;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_297;
wire n_156;
wire n_1078;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_604;
wire n_433;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_689;
wire n_738;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_152;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_146;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_833;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1419;
wire n_338;
wire n_149;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_151;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_148;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_147;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_145;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1220;
wire n_229;
wire n_437;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_246;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_135),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_95),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_61),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_130),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_75),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_18),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_55),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g154 ( 
.A(n_73),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_71),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_58),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_9),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_125),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_12),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_111),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_30),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_137),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_19),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_15),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_119),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_46),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_108),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_90),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_32),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_144),
.Y(n_171)
);

BUFx10_ASAP7_75t_L g172 ( 
.A(n_48),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_118),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_129),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_38),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_29),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_142),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_21),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_83),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_59),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_15),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_88),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_68),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_103),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_143),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_34),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_63),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_106),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_99),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_23),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_114),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_39),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_123),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_33),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_14),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_80),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_43),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_128),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_53),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_69),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_47),
.Y(n_201)
);

BUFx10_ASAP7_75t_L g202 ( 
.A(n_18),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_81),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_124),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_39),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_77),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_36),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_91),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_23),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_74),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_127),
.Y(n_211)
);

BUFx8_ASAP7_75t_SL g212 ( 
.A(n_43),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_0),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_27),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_35),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_93),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_107),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_138),
.Y(n_218)
);

BUFx10_ASAP7_75t_L g219 ( 
.A(n_101),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_29),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_60),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_44),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_76),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_64),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_96),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_34),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_14),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_9),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_8),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_37),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_121),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_100),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_11),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_37),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_52),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_8),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_44),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_19),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_120),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_94),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_24),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_70),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_36),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_66),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_25),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_31),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_116),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_78),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_102),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_45),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_6),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_46),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_140),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_41),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_5),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_50),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_72),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_86),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_30),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_17),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_21),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_47),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_132),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_131),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_5),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_26),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_41),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_25),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_139),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_133),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_85),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_105),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_28),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_42),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_56),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_0),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_49),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_104),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_27),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_10),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_79),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_12),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_4),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_10),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_82),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_89),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_87),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_22),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_166),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_176),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g291 ( 
.A(n_193),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_246),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_176),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_176),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_154),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_212),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_189),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_176),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_176),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_207),
.Y(n_300)
);

INVxp67_ASAP7_75t_SL g301 ( 
.A(n_149),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_184),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_207),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_230),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_196),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_230),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_185),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_198),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_261),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_199),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_245),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_261),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_192),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_160),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_276),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_200),
.Y(n_316)
);

INVxp33_ASAP7_75t_L g317 ( 
.A(n_152),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_189),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_203),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_160),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_258),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_219),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_204),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_276),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_288),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_206),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_162),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_208),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_219),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_172),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_154),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_172),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_157),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_190),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_217),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_195),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_218),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_209),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_213),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_172),
.Y(n_340)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_202),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_214),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_221),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_229),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_234),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_202),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_162),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_202),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_223),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_224),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_237),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_226),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_225),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_219),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_232),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_239),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_318),
.B(n_215),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_290),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_290),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_293),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_295),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_293),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_297),
.B(n_215),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_311),
.A2(n_228),
.B1(n_233),
.B2(n_241),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_297),
.B(n_258),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_294),
.Y(n_366)
);

NOR2xp67_ASAP7_75t_L g367 ( 
.A(n_307),
.B(n_235),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_294),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_298),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_289),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_292),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_298),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_299),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_299),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_307),
.Y(n_375)
);

AND2x6_ASAP7_75t_L g376 ( 
.A(n_295),
.B(n_185),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_307),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_307),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_295),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_314),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_325),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_302),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_325),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_331),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_331),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_308),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_330),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_310),
.B(n_235),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_297),
.B(n_231),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_352),
.B(n_280),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_321),
.B(n_275),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_331),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_333),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_300),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_320),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_316),
.Y(n_396)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_319),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_328),
.B(n_275),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_333),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_335),
.B(n_187),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_292),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_321),
.B(n_231),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_334),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_291),
.A2(n_256),
.B1(n_181),
.B2(n_164),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_334),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_336),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_350),
.B(n_177),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_336),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_300),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_353),
.B(n_356),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_305),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_323),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_322),
.A2(n_178),
.B1(n_170),
.B2(n_167),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_321),
.B(n_187),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_322),
.A2(n_170),
.B1(n_167),
.B2(n_165),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_347),
.B(n_164),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_303),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_338),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_303),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_371),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_358),
.Y(n_421)
);

OR2x2_ASAP7_75t_L g422 ( 
.A(n_364),
.B(n_327),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_379),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_359),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_359),
.Y(n_425)
);

OR2x6_ASAP7_75t_L g426 ( 
.A(n_397),
.B(n_191),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_358),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_358),
.Y(n_428)
);

NAND3xp33_ASAP7_75t_L g429 ( 
.A(n_414),
.B(n_313),
.C(n_191),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_379),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_388),
.B(n_301),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_369),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_360),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_365),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_369),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_365),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_407),
.B(n_249),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_372),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_360),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_360),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_373),
.Y(n_441)
);

NAND3xp33_ASAP7_75t_L g442 ( 
.A(n_357),
.B(n_339),
.C(n_338),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_397),
.B(n_329),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_379),
.Y(n_444)
);

AOI22xp33_ASAP7_75t_L g445 ( 
.A1(n_357),
.A2(n_327),
.B1(n_259),
.B2(n_283),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_379),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_398),
.B(n_326),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_376),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_373),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_376),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_397),
.B(n_329),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_372),
.Y(n_452)
);

INVx6_ASAP7_75t_L g453 ( 
.A(n_379),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_374),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_374),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_400),
.B(n_281),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_397),
.B(n_354),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_379),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_385),
.Y(n_459)
);

AND2x6_ASAP7_75t_L g460 ( 
.A(n_391),
.B(n_145),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_390),
.B(n_296),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_411),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_373),
.Y(n_463)
);

INVx2_ASAP7_75t_SL g464 ( 
.A(n_389),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_361),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_390),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_391),
.B(n_242),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_363),
.B(n_315),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_376),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_384),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_389),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_384),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_361),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_384),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_385),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_392),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_361),
.Y(n_477)
);

OAI22xp33_ASAP7_75t_L g478 ( 
.A1(n_404),
.A2(n_354),
.B1(n_175),
.B2(n_252),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_361),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_392),
.Y(n_480)
);

INVx5_ASAP7_75t_L g481 ( 
.A(n_376),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_392),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_409),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_385),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_391),
.B(n_247),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_409),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_410),
.B(n_337),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_409),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_375),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_402),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_377),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_409),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g493 ( 
.A(n_402),
.Y(n_493)
);

NAND3xp33_ASAP7_75t_L g494 ( 
.A(n_363),
.B(n_342),
.C(n_339),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_382),
.B(n_355),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_404),
.A2(n_282),
.B1(n_260),
.B2(n_262),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_386),
.B(n_343),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_377),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_370),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_409),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_409),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_417),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_377),
.Y(n_503)
);

BUFx10_ASAP7_75t_L g504 ( 
.A(n_396),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_417),
.Y(n_505)
);

BUFx8_ASAP7_75t_SL g506 ( 
.A(n_412),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_375),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_391),
.B(n_248),
.Y(n_508)
);

INVx5_ASAP7_75t_L g509 ( 
.A(n_376),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_380),
.A2(n_349),
.B1(n_341),
.B2(n_243),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_387),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_417),
.Y(n_512)
);

OAI21xp33_ASAP7_75t_SL g513 ( 
.A1(n_381),
.A2(n_324),
.B(n_315),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_381),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_401),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_383),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_417),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_413),
.A2(n_415),
.B1(n_416),
.B2(n_364),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_383),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_367),
.B(n_253),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_393),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_367),
.B(n_146),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_395),
.B(n_332),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_417),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_393),
.Y(n_525)
);

INVx6_ASAP7_75t_L g526 ( 
.A(n_377),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_362),
.B(n_153),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_376),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_417),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_399),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_419),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_419),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_399),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_403),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_377),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_387),
.B(n_340),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_419),
.Y(n_537)
);

BUFx4f_ASAP7_75t_L g538 ( 
.A(n_376),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_419),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_419),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_376),
.A2(n_265),
.B1(n_250),
.B2(n_251),
.Y(n_541)
);

BUFx6f_ASAP7_75t_SL g542 ( 
.A(n_403),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_405),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_377),
.Y(n_544)
);

AND3x2_ASAP7_75t_L g545 ( 
.A(n_405),
.B(n_348),
.C(n_346),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_362),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_413),
.B(n_317),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_415),
.B(n_324),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_419),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_406),
.Y(n_550)
);

OAI22xp33_ASAP7_75t_L g551 ( 
.A1(n_408),
.A2(n_186),
.B1(n_194),
.B2(n_197),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_408),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_418),
.B(n_304),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_416),
.B(n_231),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_362),
.Y(n_555)
);

AND3x2_ASAP7_75t_L g556 ( 
.A(n_418),
.B(n_158),
.C(n_168),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_378),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_378),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_362),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_378),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_394),
.B(n_147),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_434),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_464),
.B(n_154),
.Y(n_563)
);

NOR3xp33_ASAP7_75t_L g564 ( 
.A(n_554),
.B(n_342),
.C(n_351),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_437),
.B(n_431),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_468),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_434),
.B(n_362),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_434),
.B(n_436),
.Y(n_568)
);

O2A1O1Ixp33_ASAP7_75t_L g569 ( 
.A1(n_513),
.A2(n_255),
.B(n_266),
.C(n_268),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_436),
.B(n_362),
.Y(n_570)
);

O2A1O1Ixp5_ASAP7_75t_L g571 ( 
.A1(n_514),
.A2(n_272),
.B(n_179),
.C(n_182),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_436),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_448),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_464),
.B(n_366),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_471),
.B(n_366),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_471),
.B(n_366),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_SL g577 ( 
.A(n_504),
.B(n_240),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_490),
.B(n_366),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_490),
.B(n_366),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_489),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_448),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_456),
.B(n_148),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_489),
.Y(n_583)
);

INVxp67_ASAP7_75t_SL g584 ( 
.A(n_498),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_514),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_493),
.B(n_366),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_447),
.B(n_148),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_493),
.B(n_154),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_507),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_536),
.B(n_150),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_516),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_538),
.B(n_154),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_424),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_448),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_538),
.B(n_154),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_519),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_450),
.B(n_469),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_460),
.A2(n_211),
.B1(n_264),
.B2(n_183),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_519),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_521),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_521),
.B(n_368),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_450),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_525),
.B(n_368),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_511),
.B(n_150),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_511),
.B(n_151),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_424),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_525),
.Y(n_607)
);

INVxp33_ASAP7_75t_L g608 ( 
.A(n_548),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_468),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_530),
.B(n_533),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_530),
.B(n_368),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_533),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_534),
.B(n_543),
.Y(n_613)
);

O2A1O1Ixp33_ASAP7_75t_L g614 ( 
.A1(n_513),
.A2(n_284),
.B(n_351),
.C(n_345),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_538),
.B(n_154),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_523),
.B(n_151),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_534),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_543),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_467),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_547),
.B(n_344),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_450),
.B(n_154),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_425),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_425),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_469),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_469),
.B(n_188),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_485),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_550),
.B(n_368),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_550),
.B(n_368),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_510),
.B(n_487),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_432),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_528),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_420),
.B(n_344),
.Y(n_632)
);

A2O1A1Ixp33_ASAP7_75t_L g633 ( 
.A1(n_442),
.A2(n_345),
.B(n_210),
.C(n_244),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_552),
.B(n_278),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_499),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_552),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_435),
.B(n_286),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_435),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_438),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_515),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_528),
.B(n_287),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_553),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_515),
.B(n_304),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_508),
.A2(n_155),
.B1(n_285),
.B2(n_271),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_553),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_438),
.B(n_394),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_452),
.B(n_394),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_443),
.B(n_155),
.Y(n_648)
);

A2O1A1Ixp33_ASAP7_75t_L g649 ( 
.A1(n_442),
.A2(n_274),
.B(n_260),
.C(n_267),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_452),
.B(n_156),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_528),
.B(n_156),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_451),
.B(n_159),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_454),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_454),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_506),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_457),
.B(n_159),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_455),
.B(n_161),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_481),
.B(n_163),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_557),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_561),
.B(n_163),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_545),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_557),
.Y(n_662)
);

O2A1O1Ixp33_ASAP7_75t_L g663 ( 
.A1(n_494),
.A2(n_312),
.B(n_309),
.C(n_306),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_558),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_481),
.B(n_169),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_478),
.B(n_169),
.Y(n_666)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_542),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_426),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_504),
.B(n_306),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_422),
.Y(n_670)
);

NOR3xp33_ASAP7_75t_L g671 ( 
.A(n_466),
.B(n_236),
.C(n_201),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_481),
.B(n_509),
.Y(n_672)
);

A2O1A1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_518),
.A2(n_165),
.B(n_282),
.C(n_279),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_470),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_481),
.B(n_509),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_426),
.Y(n_676)
);

OAI221xp5_ASAP7_75t_L g677 ( 
.A1(n_445),
.A2(n_238),
.B1(n_222),
.B2(n_227),
.C(n_220),
.Y(n_677)
);

O2A1O1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_494),
.A2(n_551),
.B(n_429),
.C(n_522),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_484),
.B(n_171),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_558),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_481),
.B(n_173),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_422),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_542),
.B(n_174),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_472),
.Y(n_684)
);

NOR3x1_ASAP7_75t_L g685 ( 
.A(n_429),
.B(n_178),
.C(n_181),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_430),
.B(n_180),
.Y(n_686)
);

BUFx6f_ASAP7_75t_SL g687 ( 
.A(n_426),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_472),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_560),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_430),
.B(n_444),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_430),
.B(n_216),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_474),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_460),
.A2(n_240),
.B1(n_279),
.B2(n_277),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_444),
.B(n_216),
.Y(n_694)
);

NAND2x1p5_ASAP7_75t_L g695 ( 
.A(n_481),
.B(n_509),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_474),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_465),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_509),
.B(n_257),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_527),
.A2(n_285),
.B(n_257),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_498),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_465),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_509),
.B(n_263),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_444),
.B(n_263),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_L g704 ( 
.A1(n_426),
.A2(n_271),
.B1(n_270),
.B2(n_269),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_495),
.B(n_270),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_444),
.B(n_269),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_509),
.B(n_240),
.Y(n_707)
);

OR2x6_ASAP7_75t_L g708 ( 
.A(n_426),
.B(n_54),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_458),
.B(n_205),
.Y(n_709)
);

INVxp33_ASAP7_75t_L g710 ( 
.A(n_461),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_491),
.B(n_254),
.Y(n_711)
);

NOR2xp67_ASAP7_75t_L g712 ( 
.A(n_497),
.B(n_113),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_541),
.A2(n_277),
.B1(n_274),
.B2(n_273),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_565),
.B(n_473),
.Y(n_714)
);

INVx5_ASAP7_75t_L g715 ( 
.A(n_573),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_580),
.Y(n_716)
);

NOR2x1p5_ASAP7_75t_L g717 ( 
.A(n_655),
.B(n_462),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_608),
.B(n_462),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_573),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_593),
.B(n_473),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_609),
.B(n_556),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_583),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_655),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_R g724 ( 
.A(n_635),
.B(n_461),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_593),
.B(n_606),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_629),
.A2(n_460),
.B1(n_518),
.B2(n_520),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_666),
.A2(n_460),
.B1(n_479),
.B2(n_477),
.Y(n_727)
);

BUFx2_ASAP7_75t_L g728 ( 
.A(n_640),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_606),
.B(n_477),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_669),
.B(n_446),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_567),
.A2(n_446),
.B(n_535),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_589),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_609),
.A2(n_460),
.B1(n_479),
.B2(n_549),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_632),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_619),
.A2(n_460),
.B1(n_423),
.B2(n_458),
.Y(n_735)
);

AND2x2_ASAP7_75t_SL g736 ( 
.A(n_577),
.B(n_496),
.Y(n_736)
);

AND2x4_ASAP7_75t_L g737 ( 
.A(n_566),
.B(n_491),
.Y(n_737)
);

CKINVDCx8_ASAP7_75t_R g738 ( 
.A(n_683),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_R g739 ( 
.A(n_635),
.B(n_460),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_622),
.B(n_480),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_597),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_670),
.B(n_496),
.Y(n_742)
);

AND3x2_ASAP7_75t_SL g743 ( 
.A(n_673),
.B(n_273),
.C(n_267),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_582),
.B(n_458),
.Y(n_744)
);

INVx4_ASAP7_75t_L g745 ( 
.A(n_573),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_587),
.B(n_619),
.Y(n_746)
);

NAND3xp33_ASAP7_75t_SL g747 ( 
.A(n_705),
.B(n_262),
.C(n_512),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_626),
.A2(n_423),
.B1(n_459),
.B2(n_475),
.Y(n_748)
);

BUFx4f_ASAP7_75t_SL g749 ( 
.A(n_661),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_622),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_643),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_620),
.B(n_476),
.Y(n_752)
);

INVx5_ASAP7_75t_L g753 ( 
.A(n_573),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_623),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_642),
.B(n_491),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_623),
.B(n_480),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_630),
.B(n_482),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_630),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_626),
.A2(n_423),
.B1(n_475),
.B2(n_459),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_562),
.B(n_459),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_638),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_562),
.B(n_459),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_682),
.B(n_475),
.Y(n_763)
);

INVx4_ASAP7_75t_L g764 ( 
.A(n_581),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_638),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_639),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_590),
.B(n_482),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_572),
.B(n_475),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_604),
.B(n_446),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_645),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_667),
.Y(n_771)
);

INVx5_ASAP7_75t_L g772 ( 
.A(n_581),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_597),
.B(n_498),
.Y(n_773)
);

AOI21x1_ASAP7_75t_L g774 ( 
.A1(n_563),
.A2(n_559),
.B(n_555),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_570),
.A2(n_535),
.B(n_498),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_605),
.B(n_453),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_572),
.B(n_491),
.Y(n_777)
);

NAND3xp33_ASAP7_75t_L g778 ( 
.A(n_678),
.B(n_502),
.C(n_483),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_597),
.Y(n_779)
);

HB1xp67_ASAP7_75t_L g780 ( 
.A(n_585),
.Y(n_780)
);

BUFx4f_ASAP7_75t_L g781 ( 
.A(n_708),
.Y(n_781)
);

NOR2x1_ASAP7_75t_R g782 ( 
.A(n_711),
.B(n_526),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_653),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_709),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_591),
.B(n_544),
.Y(n_785)
);

AND2x4_ASAP7_75t_L g786 ( 
.A(n_596),
.B(n_599),
.Y(n_786)
);

INVx5_ASAP7_75t_L g787 ( 
.A(n_581),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_653),
.B(n_544),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_581),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_654),
.B(n_544),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_654),
.B(n_544),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_697),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_602),
.B(n_483),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_701),
.Y(n_794)
);

BUFx8_ASAP7_75t_L g795 ( 
.A(n_687),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_648),
.B(n_498),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_602),
.B(n_486),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_600),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_568),
.A2(n_453),
.B1(n_492),
.B2(n_549),
.Y(n_799)
);

AO22x1_ASAP7_75t_L g800 ( 
.A1(n_652),
.A2(n_501),
.B1(n_486),
.B2(n_540),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_650),
.B(n_555),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_607),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_602),
.B(n_488),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_624),
.B(n_488),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_612),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_617),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_618),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_636),
.A2(n_531),
.B1(n_500),
.B2(n_540),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_624),
.B(n_501),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_624),
.B(n_610),
.Y(n_810)
);

BUFx4f_ASAP7_75t_L g811 ( 
.A(n_708),
.Y(n_811)
);

NOR3xp33_ASAP7_75t_SL g812 ( 
.A(n_673),
.B(n_1),
.C(n_2),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_594),
.Y(n_813)
);

AND2x6_ASAP7_75t_SL g814 ( 
.A(n_616),
.B(n_1),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_594),
.B(n_631),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_613),
.B(n_631),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_674),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_656),
.B(n_453),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_677),
.B(n_453),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_659),
.B(n_502),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_668),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_662),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_668),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_664),
.B(n_505),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_680),
.Y(n_825)
);

NAND2x1p5_ASAP7_75t_L g826 ( 
.A(n_676),
.B(n_535),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_644),
.B(n_503),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_563),
.A2(n_505),
.B1(n_512),
.B2(n_539),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_584),
.A2(n_503),
.B(n_546),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_685),
.Y(n_830)
);

INVx5_ASAP7_75t_L g831 ( 
.A(n_676),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_689),
.B(n_532),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_646),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_588),
.A2(n_532),
.B1(n_517),
.B2(n_539),
.Y(n_834)
);

INVx5_ASAP7_75t_L g835 ( 
.A(n_700),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_588),
.A2(n_625),
.B1(n_641),
.B2(n_693),
.Y(n_836)
);

NAND2x1p5_ASAP7_75t_L g837 ( 
.A(n_700),
.B(n_503),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_674),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_647),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_660),
.B(n_712),
.Y(n_840)
);

INVx5_ASAP7_75t_L g841 ( 
.A(n_700),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_657),
.B(n_503),
.Y(n_842)
);

INVxp67_ASAP7_75t_L g843 ( 
.A(n_564),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_684),
.B(n_524),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_704),
.B(n_546),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_634),
.Y(n_846)
);

INVx5_ASAP7_75t_L g847 ( 
.A(n_688),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_679),
.B(n_546),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_651),
.B(n_526),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_692),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_692),
.B(n_524),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_696),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_696),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_651),
.B(n_526),
.Y(n_854)
);

OAI221xp5_ASAP7_75t_L g855 ( 
.A1(n_649),
.A2(n_449),
.B1(n_427),
.B2(n_428),
.C(n_433),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_637),
.B(n_559),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_690),
.Y(n_857)
);

INVx6_ASAP7_75t_L g858 ( 
.A(n_710),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_574),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_687),
.A2(n_537),
.B1(n_531),
.B2(n_529),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_687),
.A2(n_537),
.B1(n_529),
.B2(n_546),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_575),
.Y(n_862)
);

INVxp67_ASAP7_75t_L g863 ( 
.A(n_671),
.Y(n_863)
);

NAND2x1p5_ASAP7_75t_L g864 ( 
.A(n_672),
.B(n_675),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_649),
.B(n_546),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_576),
.B(n_463),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_578),
.B(n_463),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_579),
.B(n_449),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_586),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_601),
.Y(n_870)
);

O2A1O1Ixp5_ASAP7_75t_L g871 ( 
.A1(n_592),
.A2(n_441),
.B(n_440),
.C(n_439),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_746),
.B(n_710),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_715),
.A2(n_695),
.B(n_675),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_715),
.A2(n_695),
.B(n_672),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_752),
.B(n_686),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_786),
.B(n_625),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_767),
.B(n_691),
.Y(n_877)
);

AND2x2_ASAP7_75t_SL g878 ( 
.A(n_736),
.B(n_598),
.Y(n_878)
);

AOI21x1_ASAP7_75t_L g879 ( 
.A1(n_800),
.A2(n_796),
.B(n_848),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_726),
.A2(n_633),
.B1(n_641),
.B2(n_569),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_714),
.B(n_694),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_714),
.A2(n_706),
.B1(n_703),
.B2(n_603),
.Y(n_882)
);

BUFx2_ASAP7_75t_L g883 ( 
.A(n_728),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_734),
.B(n_751),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_813),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_833),
.B(n_633),
.Y(n_886)
);

INVx4_ASAP7_75t_L g887 ( 
.A(n_715),
.Y(n_887)
);

BUFx12f_ASAP7_75t_L g888 ( 
.A(n_795),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_718),
.B(n_713),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_813),
.Y(n_890)
);

BUFx12f_ASAP7_75t_L g891 ( 
.A(n_795),
.Y(n_891)
);

AND2x4_ASAP7_75t_L g892 ( 
.A(n_786),
.B(n_770),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_715),
.A2(n_595),
.B(n_615),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_839),
.B(n_611),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_753),
.A2(n_615),
.B(n_595),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_SL g896 ( 
.A1(n_818),
.A2(n_614),
.B(n_699),
.C(n_627),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_742),
.B(n_621),
.Y(n_897)
);

OR2x6_ASAP7_75t_L g898 ( 
.A(n_858),
.B(n_707),
.Y(n_898)
);

INVx4_ASAP7_75t_L g899 ( 
.A(n_753),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_753),
.A2(n_592),
.B(n_621),
.Y(n_900)
);

OAI22xp5_ASAP7_75t_L g901 ( 
.A1(n_781),
.A2(n_707),
.B1(n_628),
.B2(n_698),
.Y(n_901)
);

OR2x6_ASAP7_75t_L g902 ( 
.A(n_858),
.B(n_663),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_723),
.Y(n_903)
);

NAND2x1_ASAP7_75t_L g904 ( 
.A(n_745),
.B(n_441),
.Y(n_904)
);

O2A1O1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_843),
.A2(n_571),
.B(n_698),
.C(n_681),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_816),
.B(n_702),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_753),
.A2(n_702),
.B(n_681),
.Y(n_907)
);

OAI22xp5_ASAP7_75t_L g908 ( 
.A1(n_816),
.A2(n_665),
.B1(n_658),
.B2(n_440),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_846),
.B(n_665),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_781),
.A2(n_439),
.B1(n_433),
.B2(n_428),
.Y(n_910)
);

BUFx2_ASAP7_75t_L g911 ( 
.A(n_830),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_811),
.A2(n_427),
.B1(n_421),
.B2(n_6),
.Y(n_912)
);

AOI22xp33_ASAP7_75t_L g913 ( 
.A1(n_747),
.A2(n_421),
.B1(n_3),
.B2(n_7),
.Y(n_913)
);

BUFx2_ASAP7_75t_L g914 ( 
.A(n_724),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_772),
.A2(n_141),
.B(n_134),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_719),
.Y(n_916)
);

INVx4_ASAP7_75t_L g917 ( 
.A(n_772),
.Y(n_917)
);

BUFx2_ASAP7_75t_L g918 ( 
.A(n_739),
.Y(n_918)
);

O2A1O1Ixp5_ASAP7_75t_L g919 ( 
.A1(n_840),
.A2(n_126),
.B(n_122),
.C(n_117),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_815),
.B(n_3),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_772),
.A2(n_787),
.B(n_810),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_863),
.A2(n_7),
.B(n_11),
.C(n_13),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_815),
.B(n_784),
.Y(n_923)
);

AOI21x1_ASAP7_75t_L g924 ( 
.A1(n_725),
.A2(n_115),
.B(n_110),
.Y(n_924)
);

INVx1_ASAP7_75t_SL g925 ( 
.A(n_865),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_716),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_738),
.B(n_16),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_719),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_754),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_L g930 ( 
.A1(n_741),
.A2(n_98),
.B1(n_97),
.B2(n_92),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_780),
.B(n_17),
.Y(n_931)
);

O2A1O1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_763),
.A2(n_802),
.B(n_798),
.C(n_807),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_761),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_722),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_772),
.A2(n_84),
.B(n_67),
.Y(n_935)
);

INVx4_ASAP7_75t_L g936 ( 
.A(n_787),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_778),
.A2(n_65),
.B(n_62),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_766),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_732),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_779),
.B(n_57),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_805),
.B(n_20),
.Y(n_941)
);

NOR2xp67_ASAP7_75t_SL g942 ( 
.A(n_787),
.B(n_20),
.Y(n_942)
);

INVx4_ASAP7_75t_L g943 ( 
.A(n_787),
.Y(n_943)
);

NAND3xp33_ASAP7_75t_SL g944 ( 
.A(n_771),
.B(n_22),
.C(n_24),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_810),
.A2(n_51),
.B(n_28),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_865),
.Y(n_946)
);

OAI21xp33_ASAP7_75t_L g947 ( 
.A1(n_806),
.A2(n_32),
.B(n_35),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_789),
.B(n_40),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_778),
.A2(n_45),
.B(n_48),
.Y(n_949)
);

A2O1A1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_819),
.A2(n_49),
.B(n_50),
.C(n_51),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_750),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_SL g952 ( 
.A(n_811),
.B(n_745),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_731),
.A2(n_775),
.B(n_773),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_769),
.A2(n_809),
.B(n_804),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_836),
.A2(n_827),
.B1(n_725),
.B2(n_733),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_859),
.B(n_870),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_758),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_776),
.A2(n_861),
.B1(n_727),
.B2(n_860),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_721),
.B(n_755),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_765),
.Y(n_960)
);

OR2x6_ASAP7_75t_SL g961 ( 
.A(n_743),
.B(n_801),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_831),
.A2(n_854),
.B1(n_849),
.B2(n_744),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_721),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_822),
.B(n_825),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_783),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_793),
.A2(n_797),
.B(n_809),
.Y(n_966)
);

OAI21xp5_ASAP7_75t_L g967 ( 
.A1(n_871),
.A2(n_803),
.B(n_855),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_792),
.A2(n_794),
.B(n_812),
.C(n_845),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_737),
.B(n_717),
.Y(n_969)
);

BUFx4f_ASAP7_75t_L g970 ( 
.A(n_821),
.Y(n_970)
);

NAND2x1_ASAP7_75t_L g971 ( 
.A(n_764),
.B(n_789),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_803),
.A2(n_842),
.B(n_868),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_737),
.B(n_823),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_867),
.A2(n_856),
.B(n_730),
.Y(n_974)
);

BUFx3_ASAP7_75t_L g975 ( 
.A(n_749),
.Y(n_975)
);

INVx6_ASAP7_75t_L g976 ( 
.A(n_821),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_829),
.A2(n_768),
.B(n_762),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_831),
.A2(n_821),
.B1(n_823),
.B2(n_764),
.Y(n_978)
);

O2A1O1Ixp5_ASAP7_75t_L g979 ( 
.A1(n_862),
.A2(n_774),
.B(n_824),
.C(n_832),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_789),
.Y(n_980)
);

OAI21xp33_ASAP7_75t_L g981 ( 
.A1(n_720),
.A2(n_729),
.B(n_757),
.Y(n_981)
);

INVx6_ASAP7_75t_L g982 ( 
.A(n_823),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_760),
.A2(n_777),
.B(n_740),
.Y(n_983)
);

O2A1O1Ixp5_ASAP7_75t_L g984 ( 
.A1(n_862),
.A2(n_824),
.B(n_820),
.C(n_832),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_785),
.A2(n_820),
.B(n_740),
.C(n_757),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_869),
.B(n_857),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_869),
.B(n_857),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_866),
.B(n_720),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_756),
.A2(n_791),
.B(n_790),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_756),
.A2(n_791),
.B(n_790),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_903),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_872),
.B(n_831),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_964),
.Y(n_993)
);

OAI21x1_ASAP7_75t_L g994 ( 
.A1(n_953),
.A2(n_844),
.B(n_851),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_883),
.B(n_817),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_L g996 ( 
.A1(n_925),
.A2(n_831),
.B1(n_847),
.B2(n_735),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_SL g997 ( 
.A1(n_955),
.A2(n_782),
.B(n_826),
.Y(n_997)
);

BUFx12f_ASAP7_75t_L g998 ( 
.A(n_888),
.Y(n_998)
);

INVx1_ASAP7_75t_SL g999 ( 
.A(n_911),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_889),
.A2(n_748),
.B(n_759),
.C(n_729),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_877),
.B(n_866),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_R g1002 ( 
.A(n_914),
.B(n_850),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_925),
.A2(n_847),
.B1(n_826),
.B2(n_864),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_972),
.A2(n_847),
.B(n_788),
.Y(n_1004)
);

OAI21xp33_ASAP7_75t_L g1005 ( 
.A1(n_913),
.A2(n_743),
.B(n_788),
.Y(n_1005)
);

BUFx2_ASAP7_75t_L g1006 ( 
.A(n_963),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_954),
.A2(n_847),
.B(n_844),
.Y(n_1007)
);

AOI21x1_ASAP7_75t_L g1008 ( 
.A1(n_879),
.A2(n_962),
.B(n_983),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_959),
.B(n_838),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_881),
.B(n_852),
.Y(n_1010)
);

OAI21x1_ASAP7_75t_L g1011 ( 
.A1(n_989),
.A2(n_851),
.B(n_834),
.Y(n_1011)
);

NAND3xp33_ASAP7_75t_L g1012 ( 
.A(n_950),
.B(n_808),
.C(n_799),
.Y(n_1012)
);

NAND3xp33_ASAP7_75t_SL g1013 ( 
.A(n_922),
.B(n_814),
.C(n_828),
.Y(n_1013)
);

AND3x4_ASAP7_75t_L g1014 ( 
.A(n_975),
.B(n_853),
.C(n_864),
.Y(n_1014)
);

OAI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_906),
.A2(n_837),
.B(n_835),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_946),
.A2(n_835),
.B1(n_841),
.B2(n_837),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_946),
.A2(n_835),
.B1(n_841),
.B2(n_878),
.Y(n_1017)
);

NAND3x1_ASAP7_75t_L g1018 ( 
.A(n_927),
.B(n_841),
.C(n_969),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_884),
.B(n_961),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_897),
.B(n_875),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_959),
.Y(n_1021)
);

AO32x2_ASAP7_75t_L g1022 ( 
.A1(n_912),
.A2(n_880),
.A3(n_901),
.B1(n_908),
.B2(n_882),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_923),
.B(n_892),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_988),
.B(n_981),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_990),
.A2(n_985),
.B(n_981),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_892),
.B(n_973),
.Y(n_1026)
);

AO31x2_ASAP7_75t_L g1027 ( 
.A1(n_901),
.A2(n_912),
.A3(n_974),
.B(n_910),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_967),
.A2(n_896),
.B(n_893),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_894),
.B(n_886),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_967),
.A2(n_895),
.B(n_984),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_902),
.B(n_931),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_956),
.A2(n_909),
.B1(n_876),
.B2(n_918),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_902),
.B(n_876),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_L g1034 ( 
.A1(n_979),
.A2(n_921),
.B(n_907),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_905),
.A2(n_968),
.B(n_900),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_910),
.A2(n_904),
.B(n_874),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_987),
.B(n_986),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_929),
.B(n_933),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_887),
.A2(n_936),
.B(n_917),
.Y(n_1039)
);

NAND2x1p5_ASAP7_75t_L g1040 ( 
.A(n_887),
.B(n_917),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_873),
.A2(n_924),
.B(n_932),
.Y(n_1041)
);

INVx3_ASAP7_75t_L g1042 ( 
.A(n_899),
.Y(n_1042)
);

AOI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_898),
.A2(n_952),
.B1(n_940),
.B2(n_948),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_938),
.B(n_926),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_934),
.B(n_951),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_939),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_899),
.A2(n_943),
.B(n_936),
.Y(n_1047)
);

NOR2x1_ASAP7_75t_L g1048 ( 
.A(n_943),
.B(n_978),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_957),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_960),
.B(n_965),
.Y(n_1050)
);

OAI22x1_ASAP7_75t_L g1051 ( 
.A1(n_920),
.A2(n_941),
.B1(n_940),
.B2(n_949),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_885),
.B(n_890),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_947),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_937),
.A2(n_919),
.B(n_971),
.Y(n_1054)
);

AO31x2_ASAP7_75t_L g1055 ( 
.A1(n_945),
.A2(n_930),
.A3(n_935),
.B(n_915),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_898),
.B(n_885),
.Y(n_1056)
);

AND2x6_ASAP7_75t_SL g1057 ( 
.A(n_891),
.B(n_944),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_952),
.A2(n_970),
.B(n_916),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_SL g1059 ( 
.A1(n_942),
.A2(n_916),
.B(n_928),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_885),
.B(n_890),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_928),
.A2(n_980),
.B(n_976),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_928),
.B(n_980),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_980),
.B(n_976),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_982),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_887),
.Y(n_1065)
);

NAND3xp33_ASAP7_75t_L g1066 ( 
.A(n_889),
.B(n_629),
.C(n_587),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_972),
.A2(n_954),
.B(n_955),
.Y(n_1067)
);

NAND3xp33_ASAP7_75t_SL g1068 ( 
.A(n_889),
.B(n_629),
.C(n_577),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_872),
.B(n_734),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_955),
.A2(n_565),
.B(n_906),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_964),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_955),
.A2(n_565),
.B(n_906),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_877),
.B(n_565),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_877),
.B(n_565),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_883),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_877),
.B(n_565),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_964),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_872),
.B(n_608),
.Y(n_1078)
);

NOR2x1_ASAP7_75t_SL g1079 ( 
.A(n_887),
.B(n_899),
.Y(n_1079)
);

AOI21xp33_ASAP7_75t_L g1080 ( 
.A1(n_889),
.A2(n_629),
.B(n_587),
.Y(n_1080)
);

NAND2xp33_ASAP7_75t_R g1081 ( 
.A(n_903),
.B(n_462),
.Y(n_1081)
);

AO21x1_ASAP7_75t_L g1082 ( 
.A1(n_937),
.A2(n_949),
.B(n_880),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_887),
.Y(n_1083)
);

AOI21x1_ASAP7_75t_L g1084 ( 
.A1(n_879),
.A2(n_800),
.B(n_954),
.Y(n_1084)
);

AO21x2_ASAP7_75t_L g1085 ( 
.A1(n_967),
.A2(n_962),
.B(n_972),
.Y(n_1085)
);

NOR2xp67_ASAP7_75t_L g1086 ( 
.A(n_903),
.B(n_462),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_877),
.B(n_565),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_972),
.A2(n_954),
.B(n_955),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_SL g1089 ( 
.A1(n_955),
.A2(n_687),
.B(n_958),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_953),
.A2(n_977),
.B(n_966),
.Y(n_1090)
);

NAND2x1p5_ASAP7_75t_L g1091 ( 
.A(n_887),
.B(n_715),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_877),
.B(n_565),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_955),
.A2(n_565),
.B(n_906),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_964),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_964),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_872),
.B(n_734),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_872),
.B(n_608),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1073),
.B(n_1074),
.Y(n_1098)
);

BUFx12f_ASAP7_75t_L g1099 ( 
.A(n_998),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1038),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_1081),
.Y(n_1101)
);

OR2x2_ASAP7_75t_L g1102 ( 
.A(n_1020),
.B(n_1069),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1034),
.A2(n_1036),
.B(n_994),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_1042),
.Y(n_1104)
);

OR2x2_ASAP7_75t_L g1105 ( 
.A(n_1020),
.B(n_1096),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1050),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_1080),
.B(n_1078),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1050),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_1097),
.B(n_1073),
.Y(n_1109)
);

O2A1O1Ixp33_ASAP7_75t_SL g1110 ( 
.A1(n_1000),
.A2(n_1072),
.B(n_1070),
.C(n_1093),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_1074),
.A2(n_1076),
.B(n_1087),
.C(n_1092),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_1013),
.A2(n_1053),
.B1(n_1051),
.B2(n_1005),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_1033),
.B(n_1009),
.Y(n_1113)
);

OR2x2_ASAP7_75t_L g1114 ( 
.A(n_1037),
.B(n_993),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1026),
.B(n_1031),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1014),
.A2(n_1043),
.B1(n_1094),
.B2(n_1095),
.Y(n_1116)
);

AOI22xp33_ASAP7_75t_L g1117 ( 
.A1(n_1071),
.A2(n_1077),
.B1(n_1019),
.B2(n_1032),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1021),
.B(n_1023),
.Y(n_1118)
);

NOR2xp67_ASAP7_75t_L g1119 ( 
.A(n_991),
.B(n_1086),
.Y(n_1119)
);

NOR2xp67_ASAP7_75t_L g1120 ( 
.A(n_995),
.B(n_1075),
.Y(n_1120)
);

INVxp67_ASAP7_75t_SL g1121 ( 
.A(n_1037),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_1012),
.A2(n_1035),
.B1(n_1001),
.B2(n_1029),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_1001),
.B(n_1044),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_1063),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_1029),
.B(n_1010),
.Y(n_1125)
);

NAND2x1p5_ASAP7_75t_L g1126 ( 
.A(n_1048),
.B(n_1042),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1090),
.A2(n_1007),
.B(n_1004),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1007),
.A2(n_1004),
.B(n_1041),
.Y(n_1128)
);

NOR2xp67_ASAP7_75t_SL g1129 ( 
.A(n_997),
.B(n_1089),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_1063),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1044),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_999),
.A2(n_1010),
.B1(n_1018),
.B2(n_1006),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1011),
.A2(n_1084),
.B(n_1028),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1028),
.A2(n_1008),
.B(n_1088),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1046),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_1009),
.B(n_1058),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1024),
.A2(n_1015),
.B(n_1030),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_1030),
.A2(n_1054),
.B(n_1003),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1045),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_992),
.A2(n_1017),
.B(n_996),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_1002),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_1039),
.A2(n_1047),
.B(n_1016),
.Y(n_1142)
);

AO21x2_ASAP7_75t_L g1143 ( 
.A1(n_1085),
.A2(n_1059),
.B(n_1022),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1040),
.A2(n_1091),
.B(n_1045),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1040),
.A2(n_1091),
.B(n_1061),
.Y(n_1145)
);

INVx2_ASAP7_75t_SL g1146 ( 
.A(n_1064),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1065),
.A2(n_1083),
.B(n_1049),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_1065),
.A2(n_1083),
.B(n_1062),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1052),
.A2(n_1060),
.B(n_1056),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1085),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_1055),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_1079),
.B(n_1027),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_1057),
.Y(n_1153)
);

INVx1_ASAP7_75t_SL g1154 ( 
.A(n_1027),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_SL g1155 ( 
.A1(n_1080),
.A2(n_950),
.B(n_949),
.C(n_937),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1038),
.Y(n_1156)
);

O2A1O1Ixp33_ASAP7_75t_SL g1157 ( 
.A1(n_1080),
.A2(n_950),
.B(n_949),
.C(n_937),
.Y(n_1157)
);

INVx1_ASAP7_75t_SL g1158 ( 
.A(n_999),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1080),
.A2(n_1066),
.B1(n_1068),
.B2(n_736),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1080),
.A2(n_1066),
.B1(n_1068),
.B2(n_736),
.Y(n_1160)
);

OA21x2_ASAP7_75t_L g1161 ( 
.A1(n_1025),
.A2(n_1088),
.B(n_1067),
.Y(n_1161)
);

OA21x2_ASAP7_75t_L g1162 ( 
.A1(n_1025),
.A2(n_1088),
.B(n_1067),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1080),
.B(n_1066),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_1081),
.Y(n_1164)
);

O2A1O1Ixp5_ASAP7_75t_L g1165 ( 
.A1(n_1082),
.A2(n_1080),
.B(n_1066),
.C(n_1072),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_1080),
.B(n_1066),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1080),
.A2(n_1066),
.B1(n_1068),
.B2(n_736),
.Y(n_1167)
);

OA21x2_ASAP7_75t_L g1168 ( 
.A1(n_1025),
.A2(n_1088),
.B(n_1067),
.Y(n_1168)
);

INVx2_ASAP7_75t_SL g1169 ( 
.A(n_991),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_SL g1170 ( 
.A1(n_1082),
.A2(n_949),
.B(n_968),
.Y(n_1170)
);

OA21x2_ASAP7_75t_L g1171 ( 
.A1(n_1025),
.A2(n_1088),
.B(n_1067),
.Y(n_1171)
);

O2A1O1Ixp5_ASAP7_75t_L g1172 ( 
.A1(n_1082),
.A2(n_1080),
.B(n_1066),
.C(n_1072),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1038),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1038),
.Y(n_1174)
);

INVx5_ASAP7_75t_L g1175 ( 
.A(n_1042),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1034),
.A2(n_1036),
.B(n_994),
.Y(n_1176)
);

OR2x2_ASAP7_75t_L g1177 ( 
.A(n_1020),
.B(n_1069),
.Y(n_1177)
);

AOI21xp33_ASAP7_75t_L g1178 ( 
.A1(n_1066),
.A2(n_1080),
.B(n_629),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1080),
.A2(n_1066),
.B(n_1072),
.C(n_1070),
.Y(n_1179)
);

O2A1O1Ixp33_ASAP7_75t_SL g1180 ( 
.A1(n_1080),
.A2(n_950),
.B(n_949),
.C(n_937),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_1002),
.Y(n_1181)
);

NAND3xp33_ASAP7_75t_L g1182 ( 
.A(n_1066),
.B(n_1080),
.C(n_629),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1034),
.A2(n_1036),
.B(n_994),
.Y(n_1183)
);

CKINVDCx11_ASAP7_75t_R g1184 ( 
.A(n_998),
.Y(n_1184)
);

O2A1O1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1178),
.A2(n_1179),
.B(n_1166),
.C(n_1163),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1109),
.B(n_1098),
.Y(n_1186)
);

O2A1O1Ixp5_ASAP7_75t_L g1187 ( 
.A1(n_1165),
.A2(n_1172),
.B(n_1179),
.C(n_1166),
.Y(n_1187)
);

O2A1O1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1163),
.A2(n_1157),
.B(n_1155),
.C(n_1180),
.Y(n_1188)
);

O2A1O1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_1155),
.A2(n_1180),
.B(n_1157),
.C(n_1110),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1115),
.B(n_1118),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1102),
.B(n_1105),
.Y(n_1191)
);

AND2x6_ASAP7_75t_L g1192 ( 
.A(n_1136),
.B(n_1152),
.Y(n_1192)
);

INVx1_ASAP7_75t_SL g1193 ( 
.A(n_1158),
.Y(n_1193)
);

O2A1O1Ixp5_ASAP7_75t_L g1194 ( 
.A1(n_1129),
.A2(n_1182),
.B(n_1107),
.C(n_1140),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_1124),
.Y(n_1195)
);

OA21x2_ASAP7_75t_L g1196 ( 
.A1(n_1134),
.A2(n_1128),
.B(n_1127),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1154),
.B(n_1143),
.Y(n_1197)
);

CKINVDCx16_ASAP7_75t_R g1198 ( 
.A(n_1099),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1109),
.B(n_1121),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1159),
.A2(n_1160),
.B1(n_1167),
.B2(n_1117),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1159),
.A2(n_1160),
.B1(n_1167),
.B2(n_1117),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1177),
.B(n_1113),
.Y(n_1202)
);

O2A1O1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1111),
.A2(n_1116),
.B(n_1170),
.C(n_1132),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_1124),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_1143),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_1181),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1141),
.A2(n_1112),
.B1(n_1164),
.B2(n_1101),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1149),
.B(n_1114),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1111),
.B(n_1123),
.Y(n_1209)
);

AOI21x1_ASAP7_75t_SL g1210 ( 
.A1(n_1153),
.A2(n_1164),
.B(n_1101),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1100),
.B(n_1156),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1173),
.B(n_1174),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1135),
.B(n_1148),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1141),
.A2(n_1120),
.B1(n_1122),
.B2(n_1153),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1106),
.B(n_1108),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1131),
.A2(n_1119),
.B1(n_1146),
.B2(n_1125),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1139),
.B(n_1135),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1124),
.B(n_1130),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1137),
.B(n_1130),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1130),
.B(n_1104),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1126),
.A2(n_1169),
.B1(n_1130),
.B2(n_1175),
.Y(n_1221)
);

O2A1O1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1126),
.A2(n_1151),
.B(n_1150),
.C(n_1104),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_R g1223 ( 
.A(n_1184),
.B(n_1099),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_1148),
.B(n_1147),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_SL g1225 ( 
.A1(n_1161),
.A2(n_1162),
.B(n_1168),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1175),
.B(n_1144),
.Y(n_1226)
);

OA21x2_ASAP7_75t_L g1227 ( 
.A1(n_1128),
.A2(n_1127),
.B(n_1138),
.Y(n_1227)
);

OA21x2_ASAP7_75t_L g1228 ( 
.A1(n_1133),
.A2(n_1103),
.B(n_1183),
.Y(n_1228)
);

AOI21x1_ASAP7_75t_SL g1229 ( 
.A1(n_1184),
.A2(n_1142),
.B(n_1145),
.Y(n_1229)
);

CKINVDCx6p67_ASAP7_75t_R g1230 ( 
.A(n_1147),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1171),
.Y(n_1231)
);

OA21x2_ASAP7_75t_L g1232 ( 
.A1(n_1176),
.A2(n_1134),
.B(n_1128),
.Y(n_1232)
);

AOI221x1_ASAP7_75t_SL g1233 ( 
.A1(n_1178),
.A2(n_478),
.B1(n_1080),
.B2(n_1107),
.C(n_1066),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_1143),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1115),
.B(n_1118),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1115),
.B(n_1118),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1159),
.A2(n_736),
.B1(n_1066),
.B2(n_629),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_SL g1238 ( 
.A1(n_1179),
.A2(n_937),
.B(n_949),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1159),
.A2(n_736),
.B1(n_1066),
.B2(n_629),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1136),
.B(n_1149),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1159),
.A2(n_736),
.B1(n_1066),
.B2(n_629),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_SL g1242 ( 
.A(n_1141),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1163),
.A2(n_1080),
.B(n_1066),
.C(n_1166),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1115),
.B(n_1118),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1115),
.B(n_1118),
.Y(n_1245)
);

O2A1O1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1178),
.A2(n_1080),
.B(n_1068),
.C(n_629),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_1184),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1115),
.B(n_1118),
.Y(n_1248)
);

CKINVDCx20_ASAP7_75t_R g1249 ( 
.A(n_1184),
.Y(n_1249)
);

A2O1A1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1163),
.A2(n_1080),
.B(n_1066),
.C(n_1166),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_1143),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1213),
.Y(n_1252)
);

NAND3xp33_ASAP7_75t_L g1253 ( 
.A(n_1243),
.B(n_1250),
.C(n_1185),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1213),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1213),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1192),
.Y(n_1256)
);

OR2x6_ASAP7_75t_L g1257 ( 
.A(n_1238),
.B(n_1225),
.Y(n_1257)
);

OR2x6_ASAP7_75t_L g1258 ( 
.A(n_1238),
.B(n_1225),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1231),
.B(n_1240),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1205),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1208),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_1192),
.Y(n_1262)
);

INVx1_ASAP7_75t_SL g1263 ( 
.A(n_1199),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_1234),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1231),
.B(n_1240),
.Y(n_1265)
);

OR2x2_ASAP7_75t_L g1266 ( 
.A(n_1251),
.B(n_1197),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1209),
.B(n_1243),
.Y(n_1267)
);

OR2x6_ASAP7_75t_L g1268 ( 
.A(n_1240),
.B(n_1189),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1251),
.Y(n_1269)
);

AOI221xp5_ASAP7_75t_L g1270 ( 
.A1(n_1237),
.A2(n_1239),
.B1(n_1241),
.B2(n_1233),
.C(n_1200),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1224),
.Y(n_1271)
);

OR2x6_ASAP7_75t_L g1272 ( 
.A(n_1222),
.B(n_1188),
.Y(n_1272)
);

AOI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1228),
.A2(n_1232),
.B(n_1196),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1186),
.B(n_1211),
.Y(n_1274)
);

OA21x2_ASAP7_75t_L g1275 ( 
.A1(n_1187),
.A2(n_1194),
.B(n_1219),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1230),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1217),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1191),
.B(n_1192),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1226),
.Y(n_1279)
);

BUFx12f_ASAP7_75t_L g1280 ( 
.A(n_1247),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1228),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1229),
.A2(n_1227),
.B(n_1196),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1212),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1221),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1215),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1232),
.Y(n_1286)
);

OAI211xp5_ASAP7_75t_SL g1287 ( 
.A1(n_1270),
.A2(n_1246),
.B(n_1203),
.C(n_1201),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1260),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_1260),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1263),
.B(n_1216),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1264),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_1271),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1281),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1253),
.B(n_1270),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1256),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1263),
.B(n_1190),
.Y(n_1296)
);

OAI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1253),
.A2(n_1214),
.B1(n_1207),
.B2(n_1198),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1267),
.A2(n_1202),
.B1(n_1206),
.B2(n_1235),
.Y(n_1298)
);

OR2x2_ASAP7_75t_L g1299 ( 
.A(n_1266),
.B(n_1196),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1252),
.B(n_1254),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1254),
.B(n_1245),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1267),
.A2(n_1236),
.B1(n_1244),
.B2(n_1248),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1255),
.B(n_1220),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1255),
.B(n_1218),
.Y(n_1304)
);

OR2x2_ASAP7_75t_L g1305 ( 
.A(n_1266),
.B(n_1261),
.Y(n_1305)
);

INVxp67_ASAP7_75t_SL g1306 ( 
.A(n_1264),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1269),
.Y(n_1307)
);

NAND2x1p5_ASAP7_75t_L g1308 ( 
.A(n_1256),
.B(n_1262),
.Y(n_1308)
);

AO22x1_ASAP7_75t_L g1309 ( 
.A1(n_1284),
.A2(n_1247),
.B1(n_1195),
.B2(n_1204),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1286),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1288),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1294),
.B(n_1296),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1300),
.B(n_1259),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1288),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1308),
.Y(n_1315)
);

AOI221xp5_ASAP7_75t_L g1316 ( 
.A1(n_1294),
.A2(n_1274),
.B1(n_1283),
.B2(n_1285),
.C(n_1193),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1310),
.Y(n_1317)
);

OR2x6_ASAP7_75t_L g1318 ( 
.A(n_1308),
.B(n_1257),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1287),
.A2(n_1297),
.B1(n_1284),
.B2(n_1275),
.Y(n_1319)
);

OR2x2_ASAP7_75t_L g1320 ( 
.A(n_1305),
.B(n_1266),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1287),
.A2(n_1275),
.B1(n_1272),
.B2(n_1284),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1300),
.B(n_1259),
.Y(n_1322)
);

NAND3xp33_ASAP7_75t_L g1323 ( 
.A(n_1297),
.B(n_1275),
.C(n_1257),
.Y(n_1323)
);

OR2x6_ASAP7_75t_L g1324 ( 
.A(n_1308),
.B(n_1257),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1289),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1289),
.Y(n_1326)
);

OAI221xp5_ASAP7_75t_SL g1327 ( 
.A1(n_1302),
.A2(n_1272),
.B1(n_1258),
.B2(n_1257),
.C(n_1284),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1295),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1291),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1298),
.A2(n_1275),
.B1(n_1257),
.B2(n_1258),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1298),
.A2(n_1275),
.B1(n_1257),
.B2(n_1258),
.Y(n_1331)
);

NAND3xp33_ASAP7_75t_L g1332 ( 
.A(n_1290),
.B(n_1275),
.C(n_1258),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1295),
.A2(n_1258),
.B1(n_1257),
.B2(n_1272),
.Y(n_1333)
);

BUFx2_ASAP7_75t_L g1334 ( 
.A(n_1308),
.Y(n_1334)
);

A2O1A1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1290),
.A2(n_1295),
.B(n_1302),
.C(n_1256),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1304),
.B(n_1265),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_1295),
.Y(n_1337)
);

NAND3xp33_ASAP7_75t_L g1338 ( 
.A(n_1309),
.B(n_1258),
.C(n_1272),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1301),
.A2(n_1258),
.B1(n_1272),
.B2(n_1265),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1307),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1304),
.B(n_1265),
.Y(n_1341)
);

AOI221xp5_ASAP7_75t_L g1342 ( 
.A1(n_1309),
.A2(n_1274),
.B1(n_1283),
.B2(n_1285),
.C(n_1277),
.Y(n_1342)
);

OAI221xp5_ASAP7_75t_L g1343 ( 
.A1(n_1306),
.A2(n_1272),
.B1(n_1268),
.B2(n_1276),
.C(n_1279),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1304),
.B(n_1303),
.Y(n_1344)
);

OA21x2_ASAP7_75t_L g1345 ( 
.A1(n_1323),
.A2(n_1286),
.B(n_1282),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1318),
.Y(n_1346)
);

OA21x2_ASAP7_75t_L g1347 ( 
.A1(n_1323),
.A2(n_1332),
.B(n_1286),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1314),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1344),
.B(n_1292),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1311),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1311),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_1318),
.Y(n_1352)
);

OA21x2_ASAP7_75t_L g1353 ( 
.A1(n_1317),
.A2(n_1273),
.B(n_1293),
.Y(n_1353)
);

INVx1_ASAP7_75t_SL g1354 ( 
.A(n_1315),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1320),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1314),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1325),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1316),
.B(n_1278),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1325),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1326),
.B(n_1299),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1312),
.B(n_1305),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1329),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1344),
.B(n_1292),
.Y(n_1363)
);

OR2x6_ASAP7_75t_L g1364 ( 
.A(n_1318),
.B(n_1309),
.Y(n_1364)
);

INVx3_ASAP7_75t_SL g1365 ( 
.A(n_1318),
.Y(n_1365)
);

NAND3xp33_ASAP7_75t_L g1366 ( 
.A(n_1347),
.B(n_1319),
.C(n_1321),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1361),
.B(n_1280),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1346),
.B(n_1315),
.Y(n_1368)
);

OR2x2_ASAP7_75t_L g1369 ( 
.A(n_1355),
.B(n_1340),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1361),
.B(n_1316),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1356),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1346),
.B(n_1352),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_1350),
.Y(n_1373)
);

NOR2x1_ASAP7_75t_L g1374 ( 
.A(n_1358),
.B(n_1338),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1346),
.B(n_1334),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1356),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1352),
.B(n_1334),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1358),
.A2(n_1321),
.B1(n_1338),
.B2(n_1330),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1352),
.B(n_1318),
.Y(n_1379)
);

INVx1_ASAP7_75t_SL g1380 ( 
.A(n_1365),
.Y(n_1380)
);

AND2x4_ASAP7_75t_L g1381 ( 
.A(n_1364),
.B(n_1324),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1356),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1365),
.B(n_1324),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1362),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1362),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1365),
.B(n_1324),
.Y(n_1386)
);

AND2x4_ASAP7_75t_L g1387 ( 
.A(n_1364),
.B(n_1324),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1365),
.B(n_1324),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1355),
.B(n_1342),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1348),
.B(n_1342),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1364),
.B(n_1313),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1362),
.Y(n_1392)
);

INVx1_ASAP7_75t_SL g1393 ( 
.A(n_1354),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1364),
.B(n_1313),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1354),
.B(n_1280),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1353),
.Y(n_1396)
);

INVxp67_ASAP7_75t_SL g1397 ( 
.A(n_1350),
.Y(n_1397)
);

AOI21xp33_ASAP7_75t_L g1398 ( 
.A1(n_1347),
.A2(n_1335),
.B(n_1343),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1364),
.B(n_1322),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1364),
.B(n_1322),
.Y(n_1400)
);

INVxp67_ASAP7_75t_L g1401 ( 
.A(n_1357),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1357),
.B(n_1336),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1374),
.A2(n_1327),
.B1(n_1331),
.B2(n_1333),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1372),
.B(n_1364),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1390),
.B(n_1360),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1371),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1371),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1376),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1370),
.B(n_1341),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1376),
.Y(n_1410)
);

NAND4xp25_ASAP7_75t_L g1411 ( 
.A(n_1366),
.B(n_1327),
.C(n_1339),
.D(n_1343),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1382),
.Y(n_1412)
);

INVx2_ASAP7_75t_SL g1413 ( 
.A(n_1372),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1393),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1382),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1384),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1384),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1374),
.B(n_1349),
.Y(n_1418)
);

NAND2x1_ASAP7_75t_L g1419 ( 
.A(n_1381),
.B(n_1347),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1373),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1383),
.B(n_1349),
.Y(n_1421)
);

AOI21xp33_ASAP7_75t_L g1422 ( 
.A1(n_1366),
.A2(n_1347),
.B(n_1345),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1389),
.B(n_1341),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1383),
.B(n_1349),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1385),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1386),
.B(n_1363),
.Y(n_1426)
);

AOI21xp33_ASAP7_75t_L g1427 ( 
.A1(n_1380),
.A2(n_1347),
.B(n_1345),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1385),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1392),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1392),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1397),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1373),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1369),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1367),
.B(n_1359),
.Y(n_1434)
);

AOI31xp33_ASAP7_75t_L g1435 ( 
.A1(n_1378),
.A2(n_1328),
.A3(n_1337),
.B(n_1223),
.Y(n_1435)
);

NAND2x1p5_ASAP7_75t_L g1436 ( 
.A(n_1393),
.B(n_1347),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1401),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1414),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1435),
.B(n_1395),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1410),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1409),
.B(n_1280),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1403),
.A2(n_1398),
.B1(n_1381),
.B2(n_1387),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1410),
.Y(n_1443)
);

INVx1_ASAP7_75t_SL g1444 ( 
.A(n_1413),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1412),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1413),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1412),
.Y(n_1447)
);

AND3x2_ASAP7_75t_L g1448 ( 
.A(n_1437),
.B(n_1388),
.C(n_1386),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1418),
.B(n_1368),
.Y(n_1449)
);

INVx1_ASAP7_75t_SL g1450 ( 
.A(n_1418),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1420),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1415),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1411),
.A2(n_1387),
.B1(n_1381),
.B2(n_1388),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1420),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1432),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1415),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1416),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1431),
.B(n_1423),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1434),
.B(n_1249),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1405),
.B(n_1369),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1432),
.B(n_1381),
.Y(n_1461)
);

INVx1_ASAP7_75t_SL g1462 ( 
.A(n_1404),
.Y(n_1462)
);

AOI322xp5_ASAP7_75t_L g1463 ( 
.A1(n_1453),
.A2(n_1422),
.A3(n_1427),
.B1(n_1419),
.B2(n_1404),
.C1(n_1424),
.C2(n_1421),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1438),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1438),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1442),
.B(n_1436),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1440),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1459),
.B(n_1249),
.Y(n_1468)
);

INVx1_ASAP7_75t_SL g1469 ( 
.A(n_1449),
.Y(n_1469)
);

AO21x1_ASAP7_75t_L g1470 ( 
.A1(n_1446),
.A2(n_1436),
.B(n_1419),
.Y(n_1470)
);

OAI21xp33_ASAP7_75t_L g1471 ( 
.A1(n_1462),
.A2(n_1424),
.B(n_1421),
.Y(n_1471)
);

INVx1_ASAP7_75t_SL g1472 ( 
.A(n_1449),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1440),
.Y(n_1473)
);

AOI21xp33_ASAP7_75t_L g1474 ( 
.A1(n_1439),
.A2(n_1405),
.B(n_1433),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1450),
.B(n_1426),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1443),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1444),
.B(n_1426),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1443),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1448),
.B(n_1433),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1451),
.Y(n_1480)
);

INVx1_ASAP7_75t_SL g1481 ( 
.A(n_1460),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1480),
.B(n_1446),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1469),
.B(n_1458),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1480),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1472),
.B(n_1460),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1481),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1479),
.B(n_1454),
.Y(n_1487)
);

INVx1_ASAP7_75t_SL g1488 ( 
.A(n_1477),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1475),
.B(n_1454),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1464),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1471),
.B(n_1455),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1465),
.Y(n_1492)
);

NOR4xp25_ASAP7_75t_L g1493 ( 
.A(n_1487),
.B(n_1466),
.C(n_1474),
.D(n_1476),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_SL g1494 ( 
.A1(n_1482),
.A2(n_1466),
.B(n_1468),
.Y(n_1494)
);

OAI221xp5_ASAP7_75t_SL g1495 ( 
.A1(n_1491),
.A2(n_1463),
.B1(n_1485),
.B2(n_1488),
.C(n_1486),
.Y(n_1495)
);

NAND4xp25_ASAP7_75t_L g1496 ( 
.A(n_1483),
.B(n_1468),
.C(n_1441),
.D(n_1473),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1482),
.B(n_1455),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1489),
.B(n_1461),
.Y(n_1498)
);

OAI21xp33_ASAP7_75t_SL g1499 ( 
.A1(n_1484),
.A2(n_1467),
.B(n_1478),
.Y(n_1499)
);

OAI211xp5_ASAP7_75t_L g1500 ( 
.A1(n_1492),
.A2(n_1447),
.B(n_1445),
.C(n_1457),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1490),
.A2(n_1436),
.B1(n_1461),
.B2(n_1387),
.Y(n_1501)
);

AOI211xp5_ASAP7_75t_L g1502 ( 
.A1(n_1492),
.A2(n_1470),
.B(n_1461),
.C(n_1223),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1482),
.B(n_1445),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1497),
.Y(n_1504)
);

INVxp67_ASAP7_75t_SL g1505 ( 
.A(n_1503),
.Y(n_1505)
);

AOI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1493),
.A2(n_1387),
.B1(n_1379),
.B2(n_1452),
.Y(n_1506)
);

OAI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1494),
.A2(n_1456),
.B(n_1452),
.Y(n_1507)
);

AOI211xp5_ASAP7_75t_L g1508 ( 
.A1(n_1495),
.A2(n_1457),
.B(n_1456),
.C(n_1379),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1508),
.B(n_1498),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1506),
.B(n_1499),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1504),
.B(n_1368),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1507),
.Y(n_1512)
);

NOR2x1p5_ASAP7_75t_L g1513 ( 
.A(n_1505),
.B(n_1496),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1508),
.B(n_1502),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1512),
.A2(n_1500),
.B(n_1501),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1511),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1513),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1509),
.Y(n_1518)
);

AOI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1514),
.A2(n_1430),
.B1(n_1429),
.B2(n_1408),
.Y(n_1519)
);

OAI222xp33_ASAP7_75t_L g1520 ( 
.A1(n_1515),
.A2(n_1510),
.B1(n_1428),
.B2(n_1417),
.C1(n_1416),
.C2(n_1406),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1516),
.Y(n_1521)
);

NAND4xp75_ASAP7_75t_L g1522 ( 
.A(n_1517),
.B(n_1428),
.C(n_1417),
.D(n_1425),
.Y(n_1522)
);

AND3x2_ASAP7_75t_L g1523 ( 
.A(n_1521),
.B(n_1518),
.C(n_1242),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1523),
.B(n_1519),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1524),
.Y(n_1525)
);

AOI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1525),
.A2(n_1520),
.B(n_1522),
.Y(n_1526)
);

AOI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1526),
.A2(n_1407),
.B1(n_1375),
.B2(n_1377),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1527),
.Y(n_1528)
);

AOI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1527),
.A2(n_1375),
.B1(n_1377),
.B2(n_1399),
.Y(n_1529)
);

XNOR2x1_ASAP7_75t_L g1530 ( 
.A(n_1528),
.B(n_1210),
.Y(n_1530)
);

AOI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1529),
.A2(n_1394),
.B(n_1400),
.Y(n_1531)
);

OAI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1530),
.A2(n_1400),
.B(n_1399),
.Y(n_1532)
);

NOR4xp75_ASAP7_75t_L g1533 ( 
.A(n_1531),
.B(n_1391),
.C(n_1394),
.D(n_1402),
.Y(n_1533)
);

AOI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1532),
.A2(n_1391),
.B1(n_1396),
.B2(n_1351),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1533),
.Y(n_1535)
);

AOI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1535),
.A2(n_1396),
.B1(n_1351),
.B2(n_1350),
.Y(n_1536)
);

AOI211xp5_ASAP7_75t_L g1537 ( 
.A1(n_1536),
.A2(n_1534),
.B(n_1396),
.C(n_1351),
.Y(n_1537)
);


endmodule