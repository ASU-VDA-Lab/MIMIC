module fake_jpeg_19327_n_38 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_38);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_38;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_21),
.A2(n_22),
.B1(n_1),
.B2(n_2),
.Y(n_29)
);

INVx4_ASAP7_75t_SL g22 ( 
.A(n_19),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_23),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_SL g23 ( 
.A(n_16),
.B(n_0),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_6),
.C(n_12),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_24),
.B(n_7),
.Y(n_26)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_25),
.B(n_17),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_24),
.C(n_20),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_20),
.Y(n_32)
);

NAND2xp33_ASAP7_75t_R g31 ( 
.A(n_29),
.B(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_32),
.B1(n_27),
.B2(n_25),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_33),
.C(n_5),
.Y(n_37)
);

O2A1O1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_4),
.B(n_9),
.C(n_15),
.Y(n_38)
);


endmodule