module real_jpeg_10742_n_18 (n_17, n_8, n_0, n_2, n_10, n_338, n_9, n_12, n_6, n_337, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_338;
input n_9;
input n_12;
input n_6;
input n_337;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_1),
.A2(n_25),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_1),
.A2(n_30),
.B1(n_31),
.B2(n_38),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_1),
.A2(n_38),
.B1(n_67),
.B2(n_68),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_1),
.A2(n_38),
.B1(n_51),
.B2(n_52),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_2),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_2),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

AOI21xp33_ASAP7_75t_L g181 ( 
.A1(n_2),
.A2(n_12),
.B(n_31),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_3),
.A2(n_25),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_3),
.A2(n_34),
.B1(n_51),
.B2(n_52),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_3),
.A2(n_34),
.B1(n_67),
.B2(n_68),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g93 ( 
.A(n_4),
.Y(n_93)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_7),
.A2(n_30),
.B(n_49),
.C(n_50),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_7),
.B(n_30),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_7),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_9),
.A2(n_67),
.B1(n_68),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_9),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_9),
.A2(n_51),
.B1(n_52),
.B2(n_96),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_96),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_9),
.A2(n_25),
.B1(n_35),
.B2(n_96),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_10),
.A2(n_67),
.B1(n_68),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_10),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_10),
.A2(n_51),
.B1(n_52),
.B2(n_91),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_91),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_10),
.A2(n_25),
.B1(n_35),
.B2(n_91),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_12),
.A2(n_51),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_12),
.B(n_51),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_12),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_12),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_12),
.A2(n_30),
.B(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_12),
.B(n_30),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_12),
.B(n_32),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_12),
.A2(n_25),
.B1(n_35),
.B2(n_116),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_13),
.A2(n_51),
.B1(n_52),
.B2(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_13),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_13),
.A2(n_67),
.B1(n_68),
.B2(n_103),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_103),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_13),
.A2(n_25),
.B1(n_35),
.B2(n_103),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_14),
.A2(n_67),
.B1(n_68),
.B2(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_14),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_14),
.A2(n_51),
.B1(n_52),
.B2(n_132),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_132),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_14),
.A2(n_25),
.B1(n_35),
.B2(n_132),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_15),
.A2(n_25),
.B1(n_35),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_15),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_15),
.A2(n_59),
.B1(n_67),
.B2(n_68),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_15),
.A2(n_51),
.B1(n_52),
.B2(n_59),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_15),
.A2(n_30),
.B1(n_31),
.B2(n_59),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_16),
.A2(n_25),
.B1(n_35),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_16),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_16),
.A2(n_61),
.B1(n_67),
.B2(n_68),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_16),
.A2(n_51),
.B1(n_52),
.B2(n_61),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_16),
.A2(n_30),
.B1(n_31),
.B2(n_61),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_17),
.A2(n_67),
.B1(n_68),
.B2(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_17),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_17),
.A2(n_51),
.B1(n_52),
.B2(n_151),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_17),
.A2(n_30),
.B1(n_31),
.B2(n_151),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_17),
.A2(n_25),
.B1(n_35),
.B2(n_151),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_41),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_36),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_32),
.B(n_33),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_23),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_23),
.A2(n_32),
.B1(n_37),
.B2(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_23),
.A2(n_32),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_24),
.A2(n_29),
.B1(n_58),
.B2(n_60),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_24),
.A2(n_29),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_24),
.A2(n_29),
.B1(n_214),
.B2(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_24),
.A2(n_29),
.B1(n_239),
.B2(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_24),
.A2(n_29),
.B1(n_257),
.B2(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_24),
.A2(n_29),
.B1(n_58),
.B2(n_283),
.Y(n_305)
);

A2O1A1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_27),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_25),
.A2(n_27),
.B(n_116),
.C(n_181),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_29),
.Y(n_32)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_36),
.B(n_43),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_78),
.B(n_335),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_71),
.C(n_73),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_44),
.A2(n_45),
.B1(n_330),
.B2(n_332),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_56),
.C(n_62),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_46),
.A2(n_47),
.B1(n_62),
.B2(n_310),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_50),
.B1(n_54),
.B2(n_55),
.Y(n_47)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_48),
.A2(n_50),
.B1(n_140),
.B2(n_142),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_48),
.A2(n_50),
.B1(n_142),
.B2(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_48),
.A2(n_50),
.B1(n_159),
.B2(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_48),
.A2(n_50),
.B1(n_199),
.B2(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_48),
.A2(n_50),
.B1(n_210),
.B2(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_48),
.A2(n_50),
.B1(n_236),
.B2(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_48),
.A2(n_50),
.B1(n_54),
.B2(n_309),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_49),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_50),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_50),
.B(n_116),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_SL g63 ( 
.A1(n_51),
.A2(n_64),
.B(n_65),
.C(n_66),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_64),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_51),
.B(n_53),
.Y(n_146)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_52),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_55),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_56),
.A2(n_57),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_62),
.A2(n_308),
.B1(n_310),
.B2(n_311),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_62),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_66),
.B(n_70),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_63),
.A2(n_66),
.B1(n_100),
.B2(n_102),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_63),
.A2(n_66),
.B1(n_102),
.B2(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_63),
.A2(n_66),
.B1(n_129),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_63),
.A2(n_66),
.B1(n_138),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_63),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_63),
.A2(n_66),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_63),
.A2(n_66),
.B1(n_222),
.B2(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_63),
.A2(n_66),
.B1(n_231),
.B2(n_263),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_64),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_64),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_66),
.B(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_66),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_67),
.B(n_69),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_67),
.B(n_120),
.Y(n_119)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_68),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_70),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_71),
.A2(n_73),
.B1(n_74),
.B2(n_331),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_71),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_76),
.B(n_77),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_75),
.A2(n_76),
.B1(n_275),
.B2(n_276),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_328),
.B(n_334),
.Y(n_78)
);

OAI321xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_301),
.A3(n_321),
.B1(n_326),
.B2(n_327),
.C(n_337),
.Y(n_79)
);

AOI321xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_247),
.A3(n_289),
.B1(n_295),
.B2(n_300),
.C(n_338),
.Y(n_80)
);

NOR3xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_204),
.C(n_243),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_174),
.B(n_203),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_153),
.B(n_173),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_134),
.B(n_152),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_123),
.B(n_133),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_109),
.B(n_122),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_97),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_88),
.B(n_97),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_90),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_92),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_92),
.A2(n_93),
.B1(n_150),
.B2(n_164),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_93),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_95),
.A2(n_113),
.B1(n_114),
.B2(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_104),
.B2(n_108),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_98),
.B(n_108),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_101),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_104),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_117),
.B(n_121),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_115),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_113),
.A2(n_114),
.B1(n_131),
.B2(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_113),
.A2(n_114),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_113),
.A2(n_114),
.B1(n_185),
.B2(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_113),
.A2(n_114),
.B1(n_219),
.B2(n_229),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_113),
.A2(n_114),
.B(n_229),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_116),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_124),
.B(n_125),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_130),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_128),
.C(n_130),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_135),
.B(n_136),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_136),
.Y(n_154)
);

FAx1_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_139),
.CI(n_143),
.CON(n_136),
.SN(n_136)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_141),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_148),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_148),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_154),
.B(n_155),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_166),
.B2(n_167),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_169),
.C(n_171),
.Y(n_175)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_160),
.B1(n_161),
.B2(n_165),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_158),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_163),
.C(n_165),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_164),
.Y(n_184)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_171),
.B2(n_172),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_168),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_169),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_170),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_175),
.B(n_176),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_189),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_178),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_178),
.B(n_188),
.C(n_189),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_182),
.B2(n_183),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_183),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_186),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_200),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_197),
.B2(n_198),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_197),
.C(n_200),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_194),
.A2(n_196),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_195),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_202),
.Y(n_213)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

AOI21xp33_ASAP7_75t_L g296 ( 
.A1(n_205),
.A2(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_224),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_206),
.B(n_224),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_217),
.C(n_223),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_207),
.B(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_216),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_211),
.B1(n_212),
.B2(n_215),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_209),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_SL g241 ( 
.A(n_211),
.B(n_215),
.C(n_216),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_223),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_220),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_241),
.B2(n_242),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_232),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_227),
.B(n_232),
.C(n_242),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_230),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_237),
.C(n_240),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_237),
.B1(n_238),
.B2(n_240),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_235),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_241),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_244),
.B(n_245),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_266),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_248),
.B(n_266),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_259),
.C(n_265),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_249),
.A2(n_250),
.B1(n_259),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_251),
.B(n_255),
.C(n_258),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_255),
.B1(n_256),
.B2(n_258),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_253),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_254),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_259),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_264),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_260),
.A2(n_261),
.B1(n_282),
.B2(n_284),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_260),
.A2(n_282),
.B(n_285),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_262),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_262),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_263),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_293),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_287),
.B2(n_288),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_278),
.B2(n_279),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_269),
.B(n_279),
.C(n_288),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_274),
.B(n_277),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_274),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_276),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_277),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_277),
.A2(n_303),
.B1(n_312),
.B2(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_285),
.B2(n_286),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_282),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_287),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_290),
.A2(n_296),
.B(n_299),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_291),
.B(n_292),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_314),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_302),
.B(n_314),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_312),
.C(n_313),
.Y(n_302)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_303),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_304),
.A2(n_305),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_305),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_310),
.C(n_311),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_305),
.B(n_316),
.C(n_320),
.Y(n_333)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_308),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_324),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_320),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_322),
.B(n_323),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_333),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_333),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_330),
.Y(n_332)
);


endmodule