module real_jpeg_31110_n_20 (n_17, n_8, n_0, n_722, n_2, n_10, n_9, n_12, n_723, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_722;
input n_2;
input n_10;
input n_9;
input n_12;
input n_723;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_715;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_696;
wire n_657;
wire n_656;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_719;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_678;
wire n_30;
wire n_332;
wire n_149;
wire n_620;
wire n_328;
wire n_366;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_682;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_611;
wire n_221;
wire n_393;
wire n_489;
wire n_634;
wire n_104;
wire n_153;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_704;
wire n_576;
wire n_139;
wire n_33;
wire n_673;
wire n_631;
wire n_175;
wire n_718;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_707;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_710;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_703;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_411;
wire n_382;
wire n_314;
wire n_278;
wire n_689;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_697;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_716;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_712;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_714;
wire n_89;
wire n_407;
wire n_693;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_692;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_638;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_711;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_688;
wire n_342;
wire n_120;
wire n_586;
wire n_155;
wire n_405;
wire n_412;
wire n_572;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_698;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_546;
wire n_285;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_686;
wire n_391;
wire n_427;
wire n_401;
wire n_699;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_720;
wire n_600;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_708;
wire n_667;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_691;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_701;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_695;
wire n_138;
wire n_662;
wire n_217;
wire n_709;
wire n_53;
wire n_717;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_702;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_706;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_700;
wire n_94;
wire n_645;
wire n_687;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_588;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_705;
wire n_530;
wire n_361;
wire n_694;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_690;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_713;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g227 ( 
.A(n_0),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_0),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g301 ( 
.A(n_0),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_0),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_1),
.A2(n_201),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_1),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_1),
.A2(n_308),
.B1(n_369),
.B2(n_372),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_1),
.A2(n_308),
.B1(n_547),
.B2(n_550),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_1),
.A2(n_308),
.B1(n_611),
.B2(n_612),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

OAI22x1_ASAP7_75t_SL g196 ( 
.A1(n_3),
.A2(n_197),
.B1(n_198),
.B2(n_201),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_3),
.Y(n_197)
);

AOI22x1_ASAP7_75t_SL g315 ( 
.A1(n_3),
.A2(n_197),
.B1(n_316),
.B2(n_320),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_3),
.A2(n_197),
.B1(n_357),
.B2(n_361),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_3),
.A2(n_197),
.B1(n_411),
.B2(n_416),
.Y(n_410)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_4),
.A2(n_135),
.B1(n_138),
.B2(n_140),
.Y(n_134)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_4),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_4),
.A2(n_140),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_4),
.A2(n_140),
.B1(n_254),
.B2(n_256),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_4),
.A2(n_140),
.B1(n_448),
.B2(n_452),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_L g390 ( 
.A1(n_5),
.A2(n_130),
.B1(n_199),
.B2(n_391),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_5),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_5),
.A2(n_391),
.B1(n_396),
.B2(n_398),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_5),
.A2(n_391),
.B1(n_586),
.B2(n_588),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_SL g633 ( 
.A1(n_5),
.A2(n_391),
.B1(n_593),
.B2(n_634),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_6),
.A2(n_63),
.B1(n_67),
.B2(n_72),
.Y(n_62)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_6),
.Y(n_72)
);

AO22x1_ASAP7_75t_L g119 ( 
.A1(n_6),
.A2(n_72),
.B1(n_120),
.B2(n_122),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_6),
.A2(n_72),
.B1(n_174),
.B2(n_177),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_6),
.A2(n_72),
.B1(n_236),
.B2(n_239),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_7),
.A2(n_382),
.B(n_386),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_7),
.B(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_7),
.Y(n_422)
);

OAI32xp33_ASAP7_75t_L g553 ( 
.A1(n_7),
.A2(n_426),
.A3(n_554),
.B1(n_557),
.B2(n_558),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_7),
.B(n_172),
.Y(n_618)
);

OAI22xp33_ASAP7_75t_L g648 ( 
.A1(n_7),
.A2(n_228),
.B1(n_633),
.B2(n_649),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_7),
.A2(n_422),
.B1(n_674),
.B2(n_678),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_8),
.A2(n_51),
.B1(n_57),
.B2(n_60),
.Y(n_50)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_8),
.A2(n_60),
.B1(n_163),
.B2(n_167),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_8),
.A2(n_259),
.B(n_261),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_8),
.B(n_262),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_8),
.A2(n_60),
.B1(n_239),
.B2(n_303),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_10),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_11),
.Y(n_108)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_11),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_11),
.Y(n_242)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_11),
.Y(n_451)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_12),
.Y(n_713)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_13),
.Y(n_94)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_13),
.Y(n_102)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_13),
.Y(n_598)
);

OAI22xp33_ASAP7_75t_L g129 ( 
.A1(n_14),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_14),
.Y(n_131)
);

OAI22x1_ASAP7_75t_SL g273 ( 
.A1(n_14),
.A2(n_131),
.B1(n_274),
.B2(n_280),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_14),
.A2(n_131),
.B1(n_290),
.B2(n_292),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_14),
.A2(n_131),
.B1(n_404),
.B2(n_405),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_15),
.A2(n_246),
.B1(n_249),
.B2(n_250),
.Y(n_245)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_15),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_15),
.A2(n_249),
.B1(n_351),
.B2(n_354),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_15),
.A2(n_249),
.B1(n_472),
.B2(n_474),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_15),
.A2(n_249),
.B1(n_472),
.B2(n_474),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_15),
.A2(n_249),
.B1(n_562),
.B2(n_564),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g374 ( 
.A1(n_16),
.A2(n_372),
.B1(n_375),
.B2(n_378),
.Y(n_374)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_16),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_16),
.A2(n_64),
.B1(n_378),
.B2(n_481),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_16),
.A2(n_378),
.B1(n_621),
.B2(n_624),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_SL g637 ( 
.A1(n_16),
.A2(n_378),
.B1(n_638),
.B2(n_641),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_17),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_17),
.B(n_712),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_18),
.Y(n_97)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_18),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_18),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_18),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_19),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_19),
.Y(n_176)
);

OAI32xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_78),
.A3(n_712),
.B1(n_716),
.B2(n_719),
.Y(n_20)
);

AOI21xp33_ASAP7_75t_SL g719 ( 
.A1(n_21),
.A2(n_718),
.B(n_720),
.Y(n_719)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_75),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_74),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_23),
.Y(n_76)
);

NAND4xp25_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_49),
.C(n_61),
.D(n_73),
.Y(n_23)
);

NAND2xp33_ASAP7_75t_R g24 ( 
.A(n_25),
.B(n_48),
.Y(n_24)
);

NAND2xp33_ASAP7_75t_L g61 ( 
.A(n_25),
.B(n_62),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_25),
.A2(n_48),
.B(n_62),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_25),
.A2(n_48),
.B1(n_128),
.B2(n_134),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_25),
.A2(n_48),
.B1(n_50),
.B2(n_134),
.Y(n_187)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_26),
.A2(n_129),
.B1(n_196),
.B2(n_204),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_26),
.A2(n_204),
.B1(n_479),
.B2(n_484),
.Y(n_478)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_27),
.A2(n_48),
.B1(n_381),
.B2(n_390),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_27),
.A2(n_48),
.B1(n_307),
.B2(n_480),
.Y(n_498)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_28),
.B(n_245),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_28),
.A2(n_204),
.B1(n_245),
.B2(n_306),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_39),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_32),
.Y(n_137)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_32),
.Y(n_311)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_33),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_33),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_33),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_34),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_35),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_36),
.Y(n_130)
);

INVxp67_ASAP7_75t_SL g139 ( 
.A(n_36),
.Y(n_139)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_43),
.B2(n_45),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_42),
.Y(n_170)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_42),
.Y(n_181)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_43),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_43),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_44),
.Y(n_166)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_44),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_44),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_44),
.Y(n_440)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp33_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_48),
.Y(n_204)
);

NOR2x1_ASAP7_75t_L g421 ( 
.A(n_48),
.B(n_422),
.Y(n_421)
);

NAND2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_62),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_59),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g250 ( 
.A(n_65),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g133 ( 
.A(n_68),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_69),
.Y(n_200)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_70),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_71),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_74),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_76),
.B(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_76),
.B(n_214),
.Y(n_711)
);

AOI211xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_339),
.B(n_701),
.C(n_711),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI221xp5_ASAP7_75t_L g716 ( 
.A1(n_80),
.A2(n_340),
.B1(n_717),
.B2(n_718),
.C(n_723),
.Y(n_716)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AND3x1_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_213),
.C(n_215),
.Y(n_81)
);

INVxp33_ASAP7_75t_SL g710 ( 
.A(n_82),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_188),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_83),
.B(n_188),
.Y(n_706)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_182),
.B2(n_183),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_85),
.B(n_184),
.C(n_187),
.Y(n_214)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_127),
.C(n_141),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_87),
.A2(n_142),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_87),
.A2(n_192),
.B1(n_207),
.B2(n_331),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_116),
.B(n_119),
.Y(n_87)
);

OA21x2_ASAP7_75t_L g192 ( 
.A1(n_88),
.A2(n_116),
.B(n_119),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_88),
.B(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_89),
.A2(n_117),
.B1(n_253),
.B2(n_258),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_89),
.Y(n_270)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_89),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_89),
.A2(n_289),
.B1(n_356),
.B2(n_365),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_89),
.A2(n_365),
.B1(n_620),
.B2(n_626),
.Y(n_619)
);

AO21x2_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_98),
.B(n_106),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g625 ( 
.A(n_96),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_97),
.Y(n_160)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_97),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_97),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_97),
.Y(n_556)
);

INVxp33_ASAP7_75t_L g604 ( 
.A(n_98),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g363 ( 
.A(n_103),
.Y(n_363)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_104),
.Y(n_255)
);

INVx5_ASAP7_75t_L g623 ( 
.A(n_104),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g294 ( 
.A(n_105),
.Y(n_294)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_109),
.B1(n_111),
.B2(n_114),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_108),
.Y(n_408)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_108),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_108),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_108),
.Y(n_655)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_113),
.Y(n_233)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_113),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_113),
.Y(n_419)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_116),
.A2(n_119),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_116),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_116),
.B(n_296),
.Y(n_505)
);

AO22x1_ASAP7_75t_L g545 ( 
.A1(n_116),
.A2(n_349),
.B1(n_350),
.B2(n_546),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_116),
.A2(n_270),
.B1(n_546),
.B2(n_671),
.Y(n_670)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g646 ( 
.A(n_117),
.B(n_422),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_118),
.Y(n_366)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_125),
.Y(n_257)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_126),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_126),
.Y(n_584)
);

XOR2x2_ASAP7_75t_L g189 ( 
.A(n_127),
.B(n_190),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_142),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_162),
.B1(n_171),
.B2(n_173),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_143),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_143),
.A2(n_162),
.B1(n_171),
.B2(n_208),
.Y(n_207)
);

OA22x2_ASAP7_75t_L g367 ( 
.A1(n_143),
.A2(n_171),
.B1(n_368),
.B2(n_374),
.Y(n_367)
);

OAI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_143),
.A2(n_171),
.B1(n_374),
.B2(n_395),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_143),
.A2(n_171),
.B1(n_368),
.B2(n_471),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_143),
.A2(n_171),
.B1(n_315),
.B2(n_500),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g672 ( 
.A1(n_143),
.A2(n_171),
.B1(n_395),
.B2(n_673),
.Y(n_672)
);

AO21x2_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_149),
.B(n_155),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_149),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_150),
.Y(n_320)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_L g400 ( 
.A(n_151),
.Y(n_400)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_151),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_152),
.Y(n_283)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_158),
.B1(n_160),
.B2(n_161),
.Y(n_155)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_156),
.Y(n_589)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_160),
.Y(n_260)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_166),
.Y(n_679)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_SL g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_172),
.A2(n_185),
.B(n_186),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_172),
.A2(n_185),
.B1(n_209),
.B2(n_273),
.Y(n_272)
);

AOI22x1_ASAP7_75t_L g313 ( 
.A1(n_172),
.A2(n_185),
.B1(n_273),
.B2(n_314),
.Y(n_313)
);

INVxp33_ASAP7_75t_L g186 ( 
.A(n_173),
.Y(n_186)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_174),
.Y(n_210)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_176),
.Y(n_212)
);

INVx8_ASAP7_75t_L g371 ( 
.A(n_176),
.Y(n_371)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_181),
.Y(n_677)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.Y(n_183)
);

MAJx2_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_193),
.C(n_205),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_189),
.B(n_336),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_193),
.C(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_193),
.Y(n_336)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_195),
.B(n_330),
.Y(n_329)
);

AOI21x1_ASAP7_75t_L g243 ( 
.A1(n_196),
.A2(n_204),
.B(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx11_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_205),
.B(n_335),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_207),
.Y(n_331)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g709 ( 
.A(n_213),
.Y(n_709)
);

NOR2x1_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_332),
.Y(n_215)
);

NOR2xp67_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_321),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_217),
.B(n_321),
.Y(n_708)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_267),
.C(n_285),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_219),
.A2(n_267),
.B1(n_268),
.B2(n_528),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_219),
.Y(n_528)
);

OAI22x1_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_251),
.B2(n_266),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2x1_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_243),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_222),
.A2(n_323),
.B1(n_325),
.B2(n_722),
.Y(n_322)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_222),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_234),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_228),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_227),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_228),
.A2(n_235),
.B1(n_299),
.B2(n_302),
.Y(n_298)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_228),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_228),
.A2(n_302),
.B1(n_444),
.B2(n_447),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_228),
.A2(n_607),
.B1(n_609),
.B2(n_610),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_SL g632 ( 
.A1(n_228),
.A2(n_633),
.B1(n_637),
.B2(n_644),
.Y(n_632)
);

OR2x6_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

BUFx2_ASAP7_75t_R g409 ( 
.A(n_229),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_229),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_230),
.Y(n_645)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_230),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_239),
.Y(n_611)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_241),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx6_ASAP7_75t_L g415 ( 
.A(n_242),
.Y(n_415)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_242),
.Y(n_594)
);

INVxp33_ASAP7_75t_L g326 ( 
.A(n_243),
.Y(n_326)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_248),
.Y(n_432)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_251),
.Y(n_324)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_252),
.Y(n_518)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_253),
.Y(n_296)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_254),
.Y(n_550)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_257),
.Y(n_291)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx6f_ASAP7_75t_SL g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_264),
.Y(n_587)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

OAI21xp33_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_272),
.B(n_284),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_272),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_270),
.A2(n_364),
.B1(n_577),
.B2(n_585),
.Y(n_576)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVxp67_ASAP7_75t_SL g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_283),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_284),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_285),
.B(n_527),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_304),
.C(n_312),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_286),
.B(n_522),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_295),
.B(n_297),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_287),
.B(n_505),
.Y(n_504)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_289),
.Y(n_288)
);

BUFx4f_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_294),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_297),
.B(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_299),
.B(n_422),
.Y(n_651)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx8_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx8_ASAP7_75t_L g608 ( 
.A(n_301),
.Y(n_608)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_303),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_305),
.B(n_313),
.Y(n_522)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVxp33_ASAP7_75t_SL g312 ( 
.A(n_313),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_327),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_328),
.C(n_338),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g325 ( 
.A(n_326),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_329),
.Y(n_338)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_333),
.B(n_708),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_337),
.Y(n_333)
);

NOR2xp67_ASAP7_75t_SL g705 ( 
.A(n_334),
.B(n_337),
.Y(n_705)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

AO21x2_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_529),
.B(n_694),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_508),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_488),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_462),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_345),
.B(n_462),
.Y(n_697)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_392),
.C(n_423),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g532 ( 
.A(n_346),
.B(n_533),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_379),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_367),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_348),
.B(n_367),
.C(n_379),
.Y(n_467)
);

AOI22x1_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_350),
.B1(n_355),
.B2(n_364),
.Y(n_348)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_353),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx5_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_361),
.B(n_422),
.Y(n_558)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx5_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx5_ASAP7_75t_L g377 ( 
.A(n_371),
.Y(n_377)
);

INVx5_ASAP7_75t_L g397 ( 
.A(n_371),
.Y(n_397)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_371),
.Y(n_427)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx2_ASAP7_75t_SL g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g441 ( 
.A(n_386),
.Y(n_441)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_390),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_393),
.B(n_423),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_401),
.C(n_421),
.Y(n_393)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_394),
.Y(n_537)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_401),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g543 ( 
.A1(n_401),
.A2(n_538),
.B(n_539),
.Y(n_543)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g540 ( 
.A(n_402),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_403),
.A2(n_409),
.B1(n_410),
.B2(n_420),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_403),
.A2(n_420),
.B1(n_443),
.B2(n_446),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx4_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_410),
.A2(n_420),
.B1(n_561),
.B2(n_568),
.Y(n_560)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_415),
.Y(n_563)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_415),
.Y(n_603)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_415),
.Y(n_636)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_419),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_SL g658 ( 
.A1(n_420),
.A2(n_659),
.B1(n_660),
.B2(n_661),
.Y(n_658)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_421),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_421),
.B(n_542),
.Y(n_541)
);

OAI21xp33_ASAP7_75t_SL g577 ( 
.A1(n_422),
.A2(n_578),
.B(n_581),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_422),
.B(n_582),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_424),
.A2(n_442),
.B1(n_456),
.B2(n_461),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_424),
.B(n_461),
.Y(n_487)
);

OAI32xp33_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_428),
.A3(n_431),
.B1(n_433),
.B2(n_441),
.Y(n_424)
);

OAI32xp33_ASAP7_75t_L g457 ( 
.A1(n_425),
.A2(n_428),
.A3(n_433),
.B1(n_441),
.B2(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx3_ASAP7_75t_SL g426 ( 
.A(n_427),
.Y(n_426)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_437),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_442),
.Y(n_461)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx2_ASAP7_75t_SL g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_451),
.Y(n_616)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_455),
.Y(n_567)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_468),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_467),
.Y(n_463)
);

INVxp67_ASAP7_75t_SL g490 ( 
.A(n_464),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_466),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_465),
.B(n_466),
.Y(n_495)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_467),
.Y(n_491)
);

MAJx2_ASAP7_75t_L g489 ( 
.A(n_468),
.B(n_490),
.C(n_491),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_487),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_470),
.A2(n_478),
.B1(n_485),
.B2(n_486),
.Y(n_469)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_470),
.Y(n_485)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_478),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_478),
.B(n_485),
.C(n_487),
.Y(n_507)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx8_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

NAND2xp67_ASAP7_75t_SL g488 ( 
.A(n_489),
.B(n_492),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g696 ( 
.A(n_489),
.B(n_492),
.C(n_697),
.Y(n_696)
);

XOR2x2_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_507),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_494),
.A2(n_502),
.B1(n_503),
.B2(n_506),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_494),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_494),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_496),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_495),
.B(n_497),
.C(n_514),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_497),
.A2(n_498),
.B1(n_499),
.B2(n_501),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_499),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_501),
.Y(n_514)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_503),
.B(n_507),
.C(n_511),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_SL g694 ( 
.A1(n_508),
.A2(n_695),
.B(n_698),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_523),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_510),
.B(n_512),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_510),
.B(n_512),
.Y(n_699)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_515),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_513),
.B(n_516),
.C(n_525),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_521),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_517),
.A2(n_518),
.B1(n_519),
.B2(n_520),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_519),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_521),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_523),
.A2(n_699),
.B(n_700),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_526),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_524),
.B(n_526),
.Y(n_700)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

AOI21x1_ASAP7_75t_L g530 ( 
.A1(n_531),
.A2(n_570),
.B(n_693),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_532),
.B(n_534),
.Y(n_531)
);

NOR2xp67_ASAP7_75t_SL g693 ( 
.A(n_532),
.B(n_534),
.Y(n_693)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_535),
.B(n_545),
.C(n_551),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g687 ( 
.A(n_535),
.B(n_688),
.Y(n_687)
);

AOI22x1_ASAP7_75t_L g535 ( 
.A1(n_536),
.A2(n_541),
.B1(n_543),
.B2(n_544),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_537),
.B(n_538),
.Y(n_536)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_537),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_540),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_545),
.A2(n_689),
.B(n_690),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_SL g690 ( 
.A(n_545),
.B(n_552),
.Y(n_690)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_551),
.Y(n_689)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_553),
.B(n_559),
.Y(n_552)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_553),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_553),
.B(n_560),
.Y(n_684)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_559),
.Y(n_683)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_561),
.Y(n_609)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

BUFx4f_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

OAI21x1_ASAP7_75t_L g570 ( 
.A1(n_571),
.A2(n_686),
.B(n_692),
.Y(n_570)
);

AOI21x1_ASAP7_75t_L g571 ( 
.A1(n_572),
.A2(n_665),
.B(n_685),
.Y(n_571)
);

OAI21x1_ASAP7_75t_SL g572 ( 
.A1(n_573),
.A2(n_629),
.B(n_664),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_574),
.B(n_605),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_574),
.B(n_605),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_575),
.B(n_590),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_575),
.A2(n_576),
.B1(n_590),
.B2(n_591),
.Y(n_662)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g599 ( 
.A(n_581),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_585),
.Y(n_626)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_592),
.A2(n_599),
.B1(n_600),
.B2(n_604),
.Y(n_591)
);

NAND2xp33_ASAP7_75t_SL g592 ( 
.A(n_593),
.B(n_595),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_594),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_601),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_602),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g605 ( 
.A(n_606),
.B(n_617),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g666 ( 
.A(n_606),
.B(n_619),
.C(n_627),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_608),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g660 ( 
.A(n_610),
.Y(n_660)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_613),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_614),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_615),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_616),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_618),
.A2(n_619),
.B1(n_627),
.B2(n_628),
.Y(n_617)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_618),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_619),
.Y(n_628)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_620),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_622),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_623),
.Y(n_622)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_625),
.Y(n_624)
);

AOI21x1_ASAP7_75t_SL g629 ( 
.A1(n_630),
.A2(n_657),
.B(n_663),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_L g630 ( 
.A1(n_631),
.A2(n_647),
.B(n_656),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_632),
.B(n_646),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_632),
.B(n_646),
.Y(n_656)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_635),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_636),
.Y(n_635)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_637),
.Y(n_659)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_639),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_640),
.Y(n_639)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_642),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_643),
.Y(n_642)
);

INVx8_ASAP7_75t_L g644 ( 
.A(n_645),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_648),
.B(n_650),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_SL g650 ( 
.A(n_651),
.B(n_652),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_653),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_654),
.Y(n_653)
);

BUFx2_ASAP7_75t_SL g654 ( 
.A(n_655),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_658),
.B(n_662),
.Y(n_657)
);

NOR2xp67_ASAP7_75t_L g663 ( 
.A(n_658),
.B(n_662),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_666),
.B(n_667),
.Y(n_665)
);

NOR2x1_ASAP7_75t_L g685 ( 
.A(n_666),
.B(n_667),
.Y(n_685)
);

XNOR2x1_ASAP7_75t_L g667 ( 
.A(n_668),
.B(n_681),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_669),
.A2(n_670),
.B1(n_672),
.B2(n_680),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_670),
.Y(n_669)
);

MAJIxp5_ASAP7_75t_L g691 ( 
.A(n_670),
.B(n_680),
.C(n_681),
.Y(n_691)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_672),
.Y(n_680)
);

INVx1_ASAP7_75t_SL g674 ( 
.A(n_675),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_676),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_677),
.Y(n_676)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_679),
.Y(n_678)
);

AOI21x1_ASAP7_75t_L g681 ( 
.A1(n_682),
.A2(n_683),
.B(n_684),
.Y(n_681)
);

NOR2xp67_ASAP7_75t_SL g686 ( 
.A(n_687),
.B(n_691),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_687),
.B(n_691),
.Y(n_692)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_696),
.Y(n_695)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_701),
.Y(n_720)
);

INVxp67_ASAP7_75t_SL g701 ( 
.A(n_702),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_703),
.Y(n_702)
);

AOI211xp5_ASAP7_75t_L g703 ( 
.A1(n_704),
.A2(n_707),
.B(n_709),
.C(n_710),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_705),
.B(n_706),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_711),
.B(n_712),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_713),
.B(n_714),
.Y(n_712)
);

CKINVDCx11_ASAP7_75t_R g714 ( 
.A(n_715),
.Y(n_714)
);


endmodule