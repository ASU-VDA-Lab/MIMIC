module fake_aes_7946_n_266 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_266);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_266;
wire n_117;
wire n_219;
wire n_133;
wire n_149;
wire n_220;
wire n_81;
wire n_214;
wire n_221;
wire n_204;
wire n_249;
wire n_185;
wire n_203;
wire n_88;
wire n_244;
wire n_102;
wire n_141;
wire n_119;
wire n_115;
wire n_97;
wire n_80;
wire n_167;
wire n_107;
wire n_158;
wire n_114;
wire n_121;
wire n_171;
wire n_94;
wire n_196;
wire n_125;
wire n_192;
wire n_240;
wire n_254;
wire n_161;
wire n_262;
wire n_177;
wire n_130;
wire n_189;
wire n_103;
wire n_239;
wire n_87;
wire n_137;
wire n_180;
wire n_104;
wire n_160;
wire n_98;
wire n_74;
wire n_206;
wire n_154;
wire n_195;
wire n_165;
wire n_146;
wire n_85;
wire n_250;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_215;
wire n_91;
wire n_108;
wire n_116;
wire n_155;
wire n_209;
wire n_217;
wire n_139;
wire n_230;
wire n_229;
wire n_198;
wire n_169;
wire n_193;
wire n_252;
wire n_152;
wire n_113;
wire n_241;
wire n_95;
wire n_124;
wire n_156;
wire n_238;
wire n_128;
wire n_129;
wire n_120;
wire n_90;
wire n_135;
wire n_188;
wire n_78;
wire n_247;
wire n_197;
wire n_201;
wire n_242;
wire n_260;
wire n_127;
wire n_170;
wire n_111;
wire n_157;
wire n_79;
wire n_210;
wire n_202;
wire n_142;
wire n_184;
wire n_245;
wire n_265;
wire n_191;
wire n_264;
wire n_232;
wire n_208;
wire n_200;
wire n_211;
wire n_122;
wire n_187;
wire n_138;
wire n_126;
wire n_178;
wire n_118;
wire n_258;
wire n_253;
wire n_179;
wire n_84;
wire n_131;
wire n_112;
wire n_205;
wire n_86;
wire n_143;
wire n_213;
wire n_235;
wire n_243;
wire n_182;
wire n_263;
wire n_166;
wire n_162;
wire n_186;
wire n_75;
wire n_163;
wire n_226;
wire n_105;
wire n_159;
wire n_174;
wire n_227;
wire n_248;
wire n_231;
wire n_136;
wire n_89;
wire n_76;
wire n_176;
wire n_144;
wire n_183;
wire n_256;
wire n_77;
wire n_216;
wire n_147;
wire n_199;
wire n_148;
wire n_123;
wire n_83;
wire n_172;
wire n_100;
wire n_212;
wire n_228;
wire n_92;
wire n_223;
wire n_251;
wire n_236;
wire n_150;
wire n_218;
wire n_168;
wire n_194;
wire n_110;
wire n_261;
wire n_134;
wire n_222;
wire n_234;
wire n_164;
wire n_233;
wire n_82;
wire n_106;
wire n_175;
wire n_173;
wire n_190;
wire n_145;
wire n_246;
wire n_153;
wire n_259;
wire n_132;
wire n_109;
wire n_99;
wire n_93;
wire n_151;
wire n_140;
wire n_207;
wire n_257;
wire n_224;
wire n_96;
wire n_225;
INVx1_ASAP7_75t_L g74 ( .A(n_57), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_35), .Y(n_75) );
INVxp33_ASAP7_75t_L g76 ( .A(n_43), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_25), .Y(n_77) );
CKINVDCx14_ASAP7_75t_R g78 ( .A(n_52), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_21), .Y(n_79) );
INVx3_ASAP7_75t_L g80 ( .A(n_71), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_18), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_55), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_19), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_20), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_29), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_39), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_62), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_10), .Y(n_88) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_56), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_70), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_27), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_42), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_65), .Y(n_93) );
BUFx2_ASAP7_75t_L g94 ( .A(n_38), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_32), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_0), .Y(n_96) );
INVxp67_ASAP7_75t_SL g97 ( .A(n_66), .Y(n_97) );
INVxp33_ASAP7_75t_L g98 ( .A(n_64), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_44), .Y(n_99) );
INVxp67_ASAP7_75t_L g100 ( .A(n_47), .Y(n_100) );
BUFx6f_ASAP7_75t_L g101 ( .A(n_13), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_54), .Y(n_102) );
BUFx6f_ASAP7_75t_L g103 ( .A(n_59), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_34), .Y(n_104) );
INVxp67_ASAP7_75t_SL g105 ( .A(n_37), .Y(n_105) );
BUFx5_ASAP7_75t_L g106 ( .A(n_9), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_48), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_51), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_53), .Y(n_109) );
INVx3_ASAP7_75t_L g110 ( .A(n_2), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_40), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_15), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_11), .Y(n_113) );
AOI22x1_ASAP7_75t_L g114 ( .A1(n_82), .A2(n_28), .B1(n_73), .B2(n_72), .Y(n_114) );
AND2x4_ASAP7_75t_L g115 ( .A(n_110), .B(n_0), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_106), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_106), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_89), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_89), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_80), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_106), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_89), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_89), .Y(n_123) );
OAI21x1_ASAP7_75t_L g124 ( .A1(n_82), .A2(n_17), .B(n_16), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_103), .Y(n_125) );
BUFx3_ASAP7_75t_L g126 ( .A(n_94), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_103), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_106), .Y(n_128) );
BUFx2_ASAP7_75t_L g129 ( .A(n_110), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_87), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_103), .Y(n_131) );
AND2x4_ASAP7_75t_L g132 ( .A(n_87), .B(n_1), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_101), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_126), .B(n_76), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_118), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_116), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_116), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_117), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_115), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_121), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_129), .B(n_76), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_118), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_118), .Y(n_143) );
NAND3xp33_ASAP7_75t_L g144 ( .A(n_128), .B(n_75), .C(n_74), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_118), .Y(n_145) );
BUFx3_ASAP7_75t_L g146 ( .A(n_115), .Y(n_146) );
NAND2xp33_ASAP7_75t_SL g147 ( .A(n_115), .B(n_84), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_132), .B(n_104), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_120), .B(n_98), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_118), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_118), .Y(n_151) );
AND2x6_ASAP7_75t_L g152 ( .A(n_132), .B(n_77), .Y(n_152) );
AND2x6_ASAP7_75t_L g153 ( .A(n_132), .B(n_79), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_130), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_134), .B(n_109), .Y(n_155) );
BUFx3_ASAP7_75t_L g156 ( .A(n_152), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_141), .B(n_78), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_154), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_148), .B(n_90), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_146), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_139), .Y(n_161) );
A2O1A1Ixp33_ASAP7_75t_L g162 ( .A1(n_146), .A2(n_124), .B(n_88), .C(n_96), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_136), .B(n_81), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_149), .B(n_99), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_136), .B(n_100), .Y(n_165) );
BUFx3_ASAP7_75t_L g166 ( .A(n_152), .Y(n_166) );
AO21x1_ASAP7_75t_L g167 ( .A1(n_147), .A2(n_85), .B(n_83), .Y(n_167) );
NOR3xp33_ASAP7_75t_SL g168 ( .A(n_144), .B(n_113), .C(n_112), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_137), .B(n_86), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_137), .B(n_91), .Y(n_170) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_153), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_138), .B(n_92), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_144), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_138), .B(n_95), .Y(n_174) );
INVx3_ASAP7_75t_L g175 ( .A(n_140), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_140), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_161), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_160), .Y(n_178) );
O2A1O1Ixp5_ASAP7_75t_L g179 ( .A1(n_167), .A2(n_105), .B(n_107), .C(n_97), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_160), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_160), .Y(n_181) );
O2A1O1Ixp5_ASAP7_75t_L g182 ( .A1(n_162), .A2(n_93), .B(n_108), .C(n_102), .Y(n_182) );
INVx5_ASAP7_75t_L g183 ( .A(n_175), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_158), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_156), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_155), .B(n_111), .Y(n_186) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_166), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_165), .A2(n_133), .B1(n_103), .B2(n_131), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_173), .B(n_114), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_165), .A2(n_133), .B1(n_119), .B2(n_131), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_159), .A2(n_145), .B(n_143), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_163), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_169), .A2(n_151), .B(n_145), .C(n_143), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_157), .B(n_3), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_169), .A2(n_131), .B1(n_122), .B2(n_123), .Y(n_195) );
NAND2x1_ASAP7_75t_SL g196 ( .A(n_171), .B(n_4), .Y(n_196) );
O2A1O1Ixp33_ASAP7_75t_L g197 ( .A1(n_170), .A2(n_151), .B(n_145), .C(n_143), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_172), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_L g199 ( .A1(n_174), .A2(n_168), .B(n_164), .C(n_176), .Y(n_199) );
OAI21x1_ASAP7_75t_L g200 ( .A1(n_182), .A2(n_191), .B(n_189), .Y(n_200) );
OAI21x1_ASAP7_75t_L g201 ( .A1(n_189), .A2(n_123), .B(n_119), .Y(n_201) );
OAI21x1_ASAP7_75t_L g202 ( .A1(n_193), .A2(n_127), .B(n_125), .Y(n_202) );
OAI21x1_ASAP7_75t_L g203 ( .A1(n_197), .A2(n_127), .B(n_125), .Y(n_203) );
OAI21xp5_ASAP7_75t_L g204 ( .A1(n_179), .A2(n_142), .B(n_135), .Y(n_204) );
NAND3xp33_ASAP7_75t_SL g205 ( .A(n_199), .B(n_5), .C(n_6), .Y(n_205) );
INVx6_ASAP7_75t_L g206 ( .A(n_183), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_184), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_194), .A2(n_150), .B(n_7), .C(n_8), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_186), .A2(n_23), .B(n_22), .Y(n_209) );
INVx4_ASAP7_75t_SL g210 ( .A(n_185), .Y(n_210) );
OAI21x1_ASAP7_75t_L g211 ( .A1(n_178), .A2(n_49), .B(n_69), .Y(n_211) );
OAI21x1_ASAP7_75t_L g212 ( .A1(n_180), .A2(n_46), .B(n_68), .Y(n_212) );
OAI21x1_ASAP7_75t_L g213 ( .A1(n_181), .A2(n_45), .B(n_67), .Y(n_213) );
INVx4_ASAP7_75t_L g214 ( .A(n_183), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_192), .B(n_12), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_198), .B(n_14), .Y(n_216) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_188), .A2(n_41), .B(n_63), .Y(n_217) );
OA21x2_ASAP7_75t_L g218 ( .A1(n_195), .A2(n_36), .B(n_61), .Y(n_218) );
OA21x2_ASAP7_75t_L g219 ( .A1(n_190), .A2(n_50), .B(n_60), .Y(n_219) );
OAI21x1_ASAP7_75t_L g220 ( .A1(n_177), .A2(n_33), .B(n_58), .Y(n_220) );
OR2x6_ASAP7_75t_L g221 ( .A(n_187), .B(n_24), .Y(n_221) );
OA21x2_ASAP7_75t_L g222 ( .A1(n_201), .A2(n_190), .B(n_196), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_207), .B(n_26), .Y(n_223) );
AOI21xp5_ASAP7_75t_SL g224 ( .A1(n_221), .A2(n_30), .B(n_31), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_214), .Y(n_225) );
INVx3_ASAP7_75t_L g226 ( .A(n_206), .Y(n_226) );
AO31x2_ASAP7_75t_L g227 ( .A1(n_208), .A2(n_209), .A3(n_216), .B(n_215), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_204), .A2(n_215), .B(n_216), .C(n_205), .Y(n_228) );
OA21x2_ASAP7_75t_L g229 ( .A1(n_211), .A2(n_213), .B(n_212), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g230 ( .A1(n_217), .A2(n_210), .B1(n_219), .B2(n_218), .Y(n_230) );
INVx3_ASAP7_75t_L g231 ( .A(n_220), .Y(n_231) );
OA21x2_ASAP7_75t_L g232 ( .A1(n_201), .A2(n_203), .B(n_202), .Y(n_232) );
OAI21xp5_ASAP7_75t_L g233 ( .A1(n_200), .A2(n_182), .B(n_162), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_232), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_223), .Y(n_235) );
OR2x6_ASAP7_75t_L g236 ( .A(n_224), .B(n_225), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_222), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_231), .Y(n_238) );
AO21x2_ASAP7_75t_L g239 ( .A1(n_233), .A2(n_228), .B(n_230), .Y(n_239) );
OR2x2_ASAP7_75t_L g240 ( .A(n_227), .B(n_226), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_229), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_240), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_234), .Y(n_243) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_236), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_241), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_239), .B(n_235), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_243), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_243), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_246), .B(n_237), .Y(n_249) );
INVx5_ASAP7_75t_L g250 ( .A(n_244), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_242), .B(n_238), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_247), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_247), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_248), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_252), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_255), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_256), .Y(n_257) );
OAI221xp5_ASAP7_75t_L g258 ( .A1(n_257), .A2(n_250), .B1(n_253), .B2(n_252), .C(n_254), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_258), .Y(n_259) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_259), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_260), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_261), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_262), .Y(n_263) );
BUFx2_ASAP7_75t_L g264 ( .A(n_263), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_264), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_265), .A2(n_249), .B1(n_251), .B2(n_245), .Y(n_266) );
endmodule