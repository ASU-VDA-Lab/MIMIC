module fake_jpeg_12539_n_517 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_517);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_517;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_59),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_60),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_61),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_35),
.B(n_51),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_62),
.B(n_106),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_26),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_63),
.B(n_64),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_29),
.B(n_17),
.C(n_2),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_17),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_66),
.B(n_73),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_67),
.Y(n_151)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

INVx6_ASAP7_75t_SL g69 ( 
.A(n_49),
.Y(n_69)
);

INVx6_ASAP7_75t_SL g183 ( 
.A(n_69),
.Y(n_183)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_70),
.Y(n_136)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_71),
.Y(n_135)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_72),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_17),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_74),
.Y(n_153)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_75),
.Y(n_164)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_76),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_77),
.Y(n_162)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_78),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_19),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_80),
.A2(n_19),
.B1(n_44),
.B2(n_46),
.Y(n_133)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_49),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_82),
.B(n_86),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_83),
.Y(n_173)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_85),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_32),
.B(n_1),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_87),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_88),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_20),
.B(n_32),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_90),
.B(n_101),
.Y(n_163)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_91),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_36),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_92),
.A2(n_37),
.B1(n_36),
.B2(n_55),
.Y(n_149)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_18),
.Y(n_93)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_93),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_94),
.Y(n_191)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_97),
.Y(n_172)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_22),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_98),
.B(n_99),
.Y(n_167)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_23),
.Y(n_100)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_100),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_20),
.B(n_4),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_103),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

BUFx4f_ASAP7_75t_SL g160 ( 
.A(n_104),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx3_ASAP7_75t_SL g168 ( 
.A(n_105),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_41),
.B(n_4),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_22),
.Y(n_107)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_107),
.Y(n_199)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_108),
.Y(n_166)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_22),
.Y(n_109)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_109),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_111),
.Y(n_189)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_112),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_41),
.B(n_6),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_116),
.Y(n_155)
);

BUFx12f_ASAP7_75t_SL g114 ( 
.A(n_23),
.Y(n_114)
);

INVx2_ASAP7_75t_R g131 ( 
.A(n_114),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_42),
.Y(n_115)
);

BUFx4f_ASAP7_75t_L g186 ( 
.A(n_115),
.Y(n_186)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_24),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_20),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_117),
.B(n_118),
.Y(n_177)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_39),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_120),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_45),
.Y(n_120)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_33),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_45),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_122),
.B(n_96),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_100),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_125),
.B(n_127),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_59),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_L g128 ( 
.A1(n_60),
.A2(n_33),
.B1(n_19),
.B2(n_56),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_128),
.A2(n_149),
.B1(n_94),
.B2(n_45),
.Y(n_221)
);

OA22x2_ASAP7_75t_L g215 ( 
.A1(n_133),
.A2(n_139),
.B1(n_196),
.B2(n_147),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_67),
.A2(n_43),
.B1(n_56),
.B2(n_39),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_134),
.A2(n_150),
.B1(n_185),
.B2(n_95),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_61),
.A2(n_33),
.B1(n_37),
.B2(n_36),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_139),
.A2(n_196),
.B1(n_30),
.B2(n_103),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_71),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_140),
.B(n_144),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_78),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_67),
.A2(n_37),
.B1(n_53),
.B2(n_52),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_102),
.A2(n_28),
.B1(n_53),
.B2(n_52),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_152),
.A2(n_30),
.B(n_23),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_114),
.B(n_46),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_156),
.B(n_165),
.Y(n_262)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_108),
.B(n_6),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_159),
.B(n_188),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_81),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_161),
.B(n_174),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_85),
.B(n_44),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_89),
.B(n_25),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_171),
.B(n_192),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_112),
.B(n_25),
.Y(n_174)
);

CKINVDCx12_ASAP7_75t_R g179 ( 
.A(n_115),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_179),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_102),
.A2(n_27),
.B1(n_48),
.B2(n_47),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_68),
.B(n_27),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_70),
.B(n_24),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_195),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_72),
.B(n_28),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_65),
.A2(n_55),
.B1(n_48),
.B2(n_47),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_91),
.B(n_40),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_40),
.Y(n_207)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_200),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_130),
.B(n_80),
.C(n_122),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_201),
.B(n_246),
.Y(n_274)
);

BUFx2_ASAP7_75t_SL g202 ( 
.A(n_183),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_202),
.Y(n_293)
);

INVx11_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_203),
.Y(n_294)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_204),
.B(n_205),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_206),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_207),
.B(n_211),
.Y(n_279)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_198),
.Y(n_208)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_208),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_209),
.A2(n_265),
.B1(n_175),
.B2(n_172),
.Y(n_273)
);

OAI22x1_ASAP7_75t_L g308 ( 
.A1(n_210),
.A2(n_215),
.B1(n_220),
.B2(n_216),
.Y(n_308)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_199),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_166),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_212),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_213),
.B(n_240),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_149),
.A2(n_75),
.B1(n_97),
.B2(n_119),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_214),
.A2(n_224),
.B(n_243),
.Y(n_272)
);

OA22x2_ASAP7_75t_L g216 ( 
.A1(n_133),
.A2(n_121),
.B1(n_77),
.B2(n_83),
.Y(n_216)
);

HAxp5_ASAP7_75t_L g267 ( 
.A(n_216),
.B(n_254),
.CON(n_267),
.SN(n_267)
);

AOI32xp33_ASAP7_75t_L g217 ( 
.A1(n_163),
.A2(n_45),
.A3(n_120),
.B1(n_74),
.B2(n_88),
.Y(n_217)
);

AOI21xp33_ASAP7_75t_L g287 ( 
.A1(n_217),
.A2(n_250),
.B(n_160),
.Y(n_287)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_187),
.Y(n_219)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_219),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_168),
.A2(n_111),
.B1(n_110),
.B2(n_105),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_221),
.A2(n_153),
.B1(n_190),
.B2(n_181),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_129),
.Y(n_222)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_222),
.Y(n_284)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_132),
.Y(n_223)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_223),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_159),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_186),
.Y(n_225)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_225),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_148),
.B(n_7),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_227),
.B(n_248),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_129),
.Y(n_228)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_228),
.Y(n_269)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_186),
.Y(n_231)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_231),
.Y(n_271)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_232),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_182),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_233),
.B(n_234),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_167),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_143),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_235),
.B(n_236),
.Y(n_304)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_178),
.Y(n_236)
);

NAND3xp33_ASAP7_75t_L g237 ( 
.A(n_142),
.B(n_13),
.C(n_8),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_237),
.B(n_241),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_129),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_131),
.Y(n_241)
);

INVx8_ASAP7_75t_L g242 ( 
.A(n_123),
.Y(n_242)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_242),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_131),
.B(n_7),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_243),
.B(n_245),
.Y(n_285)
);

BUFx2_ASAP7_75t_SL g244 ( 
.A(n_160),
.Y(n_244)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_244),
.Y(n_313)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_126),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_167),
.B(n_13),
.C(n_10),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_166),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_247),
.B(n_252),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_197),
.B(n_10),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_128),
.A2(n_11),
.B1(n_13),
.B2(n_177),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_249),
.A2(n_172),
.B1(n_175),
.B2(n_138),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_174),
.B(n_11),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_185),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_155),
.B(n_141),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_253),
.B(n_255),
.Y(n_314)
);

OA22x2_ASAP7_75t_L g254 ( 
.A1(n_134),
.A2(n_145),
.B1(n_189),
.B2(n_170),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_157),
.B(n_193),
.Y(n_255)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_132),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_256),
.B(n_257),
.Y(n_295)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_193),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_158),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_258),
.B(n_259),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_150),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_170),
.B(n_189),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_146),
.Y(n_289)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_168),
.A2(n_145),
.B1(n_191),
.B2(n_162),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_261),
.A2(n_138),
.B1(n_147),
.B2(n_137),
.Y(n_275)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_136),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_263),
.B(n_264),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_124),
.Y(n_264)
);

OA22x2_ASAP7_75t_L g265 ( 
.A1(n_123),
.A2(n_162),
.B1(n_173),
.B2(n_137),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_268),
.A2(n_292),
.B1(n_298),
.B2(n_301),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_272),
.B(n_287),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_273),
.A2(n_278),
.B1(n_309),
.B2(n_312),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g324 ( 
.A1(n_275),
.A2(n_265),
.B1(n_254),
.B2(n_231),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_238),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_277),
.B(n_303),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_209),
.A2(n_191),
.B1(n_173),
.B2(n_146),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_252),
.A2(n_151),
.B(n_164),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_280),
.A2(n_213),
.B(n_205),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_259),
.A2(n_176),
.B1(n_180),
.B2(n_154),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_282),
.A2(n_313),
.B(n_306),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_229),
.B(n_135),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_286),
.B(n_289),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_214),
.A2(n_221),
.B1(n_201),
.B2(n_215),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_216),
.A2(n_153),
.B1(n_190),
.B2(n_124),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_216),
.A2(n_158),
.B1(n_215),
.B2(n_226),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_302),
.A2(n_311),
.B1(n_300),
.B2(n_293),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_260),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_308),
.A2(n_254),
.B1(n_240),
.B2(n_246),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_229),
.A2(n_158),
.B1(n_215),
.B2(n_250),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_251),
.A2(n_207),
.B1(n_248),
.B2(n_229),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_250),
.A2(n_265),
.B1(n_254),
.B2(n_218),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_203),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_293),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_274),
.B(n_227),
.C(n_262),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_317),
.B(n_328),
.C(n_342),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_318),
.A2(n_324),
.B1(n_294),
.B2(n_297),
.Y(n_365)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_283),
.Y(n_319)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_319),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_310),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_320),
.B(n_327),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_322),
.B(n_333),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_309),
.A2(n_267),
.B1(n_312),
.B2(n_303),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_323),
.A2(n_335),
.B1(n_336),
.B2(n_349),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_325),
.A2(n_269),
.B(n_290),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_310),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_274),
.B(n_230),
.C(n_208),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_289),
.Y(n_329)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_329),
.Y(n_361)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_291),
.Y(n_331)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_331),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_281),
.B(n_224),
.Y(n_333)
);

BUFx12f_ASAP7_75t_L g334 ( 
.A(n_316),
.Y(n_334)
);

INVx13_ASAP7_75t_L g379 ( 
.A(n_334),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_267),
.A2(n_273),
.B1(n_292),
.B2(n_302),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_267),
.A2(n_265),
.B1(n_239),
.B2(n_242),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_304),
.Y(n_337)
);

INVx13_ASAP7_75t_L g383 ( 
.A(n_337),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_277),
.B(n_263),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_338),
.B(n_337),
.Y(n_371)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_291),
.Y(n_339)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_339),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_286),
.B(n_206),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_340),
.B(n_300),
.Y(n_370)
);

OAI21xp33_ASAP7_75t_L g341 ( 
.A1(n_310),
.A2(n_257),
.B(n_247),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_341),
.A2(n_351),
.B1(n_352),
.B2(n_283),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_311),
.B(n_232),
.C(n_264),
.Y(n_342)
);

OAI32xp33_ASAP7_75t_L g343 ( 
.A1(n_314),
.A2(n_219),
.A3(n_223),
.B1(n_256),
.B2(n_225),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_343),
.B(n_347),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_281),
.B(n_222),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_344),
.B(n_350),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_266),
.B(n_228),
.C(n_296),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_346),
.B(n_307),
.C(n_315),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_304),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_270),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_348),
.B(n_299),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_308),
.A2(n_278),
.B1(n_272),
.B2(n_314),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_279),
.B(n_270),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_288),
.A2(n_275),
.B1(n_301),
.B2(n_280),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_282),
.A2(n_279),
.B1(n_268),
.B2(n_285),
.Y(n_352)
);

OAI22x1_ASAP7_75t_L g385 ( 
.A1(n_353),
.A2(n_290),
.B1(n_315),
.B2(n_305),
.Y(n_385)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_295),
.Y(n_354)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_354),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_355),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_321),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_356),
.B(n_357),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_321),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_328),
.B(n_276),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_359),
.B(n_386),
.C(n_387),
.Y(n_391)
);

AO22x1_ASAP7_75t_L g362 ( 
.A1(n_323),
.A2(n_313),
.B1(n_297),
.B2(n_294),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_362),
.A2(n_372),
.B(n_373),
.Y(n_411)
);

O2A1O1Ixp33_ASAP7_75t_L g364 ( 
.A1(n_325),
.A2(n_335),
.B(n_322),
.C(n_326),
.Y(n_364)
);

OAI21xp33_ASAP7_75t_L g409 ( 
.A1(n_364),
.A2(n_356),
.B(n_357),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_365),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g408 ( 
.A(n_370),
.B(n_384),
.Y(n_408)
);

CKINVDCx14_ASAP7_75t_R g414 ( 
.A(n_371),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_350),
.B(n_299),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_374),
.B(n_375),
.Y(n_398)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_331),
.Y(n_381)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_381),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_355),
.A2(n_269),
.B(n_284),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_382),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_317),
.B(n_284),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_385),
.B(n_336),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_340),
.B(n_305),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_376),
.A2(n_318),
.B1(n_332),
.B2(n_353),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_388),
.A2(n_390),
.B1(n_395),
.B2(n_399),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_376),
.A2(n_332),
.B1(n_329),
.B2(n_349),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_393),
.B(n_397),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_384),
.B(n_340),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_394),
.B(n_403),
.C(n_404),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_372),
.A2(n_345),
.B1(n_344),
.B2(n_330),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_383),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_361),
.A2(n_345),
.B1(n_351),
.B2(n_330),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_360),
.Y(n_400)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_400),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_383),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_402),
.B(n_405),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_377),
.B(n_326),
.C(n_342),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_377),
.B(n_326),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_369),
.Y(n_405)
);

FAx1_ASAP7_75t_SL g406 ( 
.A(n_378),
.B(n_333),
.CI(n_346),
.CON(n_406),
.SN(n_406)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_406),
.B(n_386),
.Y(n_420)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_366),
.Y(n_407)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_407),
.Y(n_418)
);

OA22x2_ASAP7_75t_L g419 ( 
.A1(n_409),
.A2(n_373),
.B1(n_362),
.B2(n_382),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_358),
.A2(n_354),
.B1(n_347),
.B2(n_352),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_410),
.B(n_412),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_361),
.A2(n_380),
.B1(n_369),
.B2(n_364),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_380),
.A2(n_343),
.B1(n_338),
.B2(n_334),
.Y(n_413)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_413),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_408),
.B(n_370),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_415),
.B(n_420),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_419),
.B(n_423),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_404),
.B(n_391),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_421),
.B(n_437),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_398),
.B(n_368),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_389),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_427),
.B(n_397),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_410),
.B(n_368),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_428),
.B(n_433),
.Y(n_449)
);

AND2x6_ASAP7_75t_L g429 ( 
.A(n_414),
.B(n_362),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_412),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_411),
.A2(n_378),
.B(n_363),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_430),
.A2(n_432),
.B(n_405),
.Y(n_440)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_389),
.Y(n_431)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_431),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_411),
.A2(n_371),
.B(n_374),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_401),
.A2(n_365),
.B1(n_387),
.B2(n_366),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_434),
.A2(n_395),
.B1(n_399),
.B2(n_413),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_391),
.B(n_359),
.C(n_381),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_435),
.B(n_438),
.C(n_403),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_401),
.A2(n_367),
.B1(n_385),
.B2(n_360),
.Y(n_436)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_436),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_408),
.B(n_367),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_394),
.B(n_339),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_439),
.B(n_440),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_443),
.A2(n_449),
.B1(n_417),
.B2(n_424),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_426),
.B(n_402),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_444),
.B(n_446),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_445),
.A2(n_417),
.B1(n_424),
.B2(n_447),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_421),
.B(n_388),
.Y(n_446)
);

NOR3xp33_ASAP7_75t_L g472 ( 
.A(n_448),
.B(n_451),
.C(n_458),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_433),
.B(n_406),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_422),
.B(n_392),
.C(n_390),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_452),
.B(n_453),
.C(n_456),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_422),
.B(n_406),
.C(n_393),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_426),
.B(n_400),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_454),
.B(n_455),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_435),
.B(n_407),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_438),
.B(n_396),
.C(n_319),
.Y(n_456)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_431),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_457),
.B(n_437),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_461),
.B(n_469),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_462),
.A2(n_470),
.B1(n_419),
.B2(n_456),
.Y(n_477)
);

FAx1_ASAP7_75t_SL g463 ( 
.A(n_453),
.B(n_432),
.CI(n_430),
.CON(n_463),
.SN(n_463)
);

A2O1A1O1Ixp25_ASAP7_75t_L g484 ( 
.A1(n_463),
.A2(n_450),
.B(n_379),
.C(n_334),
.D(n_271),
.Y(n_484)
);

BUFx24_ASAP7_75t_SL g465 ( 
.A(n_440),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_465),
.B(n_468),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_466),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_445),
.A2(n_425),
.B1(n_418),
.B2(n_429),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_443),
.A2(n_425),
.B(n_416),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_441),
.A2(n_434),
.B1(n_419),
.B2(n_416),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_457),
.B(n_415),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_471),
.B(n_473),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_442),
.A2(n_419),
.B(n_418),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_460),
.B(n_455),
.C(n_439),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_474),
.B(n_475),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_470),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_473),
.A2(n_444),
.B1(n_452),
.B2(n_454),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_476),
.A2(n_459),
.B1(n_462),
.B2(n_461),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_477),
.A2(n_464),
.B1(n_463),
.B2(n_271),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_472),
.A2(n_396),
.B1(n_400),
.B2(n_446),
.Y(n_480)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_480),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_460),
.B(n_450),
.C(n_379),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_483),
.A2(n_485),
.B(n_471),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_484),
.A2(n_483),
.B(n_477),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_464),
.B(n_307),
.C(n_334),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_474),
.B(n_467),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_486),
.B(n_491),
.Y(n_502)
);

INVxp67_ASAP7_75t_SL g497 ( 
.A(n_489),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_490),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_481),
.B(n_467),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_481),
.B(n_459),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_492),
.B(n_494),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_493),
.B(n_495),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_485),
.A2(n_463),
.B(n_271),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_486),
.B(n_478),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_499),
.B(n_500),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_487),
.B(n_491),
.C(n_492),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_488),
.B(n_479),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_501),
.B(n_476),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_500),
.B(n_502),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_505),
.B(n_506),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_498),
.B(n_493),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_507),
.A2(n_508),
.B(n_496),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_498),
.A2(n_484),
.B(n_482),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_503),
.B(n_482),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_509),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_511),
.B(n_504),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_513),
.A2(n_514),
.B(n_509),
.Y(n_515)
);

INVxp33_ASAP7_75t_SL g514 ( 
.A(n_512),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_515),
.B(n_510),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_497),
.Y(n_517)
);


endmodule