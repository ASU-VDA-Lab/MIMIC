module fake_aes_11309_n_648 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_648);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_648;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_575;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_482;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_446;
wire n_195;
wire n_420;
wire n_423;
wire n_342;
wire n_165;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g75 ( .A(n_69), .Y(n_75) );
INVx2_ASAP7_75t_L g76 ( .A(n_28), .Y(n_76) );
INVxp67_ASAP7_75t_SL g77 ( .A(n_44), .Y(n_77) );
BUFx6f_ASAP7_75t_L g78 ( .A(n_20), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_43), .Y(n_79) );
INVxp33_ASAP7_75t_SL g80 ( .A(n_2), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_59), .Y(n_81) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_67), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_30), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_62), .Y(n_84) );
HB1xp67_ASAP7_75t_L g85 ( .A(n_48), .Y(n_85) );
INVx3_ASAP7_75t_L g86 ( .A(n_34), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_45), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_39), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_23), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_12), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_0), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_8), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_2), .Y(n_93) );
INVxp33_ASAP7_75t_SL g94 ( .A(n_53), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_70), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_65), .Y(n_96) );
INVxp67_ASAP7_75t_SL g97 ( .A(n_33), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_40), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_64), .Y(n_99) );
CKINVDCx16_ASAP7_75t_R g100 ( .A(n_7), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_16), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_38), .Y(n_102) );
CKINVDCx14_ASAP7_75t_R g103 ( .A(n_68), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_49), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_18), .Y(n_105) );
INVxp67_ASAP7_75t_L g106 ( .A(n_17), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_5), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_46), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_56), .Y(n_109) );
OR2x2_ASAP7_75t_L g110 ( .A(n_54), .B(n_1), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_14), .Y(n_111) );
INVx1_ASAP7_75t_SL g112 ( .A(n_42), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_47), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_22), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_72), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_7), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_31), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_36), .Y(n_118) );
CKINVDCx14_ASAP7_75t_R g119 ( .A(n_21), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_25), .Y(n_120) );
OA21x2_ASAP7_75t_L g121 ( .A1(n_76), .A2(n_29), .B(n_73), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_75), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_103), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_85), .B(n_0), .Y(n_124) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_80), .A2(n_1), .B1(n_3), .B2(n_4), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_83), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_100), .B(n_3), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_86), .B(n_4), .Y(n_128) );
INVx3_ASAP7_75t_L g129 ( .A(n_86), .Y(n_129) );
AOI22xp5_ASAP7_75t_L g130 ( .A1(n_80), .A2(n_5), .B1(n_6), .B2(n_8), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_84), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_86), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_95), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_96), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_98), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_99), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_90), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_91), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_76), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_92), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_78), .B(n_6), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_102), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_104), .Y(n_143) );
OAI21x1_ASAP7_75t_L g144 ( .A1(n_105), .A2(n_41), .B(n_71), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_78), .Y(n_145) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_93), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_109), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_114), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_115), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_103), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_107), .B(n_9), .Y(n_151) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_116), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_119), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_118), .Y(n_154) );
OAI22xp5_ASAP7_75t_SL g155 ( .A1(n_82), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_77), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_97), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_106), .B(n_10), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_110), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_78), .Y(n_160) );
BUFx2_ASAP7_75t_L g161 ( .A(n_152), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_145), .Y(n_162) );
AND2x6_ASAP7_75t_L g163 ( .A(n_158), .B(n_78), .Y(n_163) );
INVx1_ASAP7_75t_SL g164 ( .A(n_127), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_145), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_145), .Y(n_166) );
INVxp67_ASAP7_75t_SL g167 ( .A(n_159), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_145), .Y(n_168) );
BUFx10_ASAP7_75t_L g169 ( .A(n_123), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_129), .Y(n_170) );
INVx4_ASAP7_75t_L g171 ( .A(n_129), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_159), .B(n_119), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_145), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_132), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_123), .B(n_79), .Y(n_175) );
AOI22xp33_ASAP7_75t_L g176 ( .A1(n_156), .A2(n_157), .B1(n_159), .B2(n_146), .Y(n_176) );
BUFx3_ASAP7_75t_L g177 ( .A(n_129), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_132), .Y(n_178) );
NAND3xp33_ASAP7_75t_L g179 ( .A(n_156), .B(n_79), .C(n_81), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_157), .B(n_81), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_139), .Y(n_181) );
INVx3_ASAP7_75t_L g182 ( .A(n_139), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_122), .B(n_113), .Y(n_183) );
INVx6_ASAP7_75t_L g184 ( .A(n_158), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_122), .B(n_94), .Y(n_185) );
BUFx3_ASAP7_75t_L g186 ( .A(n_121), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_137), .B(n_113), .Y(n_187) );
BUFx3_ASAP7_75t_L g188 ( .A(n_121), .Y(n_188) );
NAND2x1p5_ASAP7_75t_L g189 ( .A(n_158), .B(n_112), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_150), .B(n_94), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_121), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_160), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_121), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_160), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_147), .Y(n_195) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_150), .Y(n_196) );
AOI21x1_ASAP7_75t_L g197 ( .A1(n_128), .A2(n_120), .B(n_117), .Y(n_197) );
BUFx4f_ASAP7_75t_L g198 ( .A(n_126), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_126), .B(n_111), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_147), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_144), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_148), .Y(n_202) );
BUFx2_ASAP7_75t_L g203 ( .A(n_153), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_148), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_149), .Y(n_205) );
AND2x2_ASAP7_75t_SL g206 ( .A(n_124), .B(n_101), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_131), .B(n_108), .Y(n_207) );
NAND3x1_ASAP7_75t_L g208 ( .A(n_125), .B(n_82), .C(n_101), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_149), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_131), .B(n_89), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_154), .Y(n_211) );
AND2x4_ASAP7_75t_SL g212 ( .A(n_127), .B(n_88), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_154), .Y(n_213) );
AO22x2_ASAP7_75t_L g214 ( .A1(n_133), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_138), .B(n_87), .Y(n_215) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_161), .Y(n_216) );
BUFx4f_ASAP7_75t_L g217 ( .A(n_189), .Y(n_217) );
BUFx8_ASAP7_75t_L g218 ( .A(n_161), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_171), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_192), .Y(n_220) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_176), .A2(n_130), .B1(n_153), .B2(n_142), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_191), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_172), .B(n_133), .Y(n_223) );
INVx1_ASAP7_75t_SL g224 ( .A(n_164), .Y(n_224) );
CKINVDCx8_ASAP7_75t_R g225 ( .A(n_203), .Y(n_225) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_172), .Y(n_226) );
BUFx2_ASAP7_75t_L g227 ( .A(n_203), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_192), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_163), .A2(n_134), .B1(n_135), .B2(n_143), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_187), .B(n_134), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_177), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_185), .B(n_142), .Y(n_232) );
BUFx2_ASAP7_75t_L g233 ( .A(n_196), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_191), .Y(n_234) );
BUFx2_ASAP7_75t_L g235 ( .A(n_180), .Y(n_235) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_191), .Y(n_236) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_187), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_163), .A2(n_135), .B1(n_136), .B2(n_143), .Y(n_238) );
OAI21xp5_ASAP7_75t_L g239 ( .A1(n_186), .A2(n_144), .B(n_136), .Y(n_239) );
AND2x4_ASAP7_75t_L g240 ( .A(n_180), .B(n_140), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_177), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_163), .A2(n_151), .B1(n_155), .B2(n_141), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_167), .B(n_15), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_171), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_171), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_170), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_198), .B(n_19), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_212), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_170), .Y(n_249) );
AND2x4_ASAP7_75t_L g250 ( .A(n_215), .B(n_24), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_170), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_202), .Y(n_252) );
INVx2_ASAP7_75t_SL g253 ( .A(n_189), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_212), .Y(n_254) );
NOR3xp33_ASAP7_75t_SL g255 ( .A(n_179), .B(n_26), .C(n_27), .Y(n_255) );
NAND3xp33_ASAP7_75t_L g256 ( .A(n_179), .B(n_32), .C(n_35), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_183), .B(n_37), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_215), .B(n_50), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_202), .Y(n_259) );
INVx2_ASAP7_75t_SL g260 ( .A(n_189), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_198), .B(n_51), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_204), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_209), .Y(n_263) );
INVx5_ASAP7_75t_L g264 ( .A(n_163), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_209), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_204), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_163), .A2(n_52), .B1(n_55), .B2(n_57), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_198), .B(n_58), .Y(n_268) );
OAI22xp5_ASAP7_75t_SL g269 ( .A1(n_206), .A2(n_60), .B1(n_61), .B2(n_63), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_199), .B(n_66), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_205), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_209), .B(n_74), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_214), .Y(n_273) );
INVx2_ASAP7_75t_SL g274 ( .A(n_217), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_223), .A2(n_186), .B(n_188), .Y(n_275) );
INVxp67_ASAP7_75t_SL g276 ( .A(n_273), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_226), .Y(n_277) );
INVx5_ASAP7_75t_L g278 ( .A(n_264), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_226), .B(n_210), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_237), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_220), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_220), .Y(n_282) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_222), .Y(n_283) );
A2O1A1Ixp33_ASAP7_75t_L g284 ( .A1(n_232), .A2(n_213), .B(n_205), .C(n_178), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_239), .A2(n_188), .B(n_193), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_216), .B(n_190), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g287 ( .A(n_218), .Y(n_287) );
AO21x2_ASAP7_75t_L g288 ( .A1(n_247), .A2(n_174), .B(n_178), .Y(n_288) );
NOR2x1p5_ASAP7_75t_SL g289 ( .A(n_272), .B(n_197), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_237), .B(n_184), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_219), .Y(n_291) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_224), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_253), .B(n_197), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_240), .Y(n_294) );
AND2x4_ASAP7_75t_L g295 ( .A(n_260), .B(n_175), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_240), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_244), .A2(n_191), .B(n_193), .Y(n_297) );
AND2x4_ASAP7_75t_L g298 ( .A(n_230), .B(n_163), .Y(n_298) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_216), .Y(n_299) );
BUFx3_ASAP7_75t_L g300 ( .A(n_264), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_230), .Y(n_301) );
CKINVDCx10_ASAP7_75t_R g302 ( .A(n_218), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_227), .B(n_206), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_252), .Y(n_304) );
AND2x4_ASAP7_75t_L g305 ( .A(n_235), .B(n_163), .Y(n_305) );
CKINVDCx20_ASAP7_75t_R g306 ( .A(n_225), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_245), .A2(n_193), .B(n_191), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g308 ( .A1(n_217), .A2(n_184), .B1(n_206), .B2(n_214), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_250), .B(n_207), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_228), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_259), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_250), .B(n_201), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_221), .B(n_184), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_262), .Y(n_314) );
OR2x6_ASAP7_75t_L g315 ( .A(n_233), .B(n_208), .Y(n_315) );
OAI22xp5_ASAP7_75t_L g316 ( .A1(n_273), .A2(n_184), .B1(n_214), .B2(n_208), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_266), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_258), .B(n_213), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_271), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_281), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_304), .Y(n_321) );
OAI21x1_ASAP7_75t_L g322 ( .A1(n_285), .A2(n_261), .B(n_268), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_274), .B(n_246), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_299), .B(n_174), .Y(n_324) );
OR2x2_ASAP7_75t_L g325 ( .A(n_292), .B(n_254), .Y(n_325) );
OA21x2_ASAP7_75t_L g326 ( .A1(n_297), .A2(n_255), .B(n_256), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_313), .B(n_242), .Y(n_327) );
INVx3_ASAP7_75t_SL g328 ( .A(n_287), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_281), .Y(n_329) );
OAI21xp5_ASAP7_75t_L g330 ( .A1(n_275), .A2(n_261), .B(n_247), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_292), .B(n_248), .Y(n_331) );
OA21x2_ASAP7_75t_L g332 ( .A1(n_307), .A2(n_255), .B(n_268), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_299), .B(n_249), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_319), .Y(n_334) );
XOR2xp5_ASAP7_75t_L g335 ( .A(n_287), .B(n_242), .Y(n_335) );
NAND2xp33_ASAP7_75t_SL g336 ( .A(n_306), .B(n_269), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_311), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_303), .B(n_200), .Y(n_338) );
OAI21x1_ASAP7_75t_L g339 ( .A1(n_308), .A2(n_270), .B(n_257), .Y(n_339) );
INVx3_ASAP7_75t_L g340 ( .A(n_300), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_282), .Y(n_341) );
NAND2x1p5_ASAP7_75t_L g342 ( .A(n_278), .B(n_264), .Y(n_342) );
INVxp67_ASAP7_75t_SL g343 ( .A(n_276), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_313), .B(n_251), .Y(n_344) );
OAI21x1_ASAP7_75t_L g345 ( .A1(n_312), .A2(n_243), .B(n_267), .Y(n_345) );
OAI21x1_ASAP7_75t_L g346 ( .A1(n_312), .A2(n_267), .B(n_238), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_314), .Y(n_347) );
OA21x2_ASAP7_75t_L g348 ( .A1(n_284), .A2(n_181), .B(n_238), .Y(n_348) );
OAI21x1_ASAP7_75t_L g349 ( .A1(n_322), .A2(n_282), .B(n_310), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_343), .A2(n_276), .B1(n_316), .B2(n_309), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_321), .B(n_317), .Y(n_351) );
OAI22xp33_ASAP7_75t_L g352 ( .A1(n_328), .A2(n_315), .B1(n_306), .B2(n_279), .Y(n_352) );
AOI222xp33_ASAP7_75t_L g353 ( .A1(n_336), .A2(n_280), .B1(n_277), .B2(n_294), .C1(n_296), .C2(n_301), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_324), .B(n_290), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_320), .Y(n_355) );
NAND3xp33_ASAP7_75t_L g356 ( .A(n_330), .B(n_284), .C(n_293), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_343), .A2(n_318), .B1(n_315), .B2(n_290), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_324), .B(n_310), .Y(n_358) );
INVx2_ASAP7_75t_SL g359 ( .A(n_342), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_321), .B(n_286), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_328), .Y(n_361) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_325), .Y(n_362) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_325), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_335), .A2(n_315), .B1(n_293), .B2(n_295), .Y(n_364) );
OAI22xp33_ASAP7_75t_L g365 ( .A1(n_328), .A2(n_302), .B1(n_318), .B2(n_291), .Y(n_365) );
AOI222xp33_ASAP7_75t_L g366 ( .A1(n_327), .A2(n_214), .B1(n_295), .B2(n_305), .C1(n_298), .C2(n_181), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_337), .B(n_211), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_320), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_334), .B(n_305), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_335), .A2(n_298), .B1(n_169), .B2(n_211), .Y(n_370) );
AOI21xp5_ASAP7_75t_L g371 ( .A1(n_330), .A2(n_283), .B(n_288), .Y(n_371) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_342), .Y(n_372) );
AO21x2_ASAP7_75t_L g373 ( .A1(n_339), .A2(n_288), .B(n_289), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_320), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_368), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_358), .B(n_347), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_358), .B(n_347), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_368), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_351), .B(n_337), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_355), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_355), .Y(n_381) );
NOR2x1_ASAP7_75t_L g382 ( .A(n_365), .B(n_331), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_351), .B(n_329), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_374), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_351), .B(n_329), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_351), .B(n_329), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_374), .B(n_362), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_367), .B(n_341), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_349), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_349), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_367), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_372), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_359), .B(n_341), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_372), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_363), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_361), .Y(n_396) );
AND2x4_ASAP7_75t_L g397 ( .A(n_359), .B(n_372), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_353), .B(n_341), .Y(n_398) );
AND2x4_ASAP7_75t_L g399 ( .A(n_372), .B(n_334), .Y(n_399) );
AND2x4_ASAP7_75t_L g400 ( .A(n_372), .B(n_340), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_356), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_357), .B(n_327), .Y(n_402) );
OR2x2_ASAP7_75t_L g403 ( .A(n_354), .B(n_331), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_366), .B(n_348), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_360), .B(n_348), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_352), .B(n_338), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_356), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_381), .B(n_373), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_381), .B(n_373), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_380), .Y(n_410) );
OR2x6_ASAP7_75t_L g411 ( .A(n_402), .B(n_350), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_376), .B(n_364), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_387), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_387), .Y(n_414) );
OA21x2_ASAP7_75t_L g415 ( .A1(n_389), .A2(n_371), .B(n_339), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_388), .B(n_373), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_380), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_388), .B(n_348), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_384), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_383), .B(n_348), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_384), .B(n_344), .Y(n_421) );
AO21x2_ASAP7_75t_L g422 ( .A1(n_389), .A2(n_390), .B(n_339), .Y(n_422) );
AND2x4_ASAP7_75t_L g423 ( .A(n_392), .B(n_340), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_390), .Y(n_424) );
INVxp67_ASAP7_75t_L g425 ( .A(n_382), .Y(n_425) );
NAND3xp33_ASAP7_75t_L g426 ( .A(n_395), .B(n_361), .C(n_370), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_375), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_383), .B(n_338), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_385), .B(n_369), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_404), .A2(n_333), .B1(n_344), .B2(n_323), .Y(n_430) );
INVxp67_ASAP7_75t_SL g431 ( .A(n_375), .Y(n_431) );
NAND3xp33_ASAP7_75t_L g432 ( .A(n_401), .B(n_332), .C(n_326), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_402), .B(n_182), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_378), .Y(n_434) );
NOR3xp33_ASAP7_75t_L g435 ( .A(n_403), .B(n_182), .C(n_200), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_385), .B(n_346), .Y(n_436) );
INVx3_ASAP7_75t_L g437 ( .A(n_397), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_378), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_386), .B(n_346), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_405), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_394), .Y(n_441) );
AND2x4_ASAP7_75t_SL g442 ( .A(n_379), .B(n_340), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_386), .B(n_346), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_396), .B(n_323), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_394), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_405), .Y(n_446) );
NAND5xp2_ASAP7_75t_L g447 ( .A(n_406), .B(n_229), .C(n_342), .D(n_169), .E(n_332), .Y(n_447) );
AND2x4_ASAP7_75t_L g448 ( .A(n_392), .B(n_340), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_376), .B(n_332), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_379), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_393), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_401), .Y(n_452) );
AND2x4_ASAP7_75t_L g453 ( .A(n_397), .B(n_322), .Y(n_453) );
INVx3_ASAP7_75t_L g454 ( .A(n_397), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_440), .B(n_407), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_416), .B(n_407), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_413), .B(n_391), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_444), .B(n_396), .Y(n_458) );
NAND2x1_ASAP7_75t_L g459 ( .A(n_434), .B(n_438), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_414), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_410), .Y(n_461) );
AND2x4_ASAP7_75t_L g462 ( .A(n_437), .B(n_399), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_416), .B(n_404), .Y(n_463) );
BUFx2_ASAP7_75t_L g464 ( .A(n_431), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_410), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_424), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_447), .A2(n_398), .B1(n_391), .B2(n_399), .Y(n_467) );
NAND3xp33_ASAP7_75t_L g468 ( .A(n_425), .B(n_403), .C(n_399), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_440), .B(n_377), .Y(n_469) );
NAND3xp33_ASAP7_75t_L g470 ( .A(n_426), .B(n_398), .C(n_377), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_446), .B(n_393), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_424), .Y(n_472) );
BUFx3_ASAP7_75t_L g473 ( .A(n_442), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_417), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_450), .B(n_400), .Y(n_475) );
NOR2xp67_ASAP7_75t_L g476 ( .A(n_432), .B(n_400), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_417), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_419), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_437), .B(n_400), .Y(n_479) );
INVx4_ASAP7_75t_L g480 ( .A(n_423), .Y(n_480) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_451), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_446), .B(n_182), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_449), .B(n_332), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_419), .B(n_195), .Y(n_484) );
INVxp67_ASAP7_75t_SL g485 ( .A(n_427), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_449), .B(n_322), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_436), .B(n_326), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_427), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_436), .B(n_326), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_439), .B(n_326), .Y(n_490) );
INVx1_ASAP7_75t_SL g491 ( .A(n_442), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_434), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_452), .B(n_195), .Y(n_493) );
BUFx3_ASAP7_75t_L g494 ( .A(n_437), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_439), .B(n_345), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_438), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_443), .B(n_345), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_443), .B(n_345), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_452), .B(n_333), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_408), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_421), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_408), .B(n_333), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_412), .B(n_323), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_420), .B(n_201), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_420), .B(n_201), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_411), .A2(n_333), .B1(n_323), .B2(n_201), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_409), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_409), .Y(n_508) );
BUFx2_ASAP7_75t_L g509 ( .A(n_454), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_471), .B(n_456), .Y(n_510) );
NAND2x1_ASAP7_75t_L g511 ( .A(n_464), .B(n_411), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_460), .B(n_418), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_471), .B(n_454), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g514 ( .A1(n_482), .A2(n_435), .B(n_433), .C(n_421), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_456), .B(n_454), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_466), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_470), .A2(n_411), .B1(n_430), .B2(n_429), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_481), .B(n_418), .Y(n_518) );
NAND2xp33_ASAP7_75t_SL g519 ( .A(n_464), .B(n_433), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_466), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_501), .B(n_429), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_463), .B(n_462), .Y(n_522) );
AND2x4_ASAP7_75t_L g523 ( .A(n_480), .B(n_453), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_503), .A2(n_411), .B1(n_428), .B2(n_453), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_469), .B(n_428), .Y(n_525) );
INVx1_ASAP7_75t_SL g526 ( .A(n_491), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_467), .A2(n_411), .B1(n_448), .B2(n_423), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_463), .B(n_453), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_462), .B(n_453), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_457), .B(n_441), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_469), .B(n_441), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_502), .B(n_445), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_459), .Y(n_533) );
INVx1_ASAP7_75t_SL g534 ( .A(n_473), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_472), .Y(n_535) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_459), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_468), .B(n_448), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_507), .B(n_445), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_462), .B(n_448), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_477), .Y(n_540) );
OR2x6_ASAP7_75t_L g541 ( .A(n_473), .B(n_448), .Y(n_541) );
NOR2xp67_ASAP7_75t_L g542 ( .A(n_480), .B(n_432), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_507), .B(n_423), .Y(n_543) );
INVxp67_ASAP7_75t_L g544 ( .A(n_485), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_479), .B(n_508), .Y(n_545) );
NAND2xp33_ASAP7_75t_L g546 ( .A(n_506), .B(n_423), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_479), .B(n_422), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_477), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_502), .B(n_422), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_478), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_479), .B(n_422), .Y(n_551) );
INVxp67_ASAP7_75t_L g552 ( .A(n_509), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_500), .B(n_415), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_478), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_455), .B(n_415), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_455), .B(n_415), .Y(n_556) );
INVxp33_ASAP7_75t_L g557 ( .A(n_476), .Y(n_557) );
AND2x2_ASAP7_75t_SL g558 ( .A(n_480), .B(n_415), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_544), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_525), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_510), .B(n_500), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_526), .B(n_458), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_555), .B(n_508), .Y(n_563) );
OAI221xp5_ASAP7_75t_L g564 ( .A1(n_517), .A2(n_509), .B1(n_475), .B2(n_494), .C(n_465), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_555), .B(n_461), .Y(n_565) );
AOI22xp33_ASAP7_75t_SL g566 ( .A1(n_534), .A2(n_494), .B1(n_483), .B2(n_492), .Y(n_566) );
INVx1_ASAP7_75t_SL g567 ( .A(n_518), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_540), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_548), .Y(n_569) );
INVx1_ASAP7_75t_SL g570 ( .A(n_532), .Y(n_570) );
O2A1O1Ixp5_ASAP7_75t_L g571 ( .A1(n_519), .A2(n_474), .B(n_496), .C(n_472), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_519), .A2(n_484), .B(n_499), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_550), .Y(n_573) );
CKINVDCx20_ASAP7_75t_R g574 ( .A(n_522), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_556), .B(n_486), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_512), .B(n_486), .Y(n_576) );
OAI22xp33_ASAP7_75t_SL g577 ( .A1(n_511), .A2(n_499), .B1(n_482), .B2(n_493), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_524), .A2(n_493), .B1(n_488), .B2(n_483), .Y(n_578) );
AOI31xp33_ASAP7_75t_L g579 ( .A1(n_557), .A2(n_490), .A3(n_487), .B(n_489), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_521), .B(n_498), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_556), .B(n_487), .Y(n_581) );
CKINVDCx16_ASAP7_75t_R g582 ( .A(n_541), .Y(n_582) );
NOR4xp25_ASAP7_75t_SL g583 ( .A(n_554), .B(n_505), .C(n_504), .D(n_490), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_531), .Y(n_584) );
OAI31xp33_ASAP7_75t_L g585 ( .A1(n_527), .A2(n_489), .A3(n_495), .B(n_497), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_528), .B(n_495), .Y(n_586) );
OAI22xp33_ASAP7_75t_L g587 ( .A1(n_541), .A2(n_488), .B1(n_497), .B2(n_498), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_530), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_544), .B(n_505), .Y(n_589) );
NOR3xp33_ASAP7_75t_L g590 ( .A(n_514), .B(n_504), .C(n_263), .Y(n_590) );
AOI221xp5_ASAP7_75t_L g591 ( .A1(n_524), .A2(n_201), .B1(n_165), .B2(n_166), .C(n_168), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_538), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_515), .B(n_193), .Y(n_593) );
OAI221xp5_ASAP7_75t_L g594 ( .A1(n_585), .A2(n_537), .B1(n_546), .B2(n_542), .C(n_552), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_592), .Y(n_595) );
AND2x4_ASAP7_75t_L g596 ( .A(n_559), .B(n_551), .Y(n_596) );
INVxp67_ASAP7_75t_L g597 ( .A(n_562), .Y(n_597) );
NOR4xp25_ASAP7_75t_L g598 ( .A(n_564), .B(n_552), .C(n_537), .D(n_547), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_588), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_578), .A2(n_513), .B1(n_543), .B2(n_529), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_568), .Y(n_601) );
CKINVDCx16_ASAP7_75t_R g602 ( .A(n_582), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_574), .B(n_557), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_565), .B(n_549), .Y(n_604) );
A2O1A1Ixp33_ASAP7_75t_L g605 ( .A1(n_590), .A2(n_536), .B(n_558), .C(n_523), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_575), .B(n_545), .Y(n_606) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_566), .B(n_558), .Y(n_607) );
OA22x2_ASAP7_75t_L g608 ( .A1(n_567), .A2(n_541), .B1(n_523), .B2(n_536), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_581), .B(n_553), .Y(n_609) );
AOI211xp5_ASAP7_75t_L g610 ( .A1(n_577), .A2(n_539), .B(n_533), .C(n_535), .Y(n_610) );
XOR2x2_ASAP7_75t_L g611 ( .A(n_560), .B(n_300), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_580), .B(n_535), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_590), .A2(n_520), .B1(n_516), .B2(n_193), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_569), .Y(n_614) );
XNOR2x1_ASAP7_75t_L g615 ( .A(n_608), .B(n_611), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_595), .Y(n_616) );
NOR3xp33_ASAP7_75t_L g617 ( .A(n_594), .B(n_571), .C(n_591), .Y(n_617) );
AOI21xp33_ASAP7_75t_SL g618 ( .A1(n_602), .A2(n_579), .B(n_566), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_610), .A2(n_583), .B1(n_570), .B2(n_587), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_607), .A2(n_587), .B1(n_576), .B2(n_561), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g621 ( .A1(n_598), .A2(n_584), .B1(n_563), .B2(n_573), .C(n_571), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_605), .B(n_572), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_597), .B(n_586), .Y(n_623) );
AOI221xp5_ASAP7_75t_L g624 ( .A1(n_599), .A2(n_603), .B1(n_604), .B2(n_609), .C(n_601), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_600), .B(n_589), .Y(n_625) );
AOI21xp33_ASAP7_75t_L g626 ( .A1(n_613), .A2(n_593), .B(n_520), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_596), .A2(n_516), .B1(n_265), .B2(n_162), .Y(n_627) );
OAI22x1_ASAP7_75t_L g628 ( .A1(n_622), .A2(n_596), .B1(n_614), .B2(n_606), .Y(n_628) );
OAI311xp33_ASAP7_75t_L g629 ( .A1(n_624), .A2(n_612), .A3(n_229), .B1(n_169), .C1(n_162), .Y(n_629) );
NAND2x1_ASAP7_75t_L g630 ( .A(n_620), .B(n_619), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_618), .B(n_165), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_615), .A2(n_278), .B(n_283), .Y(n_632) );
AOI221x1_ASAP7_75t_L g633 ( .A1(n_617), .A2(n_162), .B1(n_166), .B2(n_168), .C(n_173), .Y(n_633) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_621), .A2(n_162), .B1(n_173), .B2(n_231), .C(n_241), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_630), .B(n_625), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_628), .B(n_616), .Y(n_636) );
AOI322xp5_ASAP7_75t_L g637 ( .A1(n_634), .A2(n_623), .A3(n_626), .B1(n_627), .B2(n_222), .C1(n_234), .C2(n_236), .Y(n_637) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_632), .A2(n_278), .B(n_264), .Y(n_638) );
INVxp67_ASAP7_75t_L g639 ( .A(n_635), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_636), .A2(n_631), .B1(n_629), .B2(n_633), .Y(n_640) );
NAND3xp33_ASAP7_75t_SL g641 ( .A(n_637), .B(n_638), .C(n_169), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_639), .B(n_278), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_640), .A2(n_222), .B1(n_234), .B2(n_236), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_643), .A2(n_641), .B1(n_162), .B2(n_222), .Y(n_644) );
OAI22x1_ASAP7_75t_L g645 ( .A1(n_644), .A2(n_642), .B1(n_194), .B2(n_228), .Y(n_645) );
NAND3xp33_ASAP7_75t_L g646 ( .A(n_645), .B(n_283), .C(n_234), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_646), .A2(n_194), .B1(n_234), .B2(n_236), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_647), .A2(n_283), .B(n_236), .Y(n_648) );
endmodule