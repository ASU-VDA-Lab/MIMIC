module fake_netlist_6_1692_n_1272 (n_52, n_1, n_91, n_326, n_256, n_209, n_63, n_223, n_278, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_56, n_119, n_235, n_147, n_191, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_53, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_231, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_317, n_149, n_90, n_24, n_54, n_328, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_315, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_332, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1272);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_231;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_317;
input n_149;
input n_90;
input n_24;
input n_54;
input n_328;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_332;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1272;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_509;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_447;
wire n_1172;
wire n_852;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_713;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_606;
wire n_818;
wire n_1123;
wire n_513;
wire n_645;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1068;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_354;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_487;
wire n_1107;
wire n_1014;
wire n_882;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_694;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_615;
wire n_1249;
wire n_1127;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1035;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_526;
wire n_1183;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_912;
wire n_745;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_819;
wire n_767;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_505;
wire n_537;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1224;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1267;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_385;
wire n_858;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_456;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1225;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_548;
wire n_833;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_569;
wire n_737;
wire n_1235;
wire n_1229;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_1047;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_855;
wire n_591;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1217;
wire n_751;
wire n_749;
wire n_969;
wire n_988;
wire n_1065;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1205;
wire n_1258;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_802;
wire n_561;
wire n_980;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_670;
wire n_1089;
wire n_1242;
wire n_681;
wire n_1226;
wire n_412;
wire n_640;
wire n_965;
wire n_339;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

INVx1_ASAP7_75t_L g334 ( 
.A(n_106),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_101),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_235),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_331),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_104),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_138),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_307),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_260),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_261),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_2),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_108),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_124),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_161),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_187),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_177),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_162),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_188),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_180),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_267),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_230),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_91),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_139),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_151),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_47),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_195),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_301),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_327),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_258),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_268),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_125),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_93),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_100),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_202),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_6),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_291),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_299),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_33),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_70),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_322),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_319),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_150),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_237),
.Y(n_375)
);

NOR2xp67_ASAP7_75t_L g376 ( 
.A(n_67),
.B(n_234),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_110),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_257),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_217),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_30),
.Y(n_380)
);

BUFx10_ASAP7_75t_L g381 ( 
.A(n_227),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_62),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_4),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_87),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_302),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_326),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_282),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_311),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_317),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_148),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_194),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_216),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_278),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_34),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_231),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_269),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_163),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_131),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_318),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_300),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_156),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_28),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_233),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_212),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_173),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_309),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_49),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_201),
.Y(n_408)
);

BUFx10_ASAP7_75t_L g409 ( 
.A(n_273),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_213),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_244),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_240),
.Y(n_412)
);

INVx2_ASAP7_75t_SL g413 ( 
.A(n_256),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_102),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_164),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_60),
.Y(n_416)
);

BUFx5_ASAP7_75t_L g417 ( 
.A(n_182),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_99),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_62),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_43),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_211),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_262),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_281),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_255),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_118),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_60),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_297),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_169),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_21),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_51),
.B(n_170),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_22),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_178),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_189),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_127),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_250),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_109),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_252),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_88),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_218),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_114),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_251),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_328),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_214),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_315),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_88),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_290),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_90),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_37),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_12),
.B(n_320),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_31),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_253),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_313),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_226),
.Y(n_453)
);

BUFx10_ASAP7_75t_L g454 ( 
.A(n_176),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_333),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_306),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_288),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_47),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_229),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_103),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_236),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_275),
.B(n_133),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_296),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_287),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_8),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_280),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_168),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_221),
.Y(n_468)
);

CKINVDCx14_ASAP7_75t_R g469 ( 
.A(n_285),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_154),
.Y(n_470)
);

BUFx10_ASAP7_75t_L g471 ( 
.A(n_87),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_207),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_122),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_12),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_314),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_325),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_149),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_198),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_165),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_44),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_228),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_332),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_243),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_83),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_18),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_200),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_50),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_107),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_279),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_51),
.Y(n_490)
);

BUFx5_ASAP7_75t_L g491 ( 
.A(n_57),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_196),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_79),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_2),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_310),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_81),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_117),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_271),
.Y(n_498)
);

NOR2xp67_ASAP7_75t_L g499 ( 
.A(n_175),
.B(n_242),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_491),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_491),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_379),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_335),
.B(n_0),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_379),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_364),
.Y(n_505)
);

OA21x2_ASAP7_75t_L g506 ( 
.A1(n_334),
.A2(n_0),
.B(n_1),
.Y(n_506)
);

BUFx8_ASAP7_75t_L g507 ( 
.A(n_352),
.Y(n_507)
);

AND2x6_ASAP7_75t_L g508 ( 
.A(n_379),
.B(n_105),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_491),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_422),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_363),
.B(n_435),
.Y(n_511)
);

AOI22x1_ASAP7_75t_SL g512 ( 
.A1(n_394),
.A2(n_4),
.B1(n_1),
.B2(n_3),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_369),
.B(n_3),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_491),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_491),
.Y(n_515)
);

CKINVDCx11_ASAP7_75t_R g516 ( 
.A(n_471),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_364),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_443),
.B(n_5),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_364),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_365),
.B(n_5),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_491),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_367),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_354),
.Y(n_523)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_422),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_422),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_370),
.Y(n_526)
);

INVx4_ASAP7_75t_L g527 ( 
.A(n_446),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_382),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_469),
.B(n_6),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_413),
.B(n_423),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_419),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_347),
.B(n_7),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_446),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_446),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_373),
.B(n_7),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g536 ( 
.A(n_447),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_380),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_471),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_378),
.B(n_8),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_384),
.Y(n_540)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_489),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_407),
.Y(n_542)
);

CKINVDCx6p67_ASAP7_75t_R g543 ( 
.A(n_392),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_417),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_403),
.B(n_9),
.Y(n_545)
);

BUFx12f_ASAP7_75t_L g546 ( 
.A(n_381),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_337),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_434),
.B(n_9),
.Y(n_548)
);

OA21x2_ASAP7_75t_L g549 ( 
.A1(n_338),
.A2(n_10),
.B(n_11),
.Y(n_549)
);

INVx4_ASAP7_75t_L g550 ( 
.A(n_489),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_442),
.A2(n_13),
.B1(n_10),
.B2(n_11),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_429),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_489),
.Y(n_553)
);

OA21x2_ASAP7_75t_L g554 ( 
.A1(n_341),
.A2(n_13),
.B(n_14),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_361),
.B(n_14),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_438),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_355),
.B(n_15),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_468),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_412),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_381),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_409),
.Y(n_561)
);

INVx5_ASAP7_75t_L g562 ( 
.A(n_409),
.Y(n_562)
);

BUFx8_ASAP7_75t_L g563 ( 
.A(n_430),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_454),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_480),
.Y(n_565)
);

INVx5_ASAP7_75t_L g566 ( 
.A(n_454),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_343),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_490),
.Y(n_568)
);

AOI22x1_ASAP7_75t_SL g569 ( 
.A1(n_416),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_415),
.B(n_16),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_355),
.B(n_17),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_357),
.Y(n_572)
);

INVx6_ASAP7_75t_L g573 ( 
.A(n_417),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_SL g574 ( 
.A(n_376),
.B(n_19),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_418),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_408),
.B(n_19),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_346),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_344),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_432),
.Y(n_579)
);

BUFx8_ASAP7_75t_L g580 ( 
.A(n_417),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_444),
.B(n_20),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_371),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_501),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_502),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_502),
.Y(n_585)
);

AOI21x1_ASAP7_75t_L g586 ( 
.A1(n_500),
.A2(n_348),
.B(n_345),
.Y(n_586)
);

INVx5_ASAP7_75t_L g587 ( 
.A(n_508),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_516),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_502),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_509),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_530),
.B(n_408),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_562),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_515),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_521),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_562),
.B(n_342),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_504),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_562),
.B(n_342),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_514),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_511),
.B(n_485),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_504),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_510),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_510),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_566),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_508),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_547),
.B(n_577),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_525),
.Y(n_606)
);

INVxp33_ASAP7_75t_L g607 ( 
.A(n_536),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_525),
.Y(n_608)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_508),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_525),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_533),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_572),
.B(n_459),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_533),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_566),
.B(n_475),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_533),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_534),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_566),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_513),
.B(n_377),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_534),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_558),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_561),
.B(n_377),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_561),
.B(n_564),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_553),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_559),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_564),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_505),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_559),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_505),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_558),
.B(n_495),
.Y(n_629)
);

AOI21x1_ASAP7_75t_L g630 ( 
.A1(n_544),
.A2(n_351),
.B(n_350),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_529),
.B(n_449),
.Y(n_631)
);

NAND3xp33_ASAP7_75t_L g632 ( 
.A(n_591),
.B(n_503),
.C(n_518),
.Y(n_632)
);

BUFx2_ASAP7_75t_L g633 ( 
.A(n_620),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_624),
.Y(n_634)
);

NOR3xp33_ASAP7_75t_L g635 ( 
.A(n_618),
.B(n_520),
.C(n_557),
.Y(n_635)
);

NOR3xp33_ASAP7_75t_L g636 ( 
.A(n_631),
.B(n_576),
.C(n_571),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_607),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_625),
.B(n_574),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_620),
.Y(n_639)
);

INVx8_ASAP7_75t_L g640 ( 
.A(n_599),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_605),
.B(n_543),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_625),
.B(n_567),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_627),
.B(n_612),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_621),
.B(n_560),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_601),
.B(n_524),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_622),
.B(n_563),
.Y(n_646)
);

INVxp67_ASAP7_75t_L g647 ( 
.A(n_599),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_592),
.B(n_538),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_601),
.B(n_524),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_592),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_604),
.A2(n_581),
.B1(n_570),
.B2(n_548),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_629),
.B(n_558),
.Y(n_652)
);

NOR3xp33_ASAP7_75t_L g653 ( 
.A(n_595),
.B(n_555),
.C(n_532),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_614),
.B(n_535),
.Y(n_654)
);

NAND3xp33_ASAP7_75t_SL g655 ( 
.A(n_597),
.B(n_551),
.C(n_545),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_598),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_584),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_584),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_606),
.B(n_527),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_603),
.B(n_563),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_604),
.A2(n_339),
.B1(n_340),
.B2(n_336),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_608),
.B(n_541),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_603),
.Y(n_663)
);

A2O1A1Ixp33_ASAP7_75t_L g664 ( 
.A1(n_583),
.A2(n_539),
.B(n_581),
.C(n_570),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_611),
.B(n_613),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_617),
.B(n_507),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_589),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_617),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_610),
.B(n_546),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_589),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_587),
.B(n_535),
.Y(n_671)
);

BUFx6f_ASAP7_75t_SL g672 ( 
.A(n_628),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_616),
.B(n_541),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_587),
.B(n_368),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_590),
.B(n_575),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_596),
.Y(n_676)
);

NOR3xp33_ASAP7_75t_L g677 ( 
.A(n_626),
.B(n_449),
.C(n_485),
.Y(n_677)
);

BUFx12f_ASAP7_75t_SL g678 ( 
.A(n_588),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_590),
.B(n_575),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_585),
.Y(n_680)
);

AOI221xp5_ASAP7_75t_L g681 ( 
.A1(n_626),
.A2(n_494),
.B1(n_487),
.B2(n_556),
.C(n_540),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_596),
.B(n_550),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_587),
.B(n_393),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_600),
.B(n_550),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_593),
.B(n_579),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_604),
.A2(n_549),
.B1(n_554),
.B2(n_506),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_602),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_594),
.B(n_579),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_615),
.B(n_517),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_594),
.B(n_579),
.Y(n_690)
);

AO22x1_ASAP7_75t_L g691 ( 
.A1(n_636),
.A2(n_402),
.B1(n_420),
.B2(n_383),
.Y(n_691)
);

A2O1A1Ixp33_ASAP7_75t_L g692 ( 
.A1(n_632),
.A2(n_499),
.B(n_411),
.C(n_462),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_651),
.B(n_609),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_689),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_647),
.B(n_404),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_675),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_SL g697 ( 
.A1(n_640),
.A2(n_569),
.B1(n_512),
.B2(n_467),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_639),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_654),
.B(n_619),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_661),
.A2(n_421),
.B1(n_411),
.B2(n_582),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_656),
.B(n_585),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_665),
.A2(n_366),
.B(n_362),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_633),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_679),
.Y(n_704)
);

OAI21x1_ASAP7_75t_L g705 ( 
.A1(n_686),
.A2(n_630),
.B(n_586),
.Y(n_705)
);

A2O1A1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_635),
.A2(n_375),
.B(n_387),
.C(n_372),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_653),
.A2(n_640),
.B1(n_683),
.B2(n_674),
.Y(n_707)
);

NAND2xp33_ASAP7_75t_L g708 ( 
.A(n_640),
.B(n_508),
.Y(n_708)
);

OAI21x1_ASAP7_75t_L g709 ( 
.A1(n_634),
.A2(n_630),
.B(n_586),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_681),
.B(n_349),
.Y(n_710)
);

O2A1O1Ixp5_ASAP7_75t_L g711 ( 
.A1(n_638),
.A2(n_578),
.B(n_397),
.C(n_398),
.Y(n_711)
);

OA22x2_ASAP7_75t_L g712 ( 
.A1(n_642),
.A2(n_431),
.B1(n_445),
.B2(n_426),
.Y(n_712)
);

O2A1O1Ixp33_ASAP7_75t_L g713 ( 
.A1(n_677),
.A2(n_526),
.B(n_552),
.C(n_522),
.Y(n_713)
);

BUFx4f_ASAP7_75t_L g714 ( 
.A(n_648),
.Y(n_714)
);

BUFx12f_ASAP7_75t_L g715 ( 
.A(n_680),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_657),
.B(n_623),
.Y(n_716)
);

NOR2x1_ASAP7_75t_L g717 ( 
.A(n_641),
.B(n_414),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_637),
.B(n_448),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_644),
.B(n_450),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_655),
.A2(n_549),
.B1(n_554),
.B2(n_506),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_658),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_685),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_667),
.Y(n_723)
);

O2A1O1Ixp33_ASAP7_75t_L g724 ( 
.A1(n_688),
.A2(n_568),
.B(n_565),
.C(n_542),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_670),
.B(n_676),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_687),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_652),
.B(n_650),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_690),
.A2(n_428),
.B(n_425),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_645),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_649),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_659),
.A2(n_437),
.B(n_433),
.Y(n_731)
);

A2O1A1Ixp33_ASAP7_75t_L g732 ( 
.A1(n_682),
.A2(n_684),
.B(n_439),
.C(n_440),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_663),
.B(n_537),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_662),
.B(n_673),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_668),
.B(n_537),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_SL g736 ( 
.A(n_678),
.B(n_672),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_646),
.A2(n_452),
.B(n_451),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_669),
.A2(n_455),
.B(n_453),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_660),
.B(n_458),
.Y(n_739)
);

A2O1A1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_666),
.A2(n_472),
.B(n_473),
.C(n_456),
.Y(n_740)
);

O2A1O1Ixp33_ASAP7_75t_SL g741 ( 
.A1(n_672),
.A2(n_477),
.B(n_478),
.C(n_476),
.Y(n_741)
);

BUFx4f_ASAP7_75t_L g742 ( 
.A(n_640),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_643),
.A2(n_497),
.B(n_356),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_632),
.B(n_465),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_643),
.A2(n_358),
.B(n_353),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_636),
.A2(n_360),
.B1(n_374),
.B2(n_359),
.Y(n_746)
);

OR2x2_ASAP7_75t_L g747 ( 
.A(n_637),
.B(n_542),
.Y(n_747)
);

NOR2x1_ASAP7_75t_L g748 ( 
.A(n_641),
.B(n_519),
.Y(n_748)
);

INVx1_ASAP7_75t_SL g749 ( 
.A(n_637),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_689),
.Y(n_750)
);

A2O1A1Ixp33_ASAP7_75t_L g751 ( 
.A1(n_632),
.A2(n_386),
.B(n_388),
.C(n_385),
.Y(n_751)
);

BUFx4f_ASAP7_75t_L g752 ( 
.A(n_640),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_632),
.B(n_389),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_632),
.B(n_474),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_643),
.A2(n_391),
.B(n_390),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_636),
.A2(n_396),
.B1(n_399),
.B2(n_395),
.Y(n_756)
);

OAI21xp5_ASAP7_75t_L g757 ( 
.A1(n_664),
.A2(n_401),
.B(n_400),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_643),
.A2(n_406),
.B(n_405),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_639),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_639),
.B(n_528),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_689),
.Y(n_761)
);

O2A1O1Ixp5_ASAP7_75t_L g762 ( 
.A1(n_671),
.A2(n_531),
.B(n_523),
.C(n_580),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_643),
.A2(n_424),
.B(n_410),
.Y(n_763)
);

O2A1O1Ixp33_ASAP7_75t_L g764 ( 
.A1(n_647),
.A2(n_523),
.B(n_580),
.C(n_436),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_637),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_643),
.A2(n_441),
.B(n_427),
.Y(n_766)
);

O2A1O1Ixp33_ASAP7_75t_L g767 ( 
.A1(n_647),
.A2(n_460),
.B(n_461),
.C(n_457),
.Y(n_767)
);

A2O1A1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_632),
.A2(n_464),
.B(n_466),
.C(n_463),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_651),
.B(n_470),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_637),
.B(n_484),
.Y(n_770)
);

BUFx4f_ASAP7_75t_L g771 ( 
.A(n_640),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_651),
.B(n_479),
.Y(n_772)
);

A2O1A1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_632),
.A2(n_482),
.B(n_483),
.C(n_481),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_L g774 ( 
.A1(n_632),
.A2(n_488),
.B1(n_492),
.B2(n_486),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_651),
.B(n_498),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_696),
.B(n_573),
.Y(n_776)
);

OAI21xp5_ASAP7_75t_L g777 ( 
.A1(n_693),
.A2(n_496),
.B(n_493),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_703),
.Y(n_778)
);

BUFx8_ASAP7_75t_L g779 ( 
.A(n_715),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_704),
.B(n_23),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_695),
.B(n_512),
.Y(n_781)
);

OAI21x1_ASAP7_75t_SL g782 ( 
.A1(n_764),
.A2(n_569),
.B(n_112),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_L g783 ( 
.A1(n_692),
.A2(n_113),
.B(n_111),
.Y(n_783)
);

OA21x2_ASAP7_75t_L g784 ( 
.A1(n_709),
.A2(n_116),
.B(n_115),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_698),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_722),
.B(n_729),
.Y(n_786)
);

INVxp67_ASAP7_75t_L g787 ( 
.A(n_765),
.Y(n_787)
);

NAND2x1p5_ASAP7_75t_L g788 ( 
.A(n_752),
.B(n_119),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_734),
.A2(n_121),
.B(n_120),
.Y(n_789)
);

A2O1A1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_744),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_752),
.B(n_771),
.Y(n_791)
);

AOI211x1_ASAP7_75t_L g792 ( 
.A1(n_691),
.A2(n_26),
.B(n_24),
.C(n_25),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_708),
.A2(n_126),
.B(n_123),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_730),
.B(n_26),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_699),
.A2(n_129),
.B(n_128),
.Y(n_795)
);

AO31x2_ASAP7_75t_L g796 ( 
.A1(n_706),
.A2(n_29),
.A3(n_27),
.B(n_28),
.Y(n_796)
);

AO31x2_ASAP7_75t_L g797 ( 
.A1(n_732),
.A2(n_30),
.A3(n_27),
.B(n_29),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_749),
.Y(n_798)
);

BUFx10_ASAP7_75t_L g799 ( 
.A(n_718),
.Y(n_799)
);

INVx4_ASAP7_75t_L g800 ( 
.A(n_703),
.Y(n_800)
);

OAI21x1_ASAP7_75t_L g801 ( 
.A1(n_726),
.A2(n_725),
.B(n_716),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_719),
.B(n_31),
.Y(n_802)
);

BUFx2_ASAP7_75t_L g803 ( 
.A(n_747),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_770),
.B(n_733),
.Y(n_804)
);

OR2x6_ASAP7_75t_L g805 ( 
.A(n_698),
.B(n_32),
.Y(n_805)
);

OAI21xp5_ASAP7_75t_L g806 ( 
.A1(n_754),
.A2(n_132),
.B(n_130),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_721),
.Y(n_807)
);

OAI21xp5_ASAP7_75t_L g808 ( 
.A1(n_751),
.A2(n_135),
.B(n_134),
.Y(n_808)
);

INVx1_ASAP7_75t_SL g809 ( 
.A(n_735),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_723),
.Y(n_810)
);

OAI21xp5_ASAP7_75t_L g811 ( 
.A1(n_768),
.A2(n_137),
.B(n_136),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_714),
.B(n_727),
.Y(n_812)
);

INVx4_ASAP7_75t_L g813 ( 
.A(n_742),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_769),
.A2(n_141),
.B(n_140),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_L g815 ( 
.A1(n_707),
.A2(n_143),
.B1(n_144),
.B2(n_142),
.Y(n_815)
);

O2A1O1Ixp5_ASAP7_75t_L g816 ( 
.A1(n_753),
.A2(n_146),
.B(n_147),
.C(n_145),
.Y(n_816)
);

INVx4_ASAP7_75t_L g817 ( 
.A(n_771),
.Y(n_817)
);

AO31x2_ASAP7_75t_L g818 ( 
.A1(n_773),
.A2(n_36),
.A3(n_34),
.B(n_35),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_717),
.B(n_35),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_746),
.B(n_756),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_694),
.B(n_36),
.Y(n_821)
);

NAND3xp33_ASAP7_75t_L g822 ( 
.A(n_700),
.B(n_38),
.C(n_39),
.Y(n_822)
);

OAI21xp5_ASAP7_75t_L g823 ( 
.A1(n_720),
.A2(n_153),
.B(n_152),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_772),
.B(n_155),
.Y(n_824)
);

OAI21xp5_ASAP7_75t_L g825 ( 
.A1(n_775),
.A2(n_158),
.B(n_157),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_701),
.A2(n_160),
.B(n_159),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_760),
.Y(n_827)
);

NOR2xp67_ASAP7_75t_L g828 ( 
.A(n_774),
.B(n_166),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_759),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_750),
.B(n_39),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_761),
.B(n_40),
.Y(n_831)
);

AOI21x1_ASAP7_75t_L g832 ( 
.A1(n_743),
.A2(n_171),
.B(n_167),
.Y(n_832)
);

OAI21xp33_ASAP7_75t_L g833 ( 
.A1(n_739),
.A2(n_40),
.B(n_41),
.Y(n_833)
);

OAI21x1_ASAP7_75t_L g834 ( 
.A1(n_762),
.A2(n_174),
.B(n_172),
.Y(n_834)
);

A2O1A1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_767),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_835)
);

AO31x2_ASAP7_75t_L g836 ( 
.A1(n_728),
.A2(n_45),
.A3(n_42),
.B(n_44),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_710),
.B(n_46),
.Y(n_837)
);

AOI221x1_ASAP7_75t_L g838 ( 
.A1(n_702),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.C(n_50),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_757),
.A2(n_181),
.B(n_179),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_712),
.A2(n_184),
.B1(n_185),
.B2(n_183),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_748),
.B(n_48),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_745),
.B(n_755),
.Y(n_842)
);

CKINVDCx6p67_ASAP7_75t_R g843 ( 
.A(n_759),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_758),
.A2(n_190),
.B(n_186),
.Y(n_844)
);

A2O1A1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_711),
.A2(n_52),
.B(n_53),
.C(n_54),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_741),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_763),
.B(n_52),
.Y(n_847)
);

CKINVDCx6p67_ASAP7_75t_R g848 ( 
.A(n_736),
.Y(n_848)
);

OA21x2_ASAP7_75t_L g849 ( 
.A1(n_731),
.A2(n_192),
.B(n_191),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_766),
.A2(n_247),
.B1(n_330),
.B2(n_329),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_SL g851 ( 
.A1(n_740),
.A2(n_197),
.B(n_193),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_737),
.B(n_738),
.Y(n_852)
);

AOI31xp67_ASAP7_75t_L g853 ( 
.A1(n_724),
.A2(n_248),
.A3(n_324),
.B(n_323),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_713),
.Y(n_854)
);

OAI21x1_ASAP7_75t_L g855 ( 
.A1(n_697),
.A2(n_321),
.B(n_203),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_749),
.B(n_55),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_698),
.B(n_199),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_749),
.B(n_55),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_734),
.A2(n_205),
.B(n_204),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_705),
.A2(n_208),
.B(n_206),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_698),
.Y(n_861)
);

NOR2xp67_ASAP7_75t_L g862 ( 
.A(n_765),
.B(n_209),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_752),
.B(n_210),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_696),
.B(n_56),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_696),
.B(n_56),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_696),
.B(n_57),
.Y(n_866)
);

AO31x2_ASAP7_75t_L g867 ( 
.A1(n_692),
.A2(n_58),
.A3(n_59),
.B(n_61),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_749),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_695),
.B(n_58),
.Y(n_869)
);

NOR3xp33_ASAP7_75t_L g870 ( 
.A(n_700),
.B(n_59),
.C(n_61),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_705),
.A2(n_219),
.B(n_215),
.Y(n_871)
);

INVx5_ASAP7_75t_L g872 ( 
.A(n_715),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_734),
.A2(n_259),
.B(n_316),
.Y(n_873)
);

AO31x2_ASAP7_75t_L g874 ( 
.A1(n_692),
.A2(n_63),
.A3(n_64),
.B(n_65),
.Y(n_874)
);

NAND2x1p5_ASAP7_75t_L g875 ( 
.A(n_752),
.B(n_220),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_698),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_752),
.B(n_222),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_696),
.B(n_63),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_696),
.B(n_64),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_696),
.B(n_65),
.Y(n_880)
);

A2O1A1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_744),
.A2(n_66),
.B(n_67),
.C(n_68),
.Y(n_881)
);

INVxp67_ASAP7_75t_SL g882 ( 
.A(n_693),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_698),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_696),
.B(n_66),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_734),
.A2(n_263),
.B(n_312),
.Y(n_885)
);

NOR2x1_ASAP7_75t_SL g886 ( 
.A(n_693),
.B(n_223),
.Y(n_886)
);

BUFx3_ASAP7_75t_L g887 ( 
.A(n_703),
.Y(n_887)
);

BUFx3_ASAP7_75t_L g888 ( 
.A(n_703),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_703),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_734),
.A2(n_254),
.B(n_308),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_696),
.B(n_68),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_786),
.Y(n_892)
);

CKINVDCx6p67_ASAP7_75t_R g893 ( 
.A(n_872),
.Y(n_893)
);

AOI221xp5_ASAP7_75t_L g894 ( 
.A1(n_781),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.C(n_72),
.Y(n_894)
);

AO21x2_ASAP7_75t_L g895 ( 
.A1(n_823),
.A2(n_264),
.B(n_305),
.Y(n_895)
);

OA21x2_ASAP7_75t_L g896 ( 
.A1(n_801),
.A2(n_249),
.B(n_304),
.Y(n_896)
);

OAI21xp5_ASAP7_75t_L g897 ( 
.A1(n_882),
.A2(n_246),
.B(n_303),
.Y(n_897)
);

NAND2x1p5_ASAP7_75t_L g898 ( 
.A(n_800),
.B(n_224),
.Y(n_898)
);

AO32x2_ASAP7_75t_L g899 ( 
.A1(n_840),
.A2(n_73),
.A3(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_899)
);

AO21x2_ASAP7_75t_L g900 ( 
.A1(n_839),
.A2(n_245),
.B(n_298),
.Y(n_900)
);

INVxp67_ASAP7_75t_SL g901 ( 
.A(n_798),
.Y(n_901)
);

CKINVDCx14_ASAP7_75t_R g902 ( 
.A(n_868),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_804),
.B(n_225),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_810),
.Y(n_904)
);

OAI22xp5_ASAP7_75t_L g905 ( 
.A1(n_820),
.A2(n_265),
.B1(n_295),
.B2(n_294),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_807),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_842),
.A2(n_241),
.B(n_293),
.Y(n_907)
);

AO21x2_ASAP7_75t_L g908 ( 
.A1(n_783),
.A2(n_239),
.B(n_292),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_869),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_780),
.Y(n_910)
);

BUFx12f_ASAP7_75t_L g911 ( 
.A(n_779),
.Y(n_911)
);

BUFx3_ASAP7_75t_L g912 ( 
.A(n_887),
.Y(n_912)
);

INVx5_ASAP7_75t_L g913 ( 
.A(n_785),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_864),
.Y(n_914)
);

INVx3_ASAP7_75t_SL g915 ( 
.A(n_848),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_802),
.A2(n_77),
.B(n_78),
.C(n_79),
.Y(n_916)
);

AOI22xp33_ASAP7_75t_L g917 ( 
.A1(n_870),
.A2(n_854),
.B1(n_777),
.B2(n_837),
.Y(n_917)
);

INVx8_ASAP7_75t_L g918 ( 
.A(n_872),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_865),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_866),
.Y(n_920)
);

BUFx2_ASAP7_75t_L g921 ( 
.A(n_787),
.Y(n_921)
);

OR2x2_ASAP7_75t_L g922 ( 
.A(n_778),
.B(n_77),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_L g923 ( 
.A1(n_794),
.A2(n_266),
.B(n_289),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_812),
.B(n_78),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_827),
.Y(n_925)
);

CKINVDCx16_ASAP7_75t_R g926 ( 
.A(n_888),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_878),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_879),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_880),
.A2(n_238),
.B(n_286),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_856),
.B(n_80),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_884),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_891),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_830),
.Y(n_933)
);

OAI22xp33_ASAP7_75t_L g934 ( 
.A1(n_822),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_934)
);

OA21x2_ASAP7_75t_L g935 ( 
.A1(n_860),
.A2(n_270),
.B(n_284),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_829),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_831),
.B(n_84),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_776),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_829),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_861),
.Y(n_940)
);

AOI221xp5_ASAP7_75t_L g941 ( 
.A1(n_833),
.A2(n_85),
.B1(n_86),
.B2(n_89),
.C(n_90),
.Y(n_941)
);

OAI22xp33_ASAP7_75t_L g942 ( 
.A1(n_821),
.A2(n_85),
.B1(n_86),
.B2(n_89),
.Y(n_942)
);

OA21x2_ASAP7_75t_L g943 ( 
.A1(n_871),
.A2(n_274),
.B(n_283),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_858),
.B(n_799),
.Y(n_944)
);

AOI22xp33_ASAP7_75t_SL g945 ( 
.A1(n_799),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_889),
.Y(n_946)
);

NOR2x1_ASAP7_75t_SL g947 ( 
.A(n_863),
.B(n_272),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_861),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_843),
.Y(n_949)
);

BUFx2_ASAP7_75t_R g950 ( 
.A(n_791),
.Y(n_950)
);

BUFx10_ASAP7_75t_L g951 ( 
.A(n_857),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_876),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_876),
.B(n_232),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_813),
.B(n_94),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_876),
.Y(n_955)
);

BUFx2_ASAP7_75t_L g956 ( 
.A(n_883),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_867),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_867),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_867),
.Y(n_959)
);

AOI22x1_ASAP7_75t_L g960 ( 
.A1(n_825),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_874),
.Y(n_961)
);

NAND2x1_ASAP7_75t_L g962 ( 
.A(n_817),
.B(n_276),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_857),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_872),
.B(n_277),
.Y(n_964)
);

INVx6_ASAP7_75t_SL g965 ( 
.A(n_805),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_779),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_874),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_855),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_862),
.B(n_96),
.Y(n_969)
);

OA21x2_ASAP7_75t_L g970 ( 
.A1(n_789),
.A2(n_98),
.B(n_808),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_782),
.Y(n_971)
);

CKINVDCx11_ASAP7_75t_R g972 ( 
.A(n_846),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_841),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_811),
.A2(n_828),
.B(n_806),
.Y(n_974)
);

INVxp67_ASAP7_75t_SL g975 ( 
.A(n_847),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_844),
.A2(n_819),
.B(n_790),
.C(n_881),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_797),
.Y(n_977)
);

NOR2x1_ASAP7_75t_SL g978 ( 
.A(n_877),
.B(n_815),
.Y(n_978)
);

BUFx2_ASAP7_75t_SL g979 ( 
.A(n_846),
.Y(n_979)
);

CKINVDCx11_ASAP7_75t_R g980 ( 
.A(n_852),
.Y(n_980)
);

AOI221xp5_ASAP7_75t_L g981 ( 
.A1(n_782),
.A2(n_792),
.B1(n_835),
.B2(n_845),
.C(n_890),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_788),
.B(n_875),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_L g983 ( 
.A1(n_859),
.A2(n_873),
.B1(n_885),
.B2(n_850),
.Y(n_983)
);

BUFx3_ASAP7_75t_L g984 ( 
.A(n_818),
.Y(n_984)
);

INVxp67_ASAP7_75t_L g985 ( 
.A(n_834),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_816),
.A2(n_814),
.B(n_795),
.C(n_793),
.Y(n_986)
);

BUFx2_ASAP7_75t_L g987 ( 
.A(n_818),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_796),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_826),
.A2(n_784),
.B(n_849),
.C(n_838),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_796),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_832),
.B(n_851),
.Y(n_991)
);

INVxp67_ASAP7_75t_L g992 ( 
.A(n_832),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_836),
.B(n_853),
.Y(n_993)
);

AOI22xp33_ASAP7_75t_L g994 ( 
.A1(n_836),
.A2(n_820),
.B1(n_869),
.B2(n_636),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_836),
.A2(n_882),
.B(n_823),
.Y(n_995)
);

NOR2x1_ASAP7_75t_SL g996 ( 
.A(n_824),
.B(n_842),
.Y(n_996)
);

OAI22xp33_ASAP7_75t_L g997 ( 
.A1(n_802),
.A2(n_661),
.B1(n_809),
.B2(n_632),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_786),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_786),
.B(n_804),
.Y(n_999)
);

CKINVDCx20_ASAP7_75t_R g1000 ( 
.A(n_868),
.Y(n_1000)
);

AO31x2_ASAP7_75t_L g1001 ( 
.A1(n_838),
.A2(n_886),
.A3(n_692),
.B(n_706),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_804),
.B(n_803),
.Y(n_1002)
);

AND2x2_ASAP7_75t_SL g1003 ( 
.A(n_970),
.B(n_994),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_913),
.Y(n_1004)
);

AOI22xp33_ASAP7_75t_SL g1005 ( 
.A1(n_960),
.A2(n_974),
.B1(n_970),
.B2(n_930),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_892),
.B(n_998),
.Y(n_1006)
);

NOR2x1_ASAP7_75t_SL g1007 ( 
.A(n_979),
.B(n_892),
.Y(n_1007)
);

CKINVDCx11_ASAP7_75t_R g1008 ( 
.A(n_911),
.Y(n_1008)
);

INVx2_ASAP7_75t_SL g1009 ( 
.A(n_912),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_913),
.Y(n_1010)
);

INVx11_ASAP7_75t_L g1011 ( 
.A(n_926),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_913),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_998),
.B(n_999),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_965),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_1002),
.B(n_944),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_906),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_924),
.B(n_963),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_904),
.Y(n_1018)
);

INVx2_ASAP7_75t_SL g1019 ( 
.A(n_946),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_963),
.B(n_952),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_933),
.B(n_973),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_910),
.B(n_914),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_1000),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_951),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_919),
.B(n_920),
.Y(n_1025)
);

HB1xp67_ASAP7_75t_L g1026 ( 
.A(n_901),
.Y(n_1026)
);

HB1xp67_ASAP7_75t_L g1027 ( 
.A(n_955),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_927),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_948),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_928),
.Y(n_1030)
);

OR2x2_ASAP7_75t_L g1031 ( 
.A(n_921),
.B(n_931),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_932),
.B(n_951),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_925),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_940),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_956),
.Y(n_1035)
);

NAND4xp25_ASAP7_75t_L g1036 ( 
.A(n_894),
.B(n_909),
.C(n_945),
.D(n_941),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_990),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_957),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_958),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_958),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_949),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_L g1042 ( 
.A(n_939),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_959),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_959),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_961),
.Y(n_1045)
);

OR2x6_ASAP7_75t_L g1046 ( 
.A(n_918),
.B(n_982),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_936),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_939),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_917),
.B(n_938),
.Y(n_1049)
);

INVx5_ASAP7_75t_L g1050 ( 
.A(n_939),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_967),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_977),
.Y(n_1052)
);

OR2x2_ASAP7_75t_L g1053 ( 
.A(n_937),
.B(n_997),
.Y(n_1053)
);

BUFx3_ASAP7_75t_L g1054 ( 
.A(n_918),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_988),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_902),
.B(n_954),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_984),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_962),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_965),
.Y(n_1059)
);

HB1xp67_ASAP7_75t_L g1060 ( 
.A(n_922),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_975),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_987),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_971),
.B(n_964),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_1001),
.Y(n_1064)
);

HB1xp67_ASAP7_75t_L g1065 ( 
.A(n_1001),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_899),
.Y(n_1066)
);

OAI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_960),
.A2(n_942),
.B1(n_934),
.B2(n_969),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_1001),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_968),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_980),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_899),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_947),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_947),
.Y(n_1073)
);

HB1xp67_ASAP7_75t_L g1074 ( 
.A(n_976),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_915),
.Y(n_1075)
);

INVx1_ASAP7_75t_SL g1076 ( 
.A(n_972),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_950),
.B(n_964),
.Y(n_1077)
);

OA21x2_ASAP7_75t_L g1078 ( 
.A1(n_995),
.A2(n_992),
.B(n_985),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_916),
.B(n_898),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_899),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_953),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_903),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_893),
.B(n_929),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_993),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_966),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_996),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_908),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_996),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_981),
.B(n_923),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_897),
.A2(n_905),
.B1(n_895),
.B2(n_900),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1006),
.B(n_978),
.Y(n_1091)
);

CKINVDCx20_ASAP7_75t_R g1092 ( 
.A(n_1023),
.Y(n_1092)
);

NAND2x1_ASAP7_75t_L g1093 ( 
.A(n_1058),
.B(n_983),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1006),
.B(n_978),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1015),
.B(n_935),
.Y(n_1095)
);

HB1xp67_ASAP7_75t_L g1096 ( 
.A(n_1062),
.Y(n_1096)
);

OR2x6_ASAP7_75t_L g1097 ( 
.A(n_1063),
.B(n_907),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1021),
.B(n_943),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1017),
.B(n_896),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1013),
.B(n_1074),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_1009),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_1057),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1013),
.B(n_1074),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1022),
.B(n_986),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_1063),
.Y(n_1105)
);

INVx1_ASAP7_75t_SL g1106 ( 
.A(n_1031),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1016),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_1057),
.Y(n_1108)
);

INVxp67_ASAP7_75t_L g1109 ( 
.A(n_1026),
.Y(n_1109)
);

INVx8_ASAP7_75t_L g1110 ( 
.A(n_1050),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1049),
.B(n_991),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1028),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1025),
.B(n_989),
.Y(n_1113)
);

AO221x2_ASAP7_75t_L g1114 ( 
.A1(n_1067),
.A2(n_1066),
.B1(n_1080),
.B2(n_1071),
.C(n_1049),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1089),
.B(n_1053),
.Y(n_1115)
);

INVx2_ASAP7_75t_SL g1116 ( 
.A(n_1011),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1060),
.B(n_1032),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1030),
.Y(n_1118)
);

BUFx2_ASAP7_75t_L g1119 ( 
.A(n_1029),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1038),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1039),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_1077),
.B(n_1033),
.Y(n_1122)
);

INVxp67_ASAP7_75t_R g1123 ( 
.A(n_1056),
.Y(n_1123)
);

AND2x4_ASAP7_75t_L g1124 ( 
.A(n_1020),
.B(n_1046),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1061),
.B(n_1082),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1040),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1043),
.Y(n_1127)
);

BUFx2_ASAP7_75t_SL g1128 ( 
.A(n_1023),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1044),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1029),
.B(n_1035),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_1054),
.B(n_1024),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1027),
.B(n_1018),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1045),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_1083),
.B(n_1034),
.Y(n_1134)
);

BUFx2_ASAP7_75t_L g1135 ( 
.A(n_1042),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_1019),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1082),
.B(n_1067),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_1041),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1051),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1052),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1005),
.B(n_1055),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1048),
.B(n_1047),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_1041),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_1054),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1037),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_1036),
.B(n_1081),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1114),
.B(n_1113),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1115),
.B(n_1007),
.Y(n_1148)
);

OR2x2_ASAP7_75t_L g1149 ( 
.A(n_1106),
.B(n_1084),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1115),
.B(n_1079),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1145),
.Y(n_1151)
);

OR2x2_ASAP7_75t_L g1152 ( 
.A(n_1106),
.B(n_1070),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1120),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1117),
.B(n_1134),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1146),
.B(n_1036),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1121),
.Y(n_1156)
);

NAND2x1p5_ASAP7_75t_L g1157 ( 
.A(n_1093),
.B(n_1088),
.Y(n_1157)
);

INVx1_ASAP7_75t_SL g1158 ( 
.A(n_1130),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1114),
.B(n_1064),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1114),
.B(n_1065),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1126),
.Y(n_1161)
);

NOR2x1_ASAP7_75t_L g1162 ( 
.A(n_1138),
.B(n_1086),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1127),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1098),
.B(n_1068),
.Y(n_1164)
);

OR2x2_ASAP7_75t_L g1165 ( 
.A(n_1111),
.B(n_1069),
.Y(n_1165)
);

OR2x2_ASAP7_75t_L g1166 ( 
.A(n_1111),
.B(n_1069),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1129),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1133),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1146),
.B(n_1005),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1095),
.B(n_1003),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1100),
.B(n_1103),
.Y(n_1171)
);

BUFx3_ASAP7_75t_L g1172 ( 
.A(n_1138),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1139),
.B(n_1003),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1100),
.B(n_1073),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1140),
.B(n_1078),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1103),
.B(n_1072),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1096),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1142),
.B(n_1004),
.Y(n_1178)
);

OR2x2_ASAP7_75t_L g1179 ( 
.A(n_1125),
.B(n_1076),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1125),
.B(n_1010),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_1137),
.B(n_1012),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1102),
.B(n_1087),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_1119),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1132),
.B(n_1012),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_1155),
.B(n_1150),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1177),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1154),
.B(n_1158),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1171),
.B(n_1091),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1153),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1156),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1180),
.B(n_1091),
.Y(n_1191)
);

OR2x2_ASAP7_75t_L g1192 ( 
.A(n_1170),
.B(n_1141),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1161),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1178),
.B(n_1122),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1165),
.B(n_1094),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1163),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1167),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1168),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_1182),
.B(n_1108),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1147),
.B(n_1123),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1173),
.B(n_1099),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1173),
.B(n_1135),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1166),
.B(n_1094),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1181),
.B(n_1109),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_1182),
.B(n_1175),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_1175),
.B(n_1097),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1181),
.B(n_1174),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1176),
.B(n_1109),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1155),
.B(n_1137),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1151),
.Y(n_1210)
);

OR2x2_ASAP7_75t_L g1211 ( 
.A(n_1205),
.B(n_1179),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1207),
.B(n_1169),
.Y(n_1212)
);

O2A1O1Ixp33_ASAP7_75t_SL g1213 ( 
.A1(n_1209),
.A2(n_1148),
.B(n_1185),
.C(n_1204),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1198),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_1185),
.B(n_1162),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1198),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1189),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1190),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1195),
.B(n_1183),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1193),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1203),
.B(n_1159),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1191),
.B(n_1160),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1188),
.B(n_1160),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1196),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1197),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1201),
.B(n_1164),
.Y(n_1226)
);

AOI221xp5_ASAP7_75t_L g1227 ( 
.A1(n_1208),
.A2(n_1184),
.B1(n_1112),
.B2(n_1118),
.C(n_1107),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1214),
.Y(n_1228)
);

OAI222xp33_ASAP7_75t_L g1229 ( 
.A1(n_1215),
.A2(n_1192),
.B1(n_1200),
.B2(n_1206),
.C1(n_1152),
.C2(n_1187),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1223),
.B(n_1222),
.Y(n_1230)
);

AOI211xp5_ASAP7_75t_L g1231 ( 
.A1(n_1213),
.A2(n_1076),
.B(n_1149),
.C(n_1210),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1216),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1221),
.B(n_1186),
.Y(n_1233)
);

AOI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1215),
.A2(n_1206),
.B1(n_1097),
.B2(n_1124),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1214),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1226),
.B(n_1206),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1212),
.A2(n_1227),
.B(n_1143),
.C(n_1172),
.Y(n_1237)
);

INVx1_ASAP7_75t_SL g1238 ( 
.A(n_1211),
.Y(n_1238)
);

OAI221xp5_ASAP7_75t_L g1239 ( 
.A1(n_1213),
.A2(n_1090),
.B1(n_1128),
.B2(n_1157),
.C(n_1143),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1236),
.Y(n_1240)
);

OAI32xp33_ASAP7_75t_L g1241 ( 
.A1(n_1239),
.A2(n_1219),
.A3(n_1217),
.B1(n_1220),
.B2(n_1225),
.Y(n_1241)
);

AOI211xp5_ASAP7_75t_L g1242 ( 
.A1(n_1239),
.A2(n_1237),
.B(n_1231),
.C(n_1229),
.Y(n_1242)
);

BUFx3_ASAP7_75t_L g1243 ( 
.A(n_1238),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1232),
.Y(n_1244)
);

AOI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1234),
.A2(n_1105),
.B1(n_1194),
.B2(n_1202),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1235),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1228),
.Y(n_1247)
);

OAI21xp33_ASAP7_75t_L g1248 ( 
.A1(n_1242),
.A2(n_1230),
.B(n_1233),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1243),
.B(n_1230),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1241),
.A2(n_1233),
.B(n_1224),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1245),
.A2(n_1104),
.B(n_1218),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1244),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1252),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1248),
.B(n_1240),
.Y(n_1254)
);

NAND3xp33_ASAP7_75t_L g1255 ( 
.A(n_1251),
.B(n_1245),
.C(n_1246),
.Y(n_1255)
);

OAI21xp5_ASAP7_75t_SL g1256 ( 
.A1(n_1250),
.A2(n_1090),
.B(n_1075),
.Y(n_1256)
);

NOR2x1_ASAP7_75t_L g1257 ( 
.A(n_1249),
.B(n_1092),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1248),
.A2(n_1097),
.B1(n_1247),
.B2(n_1199),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1253),
.Y(n_1259)
);

NOR2x1_ASAP7_75t_L g1260 ( 
.A(n_1257),
.B(n_1092),
.Y(n_1260)
);

NOR2x1_ASAP7_75t_L g1261 ( 
.A(n_1255),
.B(n_1254),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1261),
.B(n_1256),
.Y(n_1262)
);

NOR2x1_ASAP7_75t_L g1263 ( 
.A(n_1260),
.B(n_1101),
.Y(n_1263)
);

NOR2x1_ASAP7_75t_L g1264 ( 
.A(n_1263),
.B(n_1259),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1264),
.A2(n_1262),
.B(n_1085),
.Y(n_1265)
);

OAI22x1_ASAP7_75t_L g1266 ( 
.A1(n_1265),
.A2(n_1085),
.B1(n_1014),
.B2(n_1059),
.Y(n_1266)
);

AOI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1266),
.A2(n_1258),
.B1(n_1008),
.B2(n_1116),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1267),
.A2(n_1144),
.B(n_1101),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1268),
.A2(n_1008),
.B(n_1136),
.Y(n_1269)
);

AOI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1269),
.A2(n_1136),
.B1(n_1131),
.B2(n_1172),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_SL g1271 ( 
.A(n_1270),
.B(n_1050),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1271),
.A2(n_1010),
.B(n_1110),
.Y(n_1272)
);


endmodule