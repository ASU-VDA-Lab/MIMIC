module fake_jpeg_4163_n_344 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_20),
.Y(n_51)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_42),
.B1(n_44),
.B2(n_46),
.Y(n_59)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_51),
.B(n_58),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_38),
.B(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_54),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_27),
.B1(n_35),
.B2(n_19),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_53),
.A2(n_20),
.B1(n_28),
.B2(n_31),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_48),
.A2(n_35),
.B1(n_27),
.B2(n_19),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_17),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_63),
.Y(n_75)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_67),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_70),
.Y(n_87)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_78),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_65),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_76),
.Y(n_104)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_80),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_35),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_84),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_63),
.A2(n_49),
.B1(n_27),
.B2(n_47),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_90),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_41),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_85),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_69),
.B(n_45),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_96),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_71),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_89),
.Y(n_125)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_54),
.A2(n_40),
.B1(n_39),
.B2(n_46),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_91),
.A2(n_95),
.B1(n_18),
.B2(n_21),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_69),
.A2(n_46),
.B1(n_22),
.B2(n_28),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_41),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_41),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_99),
.C(n_101),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_57),
.B(n_45),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_100),
.A2(n_22),
.B1(n_21),
.B2(n_31),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_59),
.B(n_45),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_56),
.B(n_45),
.Y(n_102)
);

MAJx2_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_37),
.C(n_33),
.Y(n_127)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_106),
.Y(n_132)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_84),
.A2(n_30),
.B(n_23),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_108),
.A2(n_130),
.B(n_34),
.Y(n_160)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_114),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_115),
.B(n_123),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_85),
.A2(n_44),
.B1(n_42),
.B2(n_49),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_116),
.A2(n_128),
.B1(n_78),
.B2(n_93),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_73),
.A2(n_44),
.B1(n_42),
.B2(n_30),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_122),
.A2(n_72),
.B1(n_100),
.B2(n_79),
.Y(n_139)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_76),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_124),
.B(n_126),
.Y(n_153)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_74),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_101),
.A2(n_56),
.B1(n_34),
.B2(n_30),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_129),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_34),
.B(n_23),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_131),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_133),
.A2(n_143),
.B1(n_148),
.B2(n_118),
.Y(n_177)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_137),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_97),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_138),
.Y(n_166)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_139),
.A2(n_111),
.B1(n_129),
.B2(n_131),
.Y(n_165)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_149),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

INVxp67_ASAP7_75t_SL g190 ( 
.A(n_141),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_97),
.B1(n_88),
.B2(n_102),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_117),
.A2(n_99),
.B(n_96),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_146),
.B(n_103),
.Y(n_178)
);

OA21x2_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_98),
.B(n_83),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_110),
.A2(n_97),
.B1(n_89),
.B2(n_90),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_151),
.B(n_127),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_104),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_152),
.Y(n_162)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_158),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_114),
.Y(n_155)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_156),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_108),
.Y(n_157)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_94),
.C(n_80),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_125),
.C(n_33),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_160),
.A2(n_107),
.B(n_111),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_33),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_135),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_185),
.C(n_137),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_164),
.A2(n_175),
.B(n_134),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_165),
.B(n_182),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_161),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_168),
.B(n_33),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_132),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_176),
.Y(n_205)
);

MAJx2_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_112),
.C(n_123),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_171),
.B(n_26),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_149),
.A2(n_112),
.B(n_106),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_146),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_178),
.A2(n_180),
.B(n_183),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_181),
.Y(n_204)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_142),
.A2(n_118),
.B(n_23),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_133),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_184),
.B(n_187),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_139),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_189),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_143),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_191),
.Y(n_206)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_141),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_192),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_151),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_193),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_154),
.A2(n_119),
.B1(n_18),
.B2(n_29),
.Y(n_194)
);

OAI22x1_ASAP7_75t_L g207 ( 
.A1(n_194),
.A2(n_26),
.B1(n_171),
.B2(n_183),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_195),
.A2(n_199),
.B(n_208),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_186),
.A2(n_147),
.B1(n_156),
.B2(n_140),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_196),
.A2(n_172),
.B1(n_175),
.B2(n_166),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_174),
.A2(n_147),
.B1(n_151),
.B2(n_146),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_138),
.Y(n_200)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_201),
.B(n_0),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_213),
.C(n_215),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_207),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_144),
.Y(n_209)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_191),
.A2(n_144),
.B1(n_119),
.B2(n_29),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_212),
.A2(n_207),
.B1(n_199),
.B2(n_201),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_178),
.A2(n_173),
.B(n_181),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_214),
.A2(n_165),
.B1(n_166),
.B2(n_162),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_163),
.B(n_136),
.C(n_125),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_173),
.A2(n_33),
.B(n_24),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_218),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_180),
.B(n_24),
.C(n_33),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_218),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_168),
.B(n_26),
.Y(n_222)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_222),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_24),
.C(n_25),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_24),
.Y(n_241)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_192),
.Y(n_224)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_224),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_198),
.B(n_167),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_240),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_232),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_219),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_200),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_233),
.B(n_3),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_234),
.A2(n_197),
.B1(n_223),
.B2(n_25),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_172),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_235),
.A2(n_204),
.B1(n_216),
.B2(n_206),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_237),
.A2(n_239),
.B1(n_244),
.B2(n_206),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_210),
.A2(n_169),
.B1(n_164),
.B2(n_170),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_242),
.Y(n_253)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_205),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_217),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_247),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_211),
.A2(n_25),
.B1(n_2),
.B2(n_3),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_203),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_245),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_195),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_246),
.B(n_220),
.Y(n_254)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_251),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_254),
.Y(n_279)
);

BUFx24_ASAP7_75t_SL g255 ( 
.A(n_226),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_226),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_215),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_256),
.B(n_259),
.C(n_272),
.Y(n_284)
);

NAND3xp33_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_213),
.C(n_208),
.Y(n_258)
);

NOR2xp67_ASAP7_75t_SL g286 ( 
.A(n_258),
.B(n_270),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_202),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_222),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_268),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_262),
.A2(n_273),
.B(n_235),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_196),
.Y(n_264)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_264),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_238),
.B(n_221),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_266),
.B(n_269),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_267),
.A2(n_234),
.B1(n_228),
.B2(n_227),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_197),
.Y(n_268)
);

AOI21xp33_ASAP7_75t_L g270 ( 
.A1(n_251),
.A2(n_16),
.B(n_3),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_230),
.B(n_0),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_274),
.B(n_277),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_232),
.Y(n_275)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_257),
.Y(n_276)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_276),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_252),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_233),
.Y(n_278)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_278),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_229),
.Y(n_281)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_281),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_268),
.B(n_231),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_291),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_253),
.B(n_229),
.Y(n_285)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_285),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_288),
.A2(n_263),
.B1(n_257),
.B2(n_267),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_259),
.B(n_241),
.C(n_248),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_284),
.C(n_283),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_290),
.A2(n_260),
.B(n_256),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_235),
.Y(n_291)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_293),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_297),
.Y(n_308)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_290),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_304),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_272),
.C(n_7),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_300),
.A2(n_306),
.B(n_279),
.Y(n_309)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_286),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_287),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_305),
.A2(n_282),
.B1(n_280),
.B2(n_11),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_5),
.C(n_8),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_312),
.C(n_319),
.Y(n_322)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_301),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_310),
.B(n_311),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_296),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_295),
.B(n_280),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_291),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_316),
.Y(n_323)
);

OR2x6_ASAP7_75t_SL g314 ( 
.A(n_294),
.B(n_276),
.Y(n_314)
);

NOR2xp67_ASAP7_75t_SL g320 ( 
.A(n_314),
.B(n_299),
.Y(n_320)
);

INVxp33_ASAP7_75t_L g316 ( 
.A(n_302),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_293),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_317),
.B(n_318),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_298),
.A2(n_9),
.B(n_10),
.Y(n_319)
);

AOI21x1_ASAP7_75t_SL g334 ( 
.A1(n_320),
.A2(n_12),
.B(n_13),
.Y(n_334)
);

MAJx2_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_295),
.C(n_300),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_308),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_307),
.A2(n_292),
.B(n_303),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_325),
.A2(n_328),
.B(n_322),
.Y(n_335)
);

INVxp33_ASAP7_75t_L g326 ( 
.A(n_315),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_327),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_306),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_329),
.A2(n_330),
.B(n_332),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_311),
.Y(n_330)
);

O2A1O1Ixp33_ASAP7_75t_SL g332 ( 
.A1(n_324),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_332)
);

AO21x1_ASAP7_75t_L g333 ( 
.A1(n_328),
.A2(n_9),
.B(n_10),
.Y(n_333)
);

AOI222xp33_ASAP7_75t_L g336 ( 
.A1(n_333),
.A2(n_334),
.B1(n_12),
.B2(n_14),
.C1(n_15),
.C2(n_331),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_335),
.A2(n_12),
.B(n_14),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_336),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_331),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_340),
.B(n_338),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_341),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_339),
.C(n_337),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_15),
.Y(n_344)
);


endmodule