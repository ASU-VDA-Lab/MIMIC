module real_jpeg_15191_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_430, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_430;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_0),
.A2(n_14),
.B(n_427),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_0),
.B(n_428),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_1),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_1),
.Y(n_87)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_1),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_2),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_2),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g173 ( 
.A(n_2),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_2),
.Y(n_222)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_3),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_3),
.Y(n_268)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_4),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_4),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_4),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_4),
.Y(n_175)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_4),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_4),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_5),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_6),
.A2(n_39),
.B1(n_40),
.B2(n_47),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_6),
.A2(n_39),
.B1(n_270),
.B2(n_273),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_6),
.A2(n_39),
.B1(n_294),
.B2(n_297),
.Y(n_293)
);

OAI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_6),
.A2(n_39),
.B1(n_369),
.B2(n_371),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_7),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_8),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_51)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_8),
.A2(n_55),
.B1(n_280),
.B2(n_284),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_8),
.A2(n_55),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g374 ( 
.A1(n_8),
.A2(n_55),
.B1(n_375),
.B2(n_378),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_10),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_10),
.Y(n_113)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_10),
.Y(n_168)
);

BUFx4f_ASAP7_75t_L g272 ( 
.A(n_10),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_11),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_11),
.B(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_11),
.A2(n_92),
.B1(n_105),
.B2(n_109),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_11),
.A2(n_92),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_11),
.B(n_70),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_11),
.B(n_220),
.C(n_223),
.Y(n_219)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_60),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_59),
.Y(n_15)
);

OR2x2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_56),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_17),
.B(n_56),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_17),
.B(n_363),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_17),
.B(n_363),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_20),
.B1(n_37),
.B2(n_51),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_18),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_19),
.B(n_20),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_29),
.Y(n_19)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_23),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_23),
.Y(n_370)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_28),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_31),
.Y(n_152)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_33),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_38),
.A2(n_100),
.B1(n_150),
.B2(n_384),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_45),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_50),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_51),
.Y(n_57)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp33_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

AND2x4_ASAP7_75t_L g149 ( 
.A(n_58),
.B(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_361),
.B(n_421),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

AO221x1_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_252),
.B1(n_353),
.B2(n_359),
.C(n_360),
.Y(n_62)
);

AO21x2_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_202),
.B(n_251),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_178),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_65),
.B(n_178),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_147),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_119),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_67),
.B(n_119),
.C(n_147),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_99),
.C(n_101),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_68),
.A2(n_154),
.B1(n_176),
.B2(n_177),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_68),
.A2(n_176),
.B1(n_180),
.B2(n_182),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g206 ( 
.A1(n_68),
.A2(n_177),
.B(n_207),
.C(n_209),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_68),
.A2(n_319),
.B(n_324),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_68),
.B(n_319),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_69),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_69),
.B(n_154),
.Y(n_209)
);

XNOR2x1_ASAP7_75t_L g258 ( 
.A(n_69),
.B(n_149),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_69),
.B(n_149),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_69),
.B(n_149),
.Y(n_308)
);

OA21x2_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_80),
.B(n_91),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_70),
.A2(n_80),
.B1(n_91),
.B2(n_368),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_71),
.A2(n_367),
.B1(n_373),
.B2(n_374),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_71),
.Y(n_386)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_75),
.B1(n_77),
.B2(n_79),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_75),
.Y(n_157)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_76),
.Y(n_160)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_80),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B1(n_86),
.B2(n_88),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_89),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_89),
.Y(n_379)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B(n_95),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_92),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_92),
.B(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_92),
.A2(n_144),
.B(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_92),
.B(n_162),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_92),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI32xp33_ASAP7_75t_L g185 ( 
.A1(n_95),
.A2(n_186),
.A3(n_188),
.B1(n_191),
.B2(n_197),
.Y(n_185)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_99),
.A2(n_102),
.B1(n_103),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_99),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_102),
.B1(n_120),
.B2(n_146),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_101),
.B(n_185),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_101),
.B(n_214),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_101),
.B(n_177),
.C(n_216),
.Y(n_246)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_102),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_102),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_102),
.B(n_231),
.Y(n_230)
);

AND2x2_ASAP7_75t_SL g241 ( 
.A(n_102),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_102),
.B(n_120),
.Y(n_334)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_114),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_104),
.A2(n_261),
.B1(n_269),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g162 ( 
.A1(n_108),
.A2(n_163),
.B1(n_165),
.B2(n_167),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_108),
.Y(n_223)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_108),
.Y(n_264)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_108),
.Y(n_274)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_112),
.Y(n_236)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_114),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_116),
.Y(n_277)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_116),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_118),
.Y(n_240)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_127),
.B(n_135),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_126),
.Y(n_187)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_126),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_133),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_138),
.B(n_143),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_153),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_148),
.A2(n_287),
.B1(n_300),
.B2(n_316),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_148),
.B(n_366),
.C(n_380),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_148),
.B(n_389),
.C(n_395),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_148),
.A2(n_391),
.B1(n_392),
.B2(n_394),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_148),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_148),
.B(n_380),
.C(n_396),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_148),
.A2(n_394),
.B1(n_406),
.B2(n_407),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_148),
.A2(n_389),
.B1(n_390),
.B2(n_394),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_149),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_149),
.B(n_154),
.Y(n_347)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_153),
.A2(n_207),
.B1(n_208),
.B2(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_153),
.Y(n_248)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_154),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_154),
.A2(n_177),
.B1(n_183),
.B2(n_184),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_154),
.A2(n_177),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_154),
.A2(n_177),
.B1(n_218),
.B2(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_154),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_154),
.B(n_304),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_154),
.A2(n_177),
.B1(n_260),
.B2(n_332),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_154),
.A2(n_177),
.B1(n_304),
.B2(n_344),
.Y(n_343)
);

AND2x4_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_161),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_155),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_290)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_157),
.Y(n_321)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AND2x2_ASAP7_75t_SL g381 ( 
.A(n_161),
.B(n_320),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_169),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_162),
.Y(n_292)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_169),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_170)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_171),
.Y(n_323)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_177),
.B(n_218),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.C(n_201),
.Y(n_178)
);

XOR2x2_ASAP7_75t_SL g204 ( 
.A(n_179),
.B(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_180),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_193),
.Y(n_198)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_200),
.Y(n_225)
);

OAI21x1_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_210),
.B(n_250),
.Y(n_202)
);

NOR2xp67_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_204),
.B(n_206),
.Y(n_250)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

AND3x1_ASAP7_75t_L g346 ( 
.A(n_209),
.B(n_308),
.C(n_347),
.Y(n_346)
);

AOI21x1_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_245),
.B(n_249),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_226),
.B(n_244),
.Y(n_211)
);

NOR2x1_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_217),
.Y(n_244)
);

INVxp67_ASAP7_75t_SL g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_218),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_224),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NOR2x1_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_241),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_237),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_247),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_337),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_325),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_254),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_309),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_255),
.B(n_309),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_286),
.C(n_301),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_256),
.B(n_286),
.Y(n_336)
);

OAI22x1_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_259),
.B2(n_285),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_257),
.B(n_334),
.Y(n_340)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_258),
.A2(n_303),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_258),
.Y(n_329)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_259),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_259),
.A2(n_302),
.B(n_306),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_260),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_269),
.B1(n_275),
.B2(n_278),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx6_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_272),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_273),
.Y(n_284)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_289),
.B1(n_290),
.B2(n_300),
.Y(n_286)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_287),
.Y(n_300)
);

NOR2xp67_ASAP7_75t_R g314 ( 
.A(n_287),
.B(n_290),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_291),
.A2(n_292),
.B1(n_293),
.B2(n_320),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_300),
.A2(n_394),
.B1(n_412),
.B2(n_430),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_301),
.B(n_336),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_303),
.B(n_306),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_302),
.A2(n_306),
.B(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_303),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_304),
.Y(n_344)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_310),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_312),
.A2(n_313),
.B1(n_317),
.B2(n_318),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_313),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_314),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_317),
.B(n_415),
.C(n_416),
.Y(n_414)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_324),
.A2(n_404),
.B1(n_405),
.B2(n_409),
.Y(n_403)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_324),
.Y(n_409)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_325),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_335),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_326),
.B(n_335),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_331),
.C(n_333),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_328),
.B(n_331),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_333),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_349),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_348),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_339),
.B(n_348),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_340),
.B(n_343),
.C(n_345),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_343),
.B1(n_345),
.B2(n_346),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_349),
.B(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

OR2x2_ASAP7_75t_L g356 ( 
.A(n_350),
.B(n_351),
.Y(n_356)
);

A2O1A1Ixp33_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_356),
.B(n_357),
.C(n_358),
.Y(n_353)
);

NAND3xp33_ASAP7_75t_SL g361 ( 
.A(n_362),
.B(n_387),
.C(n_400),
.Y(n_361)
);

A2O1A1O1Ixp25_ASAP7_75t_L g421 ( 
.A1(n_362),
.A2(n_387),
.B(n_422),
.C(n_425),
.D(n_426),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_382),
.C(n_385),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_365),
.B(n_398),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_366),
.A2(n_380),
.B1(n_381),
.B2(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_366),
.Y(n_393)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

AO21x1_ASAP7_75t_L g385 ( 
.A1(n_373),
.A2(n_374),
.B(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_380),
.A2(n_381),
.B1(n_396),
.B2(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_381),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_382),
.A2(n_383),
.B1(n_385),
.B2(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_385),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_388),
.B(n_397),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_388),
.B(n_397),
.Y(n_425)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_395),
.B(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_396),
.Y(n_408)
);

NOR2xp67_ASAP7_75t_SL g400 ( 
.A(n_401),
.B(n_417),
.Y(n_400)
);

NOR2xp67_ASAP7_75t_SL g401 ( 
.A(n_402),
.B(n_414),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_402),
.B(n_414),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_403),
.A2(n_410),
.B1(n_411),
.B2(n_413),
.Y(n_402)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_403),
.Y(n_413)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_405),
.B(n_409),
.C(n_410),
.Y(n_420)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_417),
.A2(n_423),
.B(n_424),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_420),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_418),
.B(n_420),
.Y(n_424)
);


endmodule