module fake_netlist_5_2027_n_146 (n_16, n_0, n_12, n_9, n_25, n_18, n_22, n_1, n_8, n_10, n_24, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_20, n_5, n_14, n_2, n_23, n_13, n_3, n_6, n_146);

input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_20;
input n_5;
input n_14;
input n_2;
input n_23;
input n_13;
input n_3;
input n_6;

output n_146;

wire n_137;
wire n_91;
wire n_82;
wire n_122;
wire n_142;
wire n_140;
wire n_136;
wire n_86;
wire n_124;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_144;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_111;
wire n_108;
wire n_129;
wire n_31;
wire n_66;
wire n_98;
wire n_60;
wire n_43;
wire n_107;
wire n_58;
wire n_69;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_123;
wire n_38;
wire n_113;
wire n_139;
wire n_105;
wire n_80;
wire n_125;
wire n_35;
wire n_128;
wire n_73;
wire n_92;
wire n_120;
wire n_135;
wire n_30;
wire n_33;
wire n_126;
wire n_84;
wire n_130;
wire n_29;
wire n_79;
wire n_131;
wire n_47;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_138;
wire n_71;
wire n_109;
wire n_112;
wire n_85;
wire n_95;
wire n_119;
wire n_59;
wire n_133;
wire n_55;
wire n_99;
wire n_49;
wire n_39;
wire n_54;
wire n_67;
wire n_121;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_64;
wire n_77;
wire n_106;
wire n_102;
wire n_81;
wire n_118;
wire n_28;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_134;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_141;
wire n_145;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_19),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_22),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_46),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

AND2x6_ASAP7_75t_L g51 ( 
.A(n_29),
.B(n_12),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_28),
.B(n_1),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

AND2x4_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_15),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_1),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_3),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_4),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_7),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_61),
.B(n_65),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_65),
.B(n_35),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_64),
.B(n_56),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_64),
.B(n_35),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_52),
.B(n_37),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_56),
.B(n_62),
.Y(n_71)
);

NAND2xp33_ASAP7_75t_SL g72 ( 
.A(n_58),
.B(n_37),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_56),
.B(n_41),
.Y(n_73)
);

NAND2xp33_ASAP7_75t_SL g74 ( 
.A(n_48),
.B(n_41),
.Y(n_74)
);

NAND2xp33_ASAP7_75t_SL g75 ( 
.A(n_63),
.B(n_38),
.Y(n_75)
);

NAND2xp33_ASAP7_75t_SL g76 ( 
.A(n_54),
.B(n_32),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_60),
.B(n_18),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_23),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_60),
.B(n_24),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_55),
.B(n_57),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_55),
.B(n_57),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_78),
.B(n_51),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

OAI21x1_ASAP7_75t_L g85 ( 
.A1(n_68),
.A2(n_59),
.B(n_50),
.Y(n_85)
);

AO31x2_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_50),
.A3(n_51),
.B(n_59),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

OAI21x1_ASAP7_75t_L g88 ( 
.A1(n_71),
.A2(n_51),
.B(n_53),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_53),
.B1(n_49),
.B2(n_51),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_53),
.Y(n_91)
);

OA21x2_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_49),
.B(n_51),
.Y(n_92)
);

O2A1O1Ixp5_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_53),
.B(n_75),
.C(n_81),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

AO21x2_ASAP7_75t_L g95 ( 
.A1(n_70),
.A2(n_72),
.B(n_53),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

NAND2xp33_ASAP7_75t_R g97 ( 
.A(n_92),
.B(n_96),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_87),
.Y(n_100)
);

AND2x4_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_90),
.Y(n_101)
);

NAND2xp33_ASAP7_75t_R g102 ( 
.A(n_92),
.B(n_88),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

OR2x6_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_84),
.Y(n_104)
);

AND2x4_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_91),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_82),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

CKINVDCx5p33_ASAP7_75t_R g108 ( 
.A(n_89),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_92),
.Y(n_109)
);

BUFx10_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_86),
.Y(n_111)
);

BUFx10_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_86),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_86),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_107),
.A2(n_86),
.B1(n_88),
.B2(n_111),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_101),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_101),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_104),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_112),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_108),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_109),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_103),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_110),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_110),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_120),
.A2(n_97),
.B1(n_102),
.B2(n_103),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_97),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_120),
.A2(n_102),
.B1(n_118),
.B2(n_119),
.Y(n_130)
);

INVxp33_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_126),
.B(n_121),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_114),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_130),
.A2(n_121),
.B(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

INVxp67_ASAP7_75t_SL g136 ( 
.A(n_132),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_135),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_135),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_138),
.B(n_137),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_139),
.B(n_136),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_140),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_141),
.Y(n_143)
);

AOI31xp33_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_129),
.A3(n_127),
.B(n_128),
.Y(n_144)
);

OA22x2_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_142),
.B1(n_122),
.B2(n_115),
.Y(n_145)
);

AOI221xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_142),
.B1(n_122),
.B2(n_114),
.C(n_124),
.Y(n_146)
);


endmodule