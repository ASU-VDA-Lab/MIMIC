module real_jpeg_25105_n_17 (n_108, n_8, n_116, n_0, n_111, n_2, n_10, n_114, n_9, n_12, n_6, n_11, n_14, n_110, n_112, n_7, n_117, n_3, n_5, n_4, n_109, n_115, n_1, n_118, n_16, n_15, n_13, n_113, n_17);

input n_108;
input n_8;
input n_116;
input n_0;
input n_111;
input n_2;
input n_10;
input n_114;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_110;
input n_112;
input n_7;
input n_117;
input n_3;
input n_5;
input n_4;
input n_109;
input n_115;
input n_1;
input n_118;
input n_16;
input n_15;
input n_13;
input n_113;

output n_17;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_1),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_2),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_2),
.B(n_29),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_3),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_6),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_6),
.B(n_61),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_7),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_8),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_8),
.B(n_90),
.Y(n_97)
);

FAx1_ASAP7_75t_SL g17 ( 
.A(n_9),
.B(n_18),
.CI(n_27),
.CON(n_17),
.SN(n_17)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_11),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_11),
.B(n_93),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_12),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_13),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_13),
.B(n_39),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_14),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_14),
.B(n_78),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_15),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_16),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_20),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_25),
.B(n_102),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_26),
.B(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_26),
.B(n_68),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_32),
.B(n_105),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_99),
.B(n_104),
.Y(n_32)
);

OAI321xp33_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_89),
.A3(n_92),
.B1(n_97),
.B2(n_98),
.C(n_108),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_82),
.B(n_88),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_77),
.B(n_81),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_71),
.B(n_76),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_44),
.B(n_70),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_64),
.B(n_69),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_60),
.B(n_63),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_53),
.B(n_59),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_48),
.B(n_49),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_52),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_51),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_58),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_65),
.B(n_66),
.Y(n_69)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_72),
.B(n_73),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_83),
.B(n_84),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_85),
.B(n_91),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_103),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_109),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_110),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_111),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_112),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_113),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_114),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_115),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_116),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_117),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_118),
.Y(n_96)
);


endmodule