module fake_jpeg_8098_n_135 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx11_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_0),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_28),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_18),
.A2(n_0),
.B(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_26),
.B(n_0),
.Y(n_32)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_30),
.Y(n_39)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_32),
.A2(n_23),
.B(n_12),
.Y(n_53)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_30),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_26),
.B(n_29),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_20),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_44),
.B(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_46),
.Y(n_66)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_16),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_21),
.B(n_17),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_24),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_34),
.B(n_15),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_54),
.B(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_34),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_58),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_14),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_31),
.B1(n_30),
.B2(n_14),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_59),
.A2(n_60),
.B1(n_27),
.B2(n_22),
.Y(n_65)
);

AO22x1_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_31),
.B1(n_27),
.B2(n_20),
.Y(n_60)
);

BUFx4f_ASAP7_75t_SL g63 ( 
.A(n_45),
.Y(n_63)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_65),
.A2(n_73),
.B1(n_60),
.B2(n_59),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_23),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_50),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_76),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_28),
.B1(n_19),
.B2(n_22),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_78),
.Y(n_83)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_58),
.C(n_44),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_86),
.C(n_89),
.Y(n_96)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_85),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_77),
.B(n_62),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_53),
.C(n_60),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_91),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_78),
.C(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_67),
.B(n_21),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_12),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_93),
.A2(n_42),
.B1(n_51),
.B2(n_71),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_65),
.C(n_47),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_104),
.C(n_86),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_100),
.A2(n_101),
.B1(n_103),
.B2(n_79),
.Y(n_107)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_93),
.A2(n_72),
.B(n_17),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_82),
.C(n_13),
.Y(n_112)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_63),
.C(n_42),
.Y(n_104)
);

AOI21x1_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_9),
.B(n_2),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_109),
.C(n_108),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_107),
.A2(n_108),
.B(n_113),
.Y(n_119)
);

XNOR2x1_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_83),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_63),
.Y(n_109)
);

A2O1A1O1Ixp25_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_82),
.B(n_20),
.C(n_13),
.D(n_19),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_111),
.A2(n_112),
.B(n_98),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_117),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_116),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_109),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_95),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_118),
.A2(n_87),
.B(n_90),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_99),
.B1(n_111),
.B2(n_87),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_120),
.A2(n_70),
.B1(n_64),
.B2(n_4),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_121),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_114),
.A2(n_1),
.B(n_3),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_3),
.Y(n_127)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_125),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_1),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_127),
.Y(n_130)
);

NOR3xp33_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_6),
.C(n_7),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_126),
.B(n_7),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_132),
.B(n_133),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_131),
.A2(n_122),
.B(n_6),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_130),
.Y(n_135)
);


endmodule