module real_jpeg_7522_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_470;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_0),
.A2(n_191),
.B1(n_209),
.B2(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_0),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_0),
.A2(n_105),
.B1(n_276),
.B2(n_357),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_0),
.A2(n_97),
.B1(n_276),
.B2(n_391),
.Y(n_390)
);

OAI22xp33_ASAP7_75t_L g453 ( 
.A1(n_0),
.A2(n_143),
.B1(n_276),
.B2(n_454),
.Y(n_453)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_1),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_1),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_1),
.Y(n_242)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_1),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_1),
.Y(n_416)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g327 ( 
.A(n_2),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_2),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_2),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_2),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_3),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_90)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_3),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_3),
.A2(n_94),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_3),
.A2(n_94),
.B1(n_188),
.B2(n_367),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_3),
.A2(n_94),
.B1(n_401),
.B2(n_404),
.Y(n_400)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_4),
.A2(n_186),
.B1(n_190),
.B2(n_191),
.Y(n_185)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_4),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_4),
.A2(n_160),
.B1(n_190),
.B2(n_254),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_4),
.A2(n_190),
.B1(n_352),
.B2(n_354),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_4),
.A2(n_190),
.B1(n_346),
.B2(n_347),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_5),
.A2(n_160),
.B1(n_161),
.B2(n_165),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_5),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_5),
.B(n_175),
.C(n_178),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_5),
.B(n_82),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_5),
.B(n_204),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_5),
.B(n_127),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_5),
.B(n_260),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_6),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_7),
.A2(n_37),
.B1(n_53),
.B2(n_55),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_7),
.A2(n_55),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_7),
.A2(n_55),
.B1(n_377),
.B2(n_381),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_7),
.A2(n_55),
.B1(n_80),
.B2(n_394),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_8),
.A2(n_160),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_8),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_8),
.A2(n_186),
.B1(n_206),
.B2(n_214),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_8),
.A2(n_214),
.B1(n_293),
.B2(n_295),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_8),
.A2(n_147),
.B1(n_214),
.B2(n_420),
.Y(n_419)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_11),
.Y(n_109)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_11),
.Y(n_113)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_11),
.Y(n_118)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_12),
.Y(n_85)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_13),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_13),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_13),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_14),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_14),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_14),
.A2(n_84),
.B1(n_99),
.B2(n_129),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_14),
.A2(n_99),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_14),
.A2(n_99),
.B1(n_187),
.B2(n_372),
.Y(n_371)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_16),
.A2(n_59),
.B1(n_62),
.B2(n_65),
.Y(n_58)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g332 ( 
.A1(n_16),
.A2(n_65),
.B1(n_206),
.B2(n_333),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_16),
.A2(n_65),
.B1(n_216),
.B2(n_385),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_16),
.A2(n_65),
.B1(n_433),
.B2(n_438),
.Y(n_432)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_18),
.A2(n_130),
.B1(n_168),
.B2(n_171),
.Y(n_167)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_18),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_18),
.A2(n_171),
.B1(n_206),
.B2(n_209),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_18),
.A2(n_171),
.B1(n_266),
.B2(n_269),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_18),
.A2(n_136),
.B1(n_171),
.B2(n_346),
.Y(n_345)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_531),
.B(n_534),
.Y(n_24)
);

AO21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_149),
.B(n_530),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_141),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_27),
.B(n_141),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_132),
.C(n_138),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_28),
.A2(n_29),
.B1(n_526),
.B2(n_527),
.Y(n_525)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_66),
.C(n_100),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g517 ( 
.A(n_30),
.B(n_518),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_52),
.B1(n_56),
.B2(n_58),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_31),
.A2(n_56),
.B1(n_58),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_31),
.A2(n_56),
.B1(n_133),
.B2(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_31),
.A2(n_344),
.B(n_396),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_31),
.A2(n_42),
.B1(n_396),
.B2(n_419),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_31),
.A2(n_52),
.B1(n_56),
.B2(n_503),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_32),
.A2(n_341),
.B(n_343),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_32),
.B(n_345),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g532 ( 
.A1(n_32),
.A2(n_57),
.B(n_533),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_42),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

OAI32xp33_ASAP7_75t_L g319 ( 
.A1(n_37),
.A2(n_320),
.A3(n_321),
.B1(n_322),
.B2(n_324),
.Y(n_319)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_39),
.Y(n_143)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_40),
.Y(n_321)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_41),
.Y(n_323)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_42),
.B(n_165),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_48),
.B2(n_50),
.Y(n_42)
);

INVx6_ASAP7_75t_L g353 ( 
.A(n_44),
.Y(n_353)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_46),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_46),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_46),
.Y(n_437)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g263 ( 
.A(n_47),
.Y(n_263)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_47),
.Y(n_271)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g279 ( 
.A(n_49),
.Y(n_279)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_53),
.Y(n_137)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_53),
.Y(n_421)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_54),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_56),
.A2(n_419),
.B(n_457),
.Y(n_467)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_57),
.B(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_57),
.B(n_453),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_64),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_66),
.A2(n_100),
.B1(n_101),
.B2(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_66),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_90),
.B1(n_95),
.B2(n_96),
.Y(n_66)
);

INVx3_ASAP7_75t_SL g139 ( 
.A(n_67),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_67),
.A2(n_95),
.B1(n_292),
.B2(n_351),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_67),
.A2(n_95),
.B1(n_390),
.B2(n_393),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_67),
.A2(n_90),
.B1(n_95),
.B2(n_507),
.Y(n_506)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_82),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_74),
.B1(n_75),
.B2(n_79),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_79),
.B(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_SL g257 ( 
.A1(n_80),
.A2(n_165),
.B(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_81),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_82),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_82),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

AOI22x1_ASAP7_75t_L g422 ( 
.A1(n_82),
.A2(n_139),
.B1(n_299),
.B2(n_423),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_82),
.A2(n_139),
.B1(n_431),
.B2(n_432),
.Y(n_430)
);

AO22x2_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_86),
.B2(n_88),
.Y(n_82)
);

INVx5_ASAP7_75t_L g387 ( 
.A(n_84),
.Y(n_387)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_85),
.Y(n_160)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_85),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_85),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_87),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_87),
.Y(n_357)
);

INVx6_ASAP7_75t_L g383 ( 
.A(n_87),
.Y(n_383)
);

AOI32xp33_ASAP7_75t_L g278 ( 
.A1(n_88),
.A2(n_160),
.A3(n_259),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_89),
.Y(n_281)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_95),
.B(n_265),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_95),
.A2(n_292),
.B(n_298),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_100),
.A2(n_101),
.B1(n_505),
.B2(n_506),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_100),
.B(n_502),
.C(n_505),
.Y(n_513)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_126),
.B(n_128),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_102),
.A2(n_159),
.B(n_166),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_102),
.A2(n_126),
.B1(n_213),
.B2(n_253),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_102),
.A2(n_166),
.B(n_253),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_102),
.A2(n_126),
.B1(n_356),
.B2(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_103),
.B(n_167),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_103),
.A2(n_127),
.B1(n_376),
.B2(n_384),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_103),
.A2(n_127),
.B1(n_384),
.B2(n_400),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_103),
.A2(n_127),
.B1(n_400),
.B2(n_444),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_116),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_107),
.B1(n_110),
.B2(n_114),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx5_ASAP7_75t_L g405 ( 
.A(n_115),
.Y(n_405)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_116),
.A2(n_213),
.B(n_217),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_119),
.B1(n_123),
.B2(n_125),
.Y(n_116)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_118),
.Y(n_177)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_121),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_122),
.Y(n_182)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx8_ASAP7_75t_L g307 ( 
.A(n_124),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_126),
.A2(n_217),
.B(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_127),
.B(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_128),
.Y(n_444)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_129),
.Y(n_216)
);

INVx4_ASAP7_75t_SL g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_132),
.B(n_138),
.Y(n_527)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_139),
.A2(n_257),
.B(n_264),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_139),
.B(n_299),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_139),
.A2(n_264),
.B(n_470),
.Y(n_469)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_141),
.B(n_532),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_141),
.B(n_532),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_142),
.Y(n_533)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_524),
.B(n_529),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_496),
.B(n_521),
.Y(n_150)
);

OAI311xp33_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_360),
.A3(n_472),
.B1(n_490),
.C1(n_491),
.Y(n_151)
);

AOI21x1_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_313),
.B(n_359),
.Y(n_152)
);

AO21x1_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_283),
.B(n_312),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_247),
.B(n_282),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_220),
.B(n_246),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_183),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_157),
.B(n_183),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_172),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_158),
.A2(n_172),
.B1(n_173),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_158),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx6_ASAP7_75t_L g403 ( 
.A(n_164),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_165),
.A2(n_195),
.B(n_202),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_165),
.B(n_325),
.Y(n_324)
);

OAI21xp33_ASAP7_75t_SL g341 ( 
.A1(n_165),
.A2(n_324),
.B(n_342),
.Y(n_341)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_169),
.Y(n_254)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_210),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_184),
.B(n_211),
.C(n_219),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_195),
.B(n_202),
.Y(n_184)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_185),
.Y(n_240)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx4_ASAP7_75t_SL g192 ( 
.A(n_193),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_195),
.A2(n_277),
.B1(n_330),
.B2(n_331),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_195),
.A2(n_366),
.B1(n_369),
.B2(n_371),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_195),
.A2(n_371),
.B(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_205),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_196),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_196),
.A2(n_275),
.B1(n_303),
.B2(n_308),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_196),
.A2(n_332),
.B1(n_414),
.B2(n_415),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_198),
.Y(n_407)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g368 ( 
.A(n_201),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_203),
.Y(n_233)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_204),
.Y(n_370)
);

INVx8_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx8_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_208),
.Y(n_334)
);

BUFx5_ASAP7_75t_L g374 ( 
.A(n_208),
.Y(n_374)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_209),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_218),
.B2(n_219),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NAND2xp33_ASAP7_75t_SL g280 ( 
.A(n_215),
.B(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_237),
.B(n_245),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_230),
.B(n_236),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_229),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_228),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_235),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_235),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B(n_234),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_232),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_234),
.A2(n_274),
.B(n_277),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_243),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_243),
.Y(n_245)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_241),
.Y(n_277)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_248),
.B(n_249),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_272),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_255),
.B2(n_256),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_255),
.C(n_272),
.Y(n_284)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVxp33_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_263),
.Y(n_297)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_263),
.Y(n_441)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_265),
.Y(n_299)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx12f_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_268),
.Y(n_392)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_271),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_278),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_278),
.Y(n_289)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_284),
.B(n_285),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_290),
.B2(n_311),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_288),
.B(n_289),
.C(n_311),
.Y(n_314)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_290),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_300),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_291),
.B(n_301),
.C(n_302),
.Y(n_335)
);

INVx5_ASAP7_75t_L g354 ( 
.A(n_293),
.Y(n_354)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_303),
.Y(n_330)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx5_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_314),
.B(n_315),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_338),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_335),
.B1(n_336),
.B2(n_337),
.Y(n_316)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_317),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_319),
.B1(n_328),
.B2(n_329),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_319),
.B(n_328),
.Y(n_468)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_335),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_335),
.B(n_336),
.C(n_338),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_340),
.B1(n_349),
.B2(n_358),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_339),
.B(n_350),
.C(n_355),
.Y(n_481)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_349),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_350),
.B(n_355),
.Y(n_349)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_351),
.Y(n_470)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

NAND2xp33_ASAP7_75t_SL g360 ( 
.A(n_361),
.B(n_458),
.Y(n_360)
);

A2O1A1Ixp33_ASAP7_75t_SL g491 ( 
.A1(n_361),
.A2(n_458),
.B(n_492),
.C(n_495),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_424),
.Y(n_361)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_362),
.B(n_424),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_397),
.C(n_409),
.Y(n_362)
);

FAx1_ASAP7_75t_SL g471 ( 
.A(n_363),
.B(n_397),
.CI(n_409),
.CON(n_471),
.SN(n_471)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_388),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_364),
.B(n_389),
.C(n_395),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_375),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_365),
.B(n_375),
.Y(n_464)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_366),
.Y(n_414)
);

INVx5_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

CKINVDCx14_ASAP7_75t_R g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_376),
.Y(n_412)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx3_ASAP7_75t_SL g381 ( 
.A(n_382),
.Y(n_381)
);

INVx8_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_395),
.Y(n_388)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_390),
.Y(n_423)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_393),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_398),
.A2(n_399),
.B1(n_406),
.B2(n_408),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_399),
.B(n_406),
.Y(n_448)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_406),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_406),
.A2(n_408),
.B1(n_450),
.B2(n_451),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_406),
.A2(n_448),
.B(n_451),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_417),
.C(n_422),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_410),
.B(n_462),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_413),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_411),
.B(n_413),
.Y(n_480)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_417),
.A2(n_418),
.B1(n_422),
.B2(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_422),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_426),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_425),
.B(n_428),
.C(n_446),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_428),
.B1(n_446),
.B2(n_447),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_442),
.B(n_445),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_430),
.B(n_443),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_432),
.Y(n_507)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx4_ASAP7_75t_SL g435 ( 
.A(n_436),
.Y(n_435)
);

INVx5_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

FAx1_ASAP7_75t_SL g498 ( 
.A(n_445),
.B(n_499),
.CI(n_500),
.CON(n_498),
.SN(n_498)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_445),
.B(n_499),
.C(n_500),
.Y(n_520)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_449),
.Y(n_447)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_457),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_453),
.Y(n_503)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx8_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_471),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_459),
.B(n_471),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_464),
.C(n_465),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_460),
.A2(n_461),
.B1(n_464),
.B2(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_464),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_465),
.B(n_483),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_468),
.C(n_469),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_466),
.A2(n_467),
.B1(n_469),
.B2(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_468),
.B(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_469),
.Y(n_478)
);

BUFx24_ASAP7_75t_SL g537 ( 
.A(n_471),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_473),
.B(n_485),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_474),
.A2(n_493),
.B(n_494),
.Y(n_492)
);

NOR2x1_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_482),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_475),
.B(n_482),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_479),
.C(n_481),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_476),
.B(n_488),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_479),
.A2(n_480),
.B1(n_481),
.B2(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_481),
.Y(n_489)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_487),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_486),
.B(n_487),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_510),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_498),
.B(n_509),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_498),
.B(n_509),
.Y(n_522)
);

BUFx24_ASAP7_75t_SL g536 ( 
.A(n_498),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_501),
.A2(n_502),
.B1(n_504),
.B2(n_508),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_501),
.A2(n_502),
.B1(n_516),
.B2(n_517),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_501),
.B(n_512),
.C(n_516),
.Y(n_528)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_504),
.Y(n_508)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_510),
.A2(n_522),
.B(n_523),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g510 ( 
.A(n_511),
.B(n_520),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_511),
.B(n_520),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_512),
.A2(n_513),
.B1(n_514),
.B2(n_515),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_525),
.B(n_528),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_525),
.B(n_528),
.Y(n_529)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_535),
.Y(n_534)
);


endmodule