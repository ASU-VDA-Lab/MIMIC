module fake_jpeg_23698_n_232 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_232);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_2),
.B(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g34 ( 
.A(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_28),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_45),
.B(n_47),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_32),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_50),
.B(n_27),
.Y(n_74)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_59),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_23),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_23),
.Y(n_80)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_17),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_22),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_87),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_73),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_58),
.A2(n_19),
.B1(n_22),
.B2(n_28),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_66),
.A2(n_81),
.B1(n_88),
.B2(n_91),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_57),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_70),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_56),
.A2(n_22),
.B1(n_28),
.B2(n_19),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_74),
.B(n_82),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_77),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_78),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_51),
.A2(n_19),
.B1(n_34),
.B2(n_24),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_79),
.A2(n_90),
.B1(n_93),
.B2(n_25),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_SL g106 ( 
.A(n_80),
.B(n_36),
.C(n_35),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_58),
.A2(n_20),
.B1(n_16),
.B2(n_21),
.Y(n_81)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_41),
.C(n_37),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_36),
.C(n_35),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_59),
.B(n_31),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_86),
.B(n_30),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_42),
.B(n_38),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_55),
.A2(n_20),
.B1(n_16),
.B2(n_21),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_45),
.Y(n_89)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_43),
.A2(n_34),
.B1(n_33),
.B2(n_41),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_43),
.A2(n_25),
.B1(n_21),
.B2(n_16),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_47),
.B(n_38),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_94),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_50),
.A2(n_31),
.B1(n_30),
.B2(n_33),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_47),
.B(n_38),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_101),
.A2(n_77),
.B1(n_83),
.B2(n_76),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_63),
.B(n_34),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_118),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_71),
.C(n_64),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_90),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_114),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_36),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_115),
.Y(n_129)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_85),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_62),
.B(n_27),
.Y(n_117)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_35),
.Y(n_118)
);

NOR3xp33_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_26),
.C(n_18),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_69),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_72),
.A2(n_26),
.B1(n_18),
.B2(n_15),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_78),
.B1(n_15),
.B2(n_14),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_67),
.B(n_0),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_82),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_122),
.A2(n_123),
.B(n_95),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_69),
.C(n_62),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_135),
.Y(n_150)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_127),
.B(n_130),
.Y(n_164)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_80),
.Y(n_131)
);

XNOR2x1_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_133),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_136),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_79),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_65),
.C(n_75),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_142),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_96),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_138),
.Y(n_160)
);

OAI21xp33_ASAP7_75t_SL g162 ( 
.A1(n_139),
.A2(n_68),
.B(n_61),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_73),
.Y(n_140)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

AOI221xp5_ASAP7_75t_L g146 ( 
.A1(n_141),
.A2(n_120),
.B1(n_110),
.B2(n_116),
.C(n_101),
.Y(n_146)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_105),
.Y(n_143)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_121),
.Y(n_145)
);

NOR2x1_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_108),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_146),
.A2(n_148),
.B1(n_161),
.B2(n_130),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_112),
.B1(n_95),
.B2(n_114),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_128),
.C(n_131),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_115),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_137),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_129),
.A2(n_112),
.B(n_102),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g169 ( 
.A1(n_154),
.A2(n_155),
.B(n_157),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_123),
.A2(n_113),
.B(n_100),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_126),
.B1(n_134),
.B2(n_135),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_129),
.A2(n_108),
.B(n_1),
.Y(n_157)
);

OA21x2_ASAP7_75t_SL g158 ( 
.A1(n_133),
.A2(n_0),
.B(n_1),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_157),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_142),
.A2(n_113),
.B1(n_100),
.B2(n_98),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_162),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_182)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_164),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_167),
.B(n_168),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_175),
.C(n_178),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_172),
.Y(n_195)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_128),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_180),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_174),
.A2(n_182),
.B1(n_148),
.B2(n_159),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_122),
.C(n_125),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_176),
.A2(n_158),
.B1(n_150),
.B2(n_163),
.Y(n_185)
);

OA21x2_ASAP7_75t_SL g190 ( 
.A1(n_177),
.A2(n_183),
.B(n_152),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_144),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_166),
.Y(n_179)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_179),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_124),
.C(n_13),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_13),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_147),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_160),
.B(n_2),
.Y(n_183)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_185),
.Y(n_205)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_187),
.A2(n_189),
.B1(n_169),
.B2(n_180),
.Y(n_197)
);

AOI211xp5_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_152),
.B(n_151),
.C(n_154),
.Y(n_189)
);

AOI31xp67_ASAP7_75t_L g201 ( 
.A1(n_190),
.A2(n_189),
.A3(n_185),
.B(n_178),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_173),
.B(n_155),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_194),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_175),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_160),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_197),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_195),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_199),
.B(n_203),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_153),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_200),
.Y(n_210)
);

NOR2xp67_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_192),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_184),
.Y(n_209)
);

NOR3xp33_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_153),
.C(n_147),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_166),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_207),
.C(n_192),
.Y(n_211)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_209),
.C(n_211),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_184),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_198),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_205),
.A2(n_194),
.B1(n_159),
.B2(n_12),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_213),
.A2(n_214),
.B1(n_211),
.B2(n_5),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_220),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_210),
.A2(n_206),
.B1(n_203),
.B2(n_204),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_218),
.A2(n_209),
.B1(n_212),
.B2(n_7),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_12),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_3),
.Y(n_222)
);

NOR2x1_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_213),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_222),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_223),
.B(n_217),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_226),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_224),
.B(n_4),
.C(n_5),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_227),
.A2(n_225),
.B(n_5),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_228),
.B(n_226),
.Y(n_230)
);

AO21x1_ASAP7_75t_L g231 ( 
.A1(n_230),
.A2(n_229),
.B(n_8),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_4),
.Y(n_232)
);


endmodule