module real_jpeg_12532_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_139;
wire n_33;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_0),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_1),
.A2(n_26),
.B1(n_29),
.B2(n_39),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_1),
.A2(n_39),
.B1(n_47),
.B2(n_49),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_1),
.A2(n_39),
.B1(n_62),
.B2(n_65),
.Y(n_170)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_L g34 ( 
.A1(n_4),
.A2(n_31),
.B(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_4),
.B(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_4),
.B(n_29),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_L g148 ( 
.A1(n_4),
.A2(n_37),
.B1(n_47),
.B2(n_49),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_4),
.A2(n_49),
.B(n_59),
.C(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_4),
.B(n_90),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_4),
.B(n_76),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_4),
.B(n_68),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_L g184 ( 
.A1(n_4),
.A2(n_29),
.B(n_134),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_6),
.A2(n_47),
.B1(n_49),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_6),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_6),
.A2(n_26),
.B1(n_29),
.B2(n_56),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_6),
.A2(n_56),
.B1(n_62),
.B2(n_65),
.Y(n_137)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_9),
.A2(n_26),
.B1(n_29),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_9),
.A2(n_47),
.B1(n_49),
.B2(n_53),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_9),
.A2(n_53),
.B1(n_62),
.B2(n_65),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_10),
.A2(n_47),
.B1(n_49),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_10),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_10),
.A2(n_62),
.B1(n_65),
.B2(n_67),
.Y(n_94)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_12),
.A2(n_62),
.B1(n_65),
.B2(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_12),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_13),
.A2(n_62),
.B1(n_65),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_13),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_13),
.A2(n_47),
.B1(n_49),
.B2(n_78),
.Y(n_102)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_15),
.A2(n_62),
.B1(n_65),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_15),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_16),
.A2(n_26),
.B1(n_29),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_16),
.A2(n_31),
.B1(n_32),
.B2(n_51),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_16),
.A2(n_47),
.B1(n_49),
.B2(n_51),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_16),
.A2(n_51),
.B1(n_62),
.B2(n_65),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_121),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_120),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_95),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_20),
.B(n_95),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_71),
.C(n_84),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_21),
.A2(n_22),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_23),
.B(n_41),
.C(n_70),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_34),
.B2(n_38),
.Y(n_23)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_24),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_26),
.A2(n_29),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

OAI32xp33_ASAP7_75t_L g82 ( 
.A1(n_26),
.A2(n_28),
.A3(n_31),
.B1(n_36),
.B2(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_27),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_27),
.B(n_29),
.Y(n_83)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI32xp33_ASAP7_75t_L g132 ( 
.A1(n_29),
.A2(n_44),
.A3(n_47),
.B1(n_133),
.B2(n_135),
.Y(n_132)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_32),
.B(n_37),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_37),
.A2(n_60),
.B(n_65),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_37),
.A2(n_74),
.B1(n_76),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_38),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_54),
.B1(n_69),
.B2(n_70),
.Y(n_40)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_46),
.B1(n_50),
.B2(n_52),
.Y(n_41)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_42),
.A2(n_46),
.B1(n_87),
.B2(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_45),
.B1(n_47),
.B2(n_49),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_45),
.B(n_49),
.Y(n_135)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_49),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_57),
.B1(n_66),
.B2(n_68),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_55),
.A2(n_57),
.B1(n_68),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_57),
.A2(n_68),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_57),
.A2(n_68),
.B1(n_149),
.B2(n_156),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_65),
.Y(n_61)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_61),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_61),
.A2(n_101),
.B1(n_128),
.B2(n_186),
.Y(n_185)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_62),
.B(n_172),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_66),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_71),
.B(n_84),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_81),
.B2(n_82),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_72),
.B(n_82),
.Y(n_119)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_76),
.B1(n_77),
.B2(n_79),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_76),
.B1(n_77),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_74),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_74),
.A2(n_76),
.B1(n_94),
.B2(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_74),
.A2(n_76),
.B1(n_137),
.B2(n_158),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_74),
.A2(n_76),
.B1(n_163),
.B2(n_170),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_75),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_75),
.A2(n_104),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_91),
.C(n_93),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_85),
.B(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_90),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_93),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_92),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_108),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_119),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_141),
.B(n_196),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_138),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_123),
.B(n_138),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.C(n_129),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_124),
.B(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_126),
.A2(n_129),
.B1(n_130),
.B2(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_126),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_136),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_131),
.A2(n_132),
.B1(n_136),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_136),
.Y(n_188)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_190),
.B(n_195),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_179),
.B(n_189),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_159),
.B(n_178),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_152),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_145),
.B(n_152),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_150),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_146),
.A2(n_147),
.B1(n_150),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_157),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_155),
.C(n_157),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_158),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_167),
.B(n_177),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_161),
.B(n_165),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_173),
.B(n_176),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_174),
.B(n_175),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_180),
.B(n_181),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_187),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_185),
.C(n_187),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_191),
.B(n_192),
.Y(n_195)
);


endmodule