module fake_jpeg_1907_n_136 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_136);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_46),
.Y(n_57)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

NAND2x1_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_52),
.Y(n_58)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_46),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_45),
.B1(n_35),
.B2(n_46),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_35),
.B1(n_45),
.B2(n_39),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_50),
.B(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_43),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_63),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_69),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_61),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_68),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_58),
.A2(n_49),
.B(n_43),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_72),
.C(n_70),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_61),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_71),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_41),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_41),
.C(n_44),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_73),
.A2(n_38),
.B(n_57),
.C(n_62),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_44),
.B1(n_42),
.B2(n_40),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_75),
.A2(n_58),
.B1(n_55),
.B2(n_57),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_79),
.B1(n_85),
.B2(n_1),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_60),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_80),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_61),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_84),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_53),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_70),
.A2(n_62),
.B1(n_1),
.B2(n_2),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_25),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_0),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_81),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_100),
.Y(n_104)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_93),
.Y(n_114)
);

AOI221xp5_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_112)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_87),
.B(n_62),
.Y(n_94)
);

NOR2x1_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_23),
.Y(n_111)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_32),
.C(n_30),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_101),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_77),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_85),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_102),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_2),
.B(n_3),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_103),
.B(n_105),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_92),
.A2(n_3),
.B(n_4),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_91),
.B(n_4),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_115),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_29),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_96),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_99),
.C(n_98),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_99),
.B1(n_91),
.B2(n_11),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_94),
.A2(n_28),
.B(n_21),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_119),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_105),
.B1(n_108),
.B2(n_110),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_18),
.C(n_17),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_103),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_118),
.Y(n_123)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_125),
.C(n_126),
.Y(n_128)
);

AOI321xp33_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_104),
.A3(n_111),
.B1(n_109),
.B2(n_106),
.C(n_114),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_125),
.C(n_117),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_129),
.A2(n_128),
.B1(n_130),
.B2(n_117),
.Y(n_131)
);

XOR2x2_ASAP7_75t_SL g133 ( 
.A(n_131),
.B(n_132),
.Y(n_133)
);

NOR3xp33_ASAP7_75t_SL g132 ( 
.A(n_130),
.B(n_9),
.C(n_10),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_133),
.A2(n_9),
.B(n_10),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_12),
.C(n_13),
.Y(n_136)
);


endmodule