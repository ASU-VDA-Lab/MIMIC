module fake_jpeg_12792_n_220 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_220);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_220;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_44),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_0),
.C(n_1),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_29),
.B1(n_32),
.B2(n_25),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_SL g90 ( 
.A1(n_50),
.A2(n_40),
.B(n_19),
.C(n_45),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_23),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_53),
.B(n_61),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_26),
.B1(n_32),
.B2(n_24),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_55),
.A2(n_45),
.B1(n_43),
.B2(n_39),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_47),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_67),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_44),
.B(n_18),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_58),
.B(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_18),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_31),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_62),
.B(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_31),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_30),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_65),
.B(n_66),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_30),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_19),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_28),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_71),
.A2(n_90),
.B1(n_37),
.B2(n_56),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_24),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_83),
.Y(n_100)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_38),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_77),
.Y(n_97)
);

AND2x4_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_33),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_86),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_28),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_79),
.B(n_82),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_26),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_35),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_35),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_77),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_64),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

NAND2xp33_ASAP7_75t_SL g92 ( 
.A(n_67),
.B(n_40),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_92),
.A2(n_40),
.B(n_64),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_17),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_94),
.B(n_56),
.Y(n_112)
);

AO22x1_ASAP7_75t_SL g95 ( 
.A1(n_50),
.A2(n_40),
.B1(n_37),
.B2(n_43),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_48),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_98),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_SL g98 ( 
.A(n_72),
.B(n_1),
.C(n_2),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_83),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_112),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_17),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_104),
.B(n_107),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_120),
.B1(n_84),
.B2(n_90),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_60),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_117),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_85),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_116),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_73),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_60),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_77),
.Y(n_127)
);

NOR2x1_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_91),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

INVxp33_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_133),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_127),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_132),
.B1(n_106),
.B2(n_120),
.Y(n_146)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_116),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_106),
.A2(n_71),
.B1(n_95),
.B2(n_90),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_100),
.B(n_89),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_84),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_138),
.Y(n_148)
);

OA22x2_ASAP7_75t_L g138 ( 
.A1(n_102),
.A2(n_95),
.B1(n_90),
.B2(n_74),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_100),
.B(n_84),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_139),
.B(n_142),
.Y(n_156)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_141),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_92),
.Y(n_142)
);

FAx1_ASAP7_75t_SL g144 ( 
.A(n_139),
.B(n_97),
.CI(n_107),
.CON(n_144),
.SN(n_144)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_147),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_146),
.A2(n_150),
.B1(n_68),
.B2(n_48),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_140),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_118),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_160),
.C(n_155),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_128),
.A2(n_60),
.B1(n_68),
.B2(n_109),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_109),
.B(n_110),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_151),
.A2(n_155),
.B(n_103),
.Y(n_174)
);

FAx1_ASAP7_75t_SL g152 ( 
.A(n_136),
.B(n_98),
.CI(n_110),
.CON(n_152),
.SN(n_152)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_138),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_119),
.B(n_87),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_119),
.C(n_81),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_126),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_165),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_150),
.A2(n_123),
.B1(n_143),
.B2(n_125),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_176),
.B1(n_159),
.B2(n_153),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_145),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_166),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_126),
.C(n_124),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_171),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_162),
.A2(n_142),
.B(n_138),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_168),
.A2(n_148),
.B(n_151),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_156),
.B(n_121),
.Y(n_170)
);

AOI21xp33_ASAP7_75t_L g185 ( 
.A1(n_170),
.A2(n_172),
.B(n_173),
.Y(n_185)
);

NOR2x1_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_129),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g173 ( 
.A1(n_152),
.A2(n_138),
.A3(n_141),
.B1(n_21),
.B2(n_131),
.C1(n_75),
.C2(n_25),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_174),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_103),
.Y(n_175)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_175),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_157),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_161),
.Y(n_189)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_161),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_181),
.Y(n_194)
);

OAI21x1_ASAP7_75t_SL g197 ( 
.A1(n_183),
.A2(n_188),
.B(n_168),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_175),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_189),
.B(n_169),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_148),
.B1(n_152),
.B2(n_154),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_190),
.A2(n_144),
.B1(n_176),
.B2(n_154),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_192),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_167),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_163),
.Y(n_193)
);

XOR2x2_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_179),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_170),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_199),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_186),
.A2(n_174),
.B(n_178),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_196),
.B(n_198),
.Y(n_205)
);

OAI221xp5_ASAP7_75t_SL g200 ( 
.A1(n_197),
.A2(n_188),
.B1(n_183),
.B2(n_194),
.C(n_195),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_158),
.Y(n_199)
);

NOR5xp2_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_1),
.C(n_2),
.D(n_4),
.E(n_5),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_204),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_SL g202 ( 
.A(n_192),
.B(n_185),
.C(n_181),
.Y(n_202)
);

AOI31xp33_ASAP7_75t_L g208 ( 
.A1(n_202),
.A2(n_7),
.A3(n_11),
.B(n_8),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_193),
.A2(n_187),
.B1(n_158),
.B2(n_144),
.Y(n_204)
);

OAI211xp5_ASAP7_75t_L g207 ( 
.A1(n_205),
.A2(n_9),
.B(n_15),
.C(n_13),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_207),
.B(n_209),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_208),
.B(n_205),
.Y(n_212)
);

NAND4xp25_ASAP7_75t_SL g209 ( 
.A(n_203),
.B(n_8),
.C(n_11),
.D(n_4),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_210),
.A2(n_206),
.B1(n_5),
.B2(n_6),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_212),
.A2(n_215),
.B(n_64),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_213),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_211),
.A2(n_52),
.B(n_56),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_214),
.C(n_64),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_219),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_216),
.A2(n_2),
.B(n_6),
.Y(n_219)
);


endmodule