module fake_netlist_5_220_n_72 (n_8, n_10, n_4, n_5, n_7, n_0, n_12, n_9, n_14, n_2, n_16, n_13, n_3, n_11, n_17, n_15, n_6, n_1, n_72);

input n_8;
input n_10;
input n_4;
input n_5;
input n_7;
input n_0;
input n_12;
input n_9;
input n_14;
input n_2;
input n_16;
input n_13;
input n_3;
input n_11;
input n_17;
input n_15;
input n_6;
input n_1;

output n_72;

wire n_54;
wire n_29;
wire n_43;
wire n_47;
wire n_58;
wire n_67;
wire n_69;
wire n_36;
wire n_25;
wire n_53;
wire n_18;
wire n_27;
wire n_42;
wire n_64;
wire n_22;
wire n_45;
wire n_24;
wire n_28;
wire n_46;
wire n_21;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_70;
wire n_38;
wire n_71;
wire n_61;
wire n_68;
wire n_35;
wire n_32;
wire n_41;
wire n_65;
wire n_56;
wire n_51;
wire n_63;
wire n_19;
wire n_57;
wire n_37;
wire n_59;
wire n_26;
wire n_30;
wire n_20;
wire n_33;
wire n_55;
wire n_48;
wire n_31;
wire n_23;
wire n_50;
wire n_66;
wire n_49;
wire n_52;
wire n_60;
wire n_39;

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_8),
.B(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_6),
.B(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

AND2x4_ASAP7_75t_L g29 ( 
.A(n_1),
.B(n_12),
.Y(n_29)
);

OAI22x1_ASAP7_75t_L g30 ( 
.A1(n_1),
.A2(n_9),
.B1(n_0),
.B2(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_0),
.Y(n_33)
);

INVxp67_ASAP7_75t_SL g34 ( 
.A(n_24),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_3),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_18),
.A2(n_29),
.B1(n_21),
.B2(n_19),
.Y(n_36)
);

OAI21x1_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_35),
.B(n_22),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_22),
.B(n_20),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_29),
.B(n_28),
.C(n_25),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_47),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_46),
.Y(n_59)
);

OA21x2_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_54),
.B(n_48),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_SL g61 ( 
.A1(n_55),
.A2(n_45),
.B(n_44),
.Y(n_61)
);

AOI221xp5_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_45),
.B1(n_55),
.B2(n_58),
.C(n_49),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_53),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_44),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_23),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_63),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_26),
.B1(n_23),
.B2(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_71),
.A2(n_69),
.B1(n_23),
.B2(n_60),
.Y(n_72)
);


endmodule