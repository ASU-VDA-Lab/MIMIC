module real_aes_6734_n_350 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_350);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_350;
wire n_480;
wire n_476;
wire n_758;
wire n_887;
wire n_436;
wire n_599;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_979;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_1014;
wire n_364;
wire n_421;
wire n_555;
wire n_852;
wire n_766;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_923;
wire n_894;
wire n_1034;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_742;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_353;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_537;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_478;
wire n_356;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_994;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_981;
wire n_791;
wire n_976;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_755;
wire n_532;
wire n_656;
wire n_746;
wire n_1025;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_973;
wire n_504;
wire n_725;
wire n_671;
wire n_960;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_398;
wire n_688;
wire n_609;
wire n_425;
wire n_1042;
wire n_879;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1031;
wire n_1037;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_488;
wire n_501;
wire n_1041;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_1028;
wire n_366;
wire n_727;
wire n_397;
wire n_358;
wire n_385;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_354;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_365;
wire n_899;
wire n_526;
wire n_928;
wire n_637;
wire n_653;
wire n_692;
wire n_789;
wire n_544;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_922;
wire n_633;
wire n_482;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_575;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_888;
wire n_836;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1024;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g780 ( .A1(n_0), .A2(n_151), .B1(n_781), .B2(n_782), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_1), .B(n_417), .Y(n_500) );
XOR2x2_ASAP7_75t_L g457 ( .A(n_2), .B(n_458), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_3), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g945 ( .A1(n_4), .A2(n_260), .B1(n_394), .B2(n_652), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_5), .A2(n_320), .B1(n_709), .B2(n_719), .Y(n_798) );
CKINVDCx20_ASAP7_75t_R g679 ( .A(n_6), .Y(n_679) );
AO22x2_ASAP7_75t_L g372 ( .A1(n_7), .A2(n_193), .B1(n_373), .B2(n_374), .Y(n_372) );
INVx1_ASAP7_75t_L g998 ( .A(n_7), .Y(n_998) );
AOI22xp33_ASAP7_75t_SL g860 ( .A1(n_8), .A2(n_179), .B1(n_464), .B2(n_861), .Y(n_860) );
AOI22xp5_ASAP7_75t_SL g1020 ( .A1(n_9), .A2(n_347), .B1(n_568), .B2(n_782), .Y(n_1020) );
AOI222xp33_ASAP7_75t_L g590 ( .A1(n_10), .A2(n_50), .B1(n_293), .B2(n_591), .C1(n_592), .C2(n_593), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g495 ( .A1(n_11), .A2(n_270), .B1(n_404), .B2(n_496), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_12), .A2(n_55), .B1(n_628), .B2(n_923), .Y(n_922) );
AOI22xp5_ASAP7_75t_SL g1016 ( .A1(n_13), .A2(n_220), .B1(n_655), .B2(n_976), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_14), .A2(n_93), .B1(n_446), .B2(n_572), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_15), .A2(n_20), .B1(n_652), .B2(n_805), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_16), .A2(n_349), .B1(n_472), .B2(n_723), .Y(n_867) );
CKINVDCx20_ASAP7_75t_R g953 ( .A(n_17), .Y(n_953) );
CKINVDCx20_ASAP7_75t_R g847 ( .A(n_18), .Y(n_847) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_19), .A2(n_339), .B1(n_468), .B2(n_469), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_21), .A2(n_236), .B1(n_442), .B2(n_507), .Y(n_952) );
INVx1_ASAP7_75t_L g482 ( .A(n_22), .Y(n_482) );
AOI221xp5_ASAP7_75t_L g583 ( .A1(n_23), .A2(n_221), .B1(n_476), .B2(n_584), .C(n_585), .Y(n_583) );
AOI22xp33_ASAP7_75t_SL g1013 ( .A1(n_24), .A2(n_154), .B1(n_478), .B2(n_1014), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_25), .A2(n_309), .B1(n_514), .B2(n_515), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_26), .A2(n_86), .B1(n_395), .B2(n_484), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_27), .A2(n_564), .B1(n_594), .B2(n_595), .Y(n_563) );
INVx1_ASAP7_75t_L g594 ( .A(n_27), .Y(n_594) );
AOI22xp33_ASAP7_75t_SL g934 ( .A1(n_28), .A2(n_46), .B1(n_607), .B2(n_657), .Y(n_934) );
AO22x2_ASAP7_75t_L g376 ( .A1(n_29), .A2(n_98), .B1(n_373), .B2(n_377), .Y(n_376) );
AOI22xp33_ASAP7_75t_SL g834 ( .A1(n_30), .A2(n_231), .B1(n_548), .B2(n_835), .Y(n_834) );
AOI22xp33_ASAP7_75t_SL g967 ( .A1(n_31), .A2(n_90), .B1(n_592), .B2(n_628), .Y(n_967) );
CKINVDCx20_ASAP7_75t_R g588 ( .A(n_32), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_33), .A2(n_248), .B1(n_424), .B2(n_572), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_34), .A2(n_226), .B1(n_409), .B2(n_416), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_35), .Y(n_705) );
AOI22xp33_ASAP7_75t_SL g399 ( .A1(n_36), .A2(n_304), .B1(n_400), .B2(n_404), .Y(n_399) );
AOI22xp33_ASAP7_75t_SL g783 ( .A1(n_37), .A2(n_297), .B1(n_553), .B2(n_714), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_38), .A2(n_198), .B1(n_642), .B2(n_643), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g391 ( .A(n_39), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_40), .B(n_416), .Y(n_926) );
AOI22xp33_ASAP7_75t_SL g940 ( .A1(n_41), .A2(n_243), .B1(n_422), .B2(n_713), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_42), .A2(n_240), .B1(n_393), .B2(n_533), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g620 ( .A(n_43), .Y(n_620) );
AOI22xp33_ASAP7_75t_SL g768 ( .A1(n_44), .A2(n_171), .B1(n_393), .B2(n_769), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_45), .A2(n_124), .B1(n_465), .B2(n_655), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_47), .B(n_481), .Y(n_677) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_48), .Y(n_819) );
AOI22xp33_ASAP7_75t_SL g740 ( .A1(n_49), .A2(n_302), .B1(n_717), .B2(n_741), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_51), .A2(n_188), .B1(n_472), .B2(n_612), .Y(n_611) );
CKINVDCx20_ASAP7_75t_R g577 ( .A(n_52), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_53), .A2(n_165), .B1(n_423), .B2(n_609), .Y(n_608) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_54), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_56), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_57), .A2(n_336), .B1(n_507), .B2(n_508), .Y(n_506) );
AOI22xp33_ASAP7_75t_SL g504 ( .A1(n_58), .A2(n_267), .B1(n_442), .B2(n_505), .Y(n_504) );
AOI22xp5_ASAP7_75t_SL g726 ( .A1(n_59), .A2(n_727), .B1(n_747), .B2(n_748), .Y(n_726) );
CKINVDCx16_ASAP7_75t_R g748 ( .A(n_59), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_60), .A2(n_180), .B1(n_606), .B2(n_722), .Y(n_839) );
AOI222xp33_ASAP7_75t_L g659 ( .A1(n_61), .A2(n_178), .B1(n_211), .B2(n_660), .C1(n_661), .C2(n_662), .Y(n_659) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_62), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_63), .Y(n_737) );
AOI22xp33_ASAP7_75t_SL g428 ( .A1(n_64), .A2(n_67), .B1(n_429), .B2(n_433), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_65), .A2(n_251), .B1(n_606), .B2(n_607), .Y(n_605) );
AOI22xp33_ASAP7_75t_SL g787 ( .A1(n_66), .A2(n_241), .B1(n_469), .B2(n_788), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_68), .A2(n_227), .B1(n_386), .B2(n_401), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_69), .A2(n_206), .B1(n_446), .B2(n_642), .Y(n_903) );
AOI22xp33_ASAP7_75t_SL g420 ( .A1(n_70), .A2(n_212), .B1(n_421), .B2(n_423), .Y(n_420) );
AOI22xp5_ASAP7_75t_SL g1017 ( .A1(n_71), .A2(n_224), .B1(n_465), .B2(n_1018), .Y(n_1017) );
AOI22xp33_ASAP7_75t_SL g927 ( .A1(n_72), .A2(n_199), .B1(n_484), .B2(n_928), .Y(n_927) );
OA22x2_ASAP7_75t_L g363 ( .A1(n_73), .A2(n_364), .B1(n_365), .B2(n_452), .Y(n_363) );
CKINVDCx20_ASAP7_75t_R g364 ( .A(n_73), .Y(n_364) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_74), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_75), .A2(n_222), .B1(n_469), .B2(n_561), .Y(n_560) );
AOI22xp33_ASAP7_75t_SL g746 ( .A1(n_76), .A2(n_113), .B1(n_465), .B2(n_657), .Y(n_746) );
AOI22xp33_ASAP7_75t_SL g557 ( .A1(n_77), .A2(n_250), .B1(n_505), .B2(n_558), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_78), .A2(n_274), .B1(n_472), .B2(n_645), .Y(n_858) );
AOI22xp33_ASAP7_75t_SL g552 ( .A1(n_79), .A2(n_190), .B1(n_553), .B2(n_555), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_80), .A2(n_103), .B1(n_607), .B2(n_655), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g944 ( .A(n_81), .Y(n_944) );
AO22x2_ASAP7_75t_L g382 ( .A1(n_82), .A2(n_230), .B1(n_373), .B2(n_374), .Y(n_382) );
INVx1_ASAP7_75t_L g995 ( .A(n_82), .Y(n_995) );
CKINVDCx20_ASAP7_75t_R g1035 ( .A(n_83), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_84), .A2(n_87), .B1(n_548), .B2(n_550), .Y(n_547) );
AOI22xp33_ASAP7_75t_SL g974 ( .A1(n_85), .A2(n_288), .B1(n_449), .B2(n_558), .Y(n_974) );
AOI22xp5_ASAP7_75t_SL g1021 ( .A1(n_88), .A2(n_184), .B1(n_606), .B2(n_788), .Y(n_1021) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_89), .A2(n_268), .B1(n_657), .B2(n_658), .Y(n_656) );
AOI211xp5_ASAP7_75t_L g975 ( .A1(n_91), .A2(n_976), .B(n_977), .C(n_980), .Y(n_975) );
AOI22xp33_ASAP7_75t_SL g969 ( .A1(n_92), .A2(n_256), .B1(n_400), .B2(n_404), .Y(n_969) );
CKINVDCx20_ASAP7_75t_R g908 ( .A(n_94), .Y(n_908) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_95), .A2(n_602), .B1(n_633), .B2(n_634), .Y(n_601) );
INVx1_ASAP7_75t_L g633 ( .A(n_95), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_96), .A2(n_102), .B1(n_661), .B2(n_662), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_97), .A2(n_157), .B1(n_401), .B2(n_876), .Y(n_875) );
INVx1_ASAP7_75t_L g999 ( .A(n_98), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_99), .B(n_627), .Y(n_626) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_100), .Y(n_695) );
CKINVDCx20_ASAP7_75t_R g586 ( .A(n_101), .Y(n_586) );
AOI22xp33_ASAP7_75t_SL g651 ( .A1(n_104), .A2(n_305), .B1(n_401), .B2(n_652), .Y(n_651) );
AOI22xp33_ASAP7_75t_SL g785 ( .A1(n_105), .A2(n_175), .B1(n_741), .B2(n_786), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_106), .B(n_409), .Y(n_947) );
AOI22xp33_ASAP7_75t_SL g774 ( .A1(n_107), .A2(n_182), .B1(n_775), .B2(n_777), .Y(n_774) );
AOI22xp33_ASAP7_75t_SL g438 ( .A1(n_108), .A2(n_242), .B1(n_439), .B2(n_442), .Y(n_438) );
AOI22xp33_ASAP7_75t_SL g1040 ( .A1(n_109), .A2(n_155), .B1(n_533), .B2(n_928), .Y(n_1040) );
AOI22xp33_ASAP7_75t_SL g1043 ( .A1(n_110), .A2(n_275), .B1(n_465), .B2(n_655), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_111), .A2(n_121), .B1(n_496), .B2(n_533), .Y(n_676) );
AOI22xp33_ASAP7_75t_SL g931 ( .A1(n_112), .A2(n_162), .B1(n_424), .B2(n_835), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_114), .A2(n_306), .B1(n_657), .B2(n_796), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_115), .A2(n_214), .B1(n_401), .B2(n_484), .Y(n_501) );
AOI22xp33_ASAP7_75t_SL g1008 ( .A1(n_116), .A2(n_314), .B1(n_496), .B2(n_769), .Y(n_1008) );
AOI22xp33_ASAP7_75t_SL g445 ( .A1(n_117), .A2(n_132), .B1(n_446), .B2(n_449), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_118), .A2(n_167), .B1(n_409), .B2(n_802), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_119), .A2(n_334), .B1(n_719), .B2(n_722), .Y(n_718) );
XNOR2x2_ASAP7_75t_L g791 ( .A(n_120), .B(n_792), .Y(n_791) );
AOI221xp5_ASAP7_75t_L g565 ( .A1(n_122), .A2(n_186), .B1(n_548), .B2(n_566), .C(n_569), .Y(n_565) );
INVx1_ASAP7_75t_L g517 ( .A(n_123), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g948 ( .A(n_125), .B(n_417), .Y(n_948) );
AND2x6_ASAP7_75t_L g355 ( .A(n_126), .B(n_356), .Y(n_355) );
HB1xp67_ASAP7_75t_L g992 ( .A(n_126), .Y(n_992) );
AOI22xp33_ASAP7_75t_SL g685 ( .A1(n_127), .A2(n_338), .B1(n_472), .B2(n_568), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_128), .A2(n_164), .B1(n_511), .B2(n_741), .Y(n_840) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_129), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g773 ( .A(n_130), .B(n_650), .Y(n_773) );
AOI22xp33_ASAP7_75t_SL g686 ( .A1(n_131), .A2(n_322), .B1(n_421), .B2(n_469), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_133), .A2(n_168), .B1(n_424), .B2(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g772 ( .A(n_134), .B(n_416), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g647 ( .A(n_135), .Y(n_647) );
AOI22xp33_ASAP7_75t_SL g878 ( .A1(n_136), .A2(n_158), .B1(n_511), .B2(n_879), .Y(n_878) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_137), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_138), .B(n_499), .Y(n_925) );
CKINVDCx20_ASAP7_75t_R g854 ( .A(n_139), .Y(n_854) );
AOI222xp33_ASAP7_75t_L g806 ( .A1(n_140), .A2(n_181), .B1(n_310), .B2(n_481), .C1(n_593), .C2(n_807), .Y(n_806) );
NAND2xp5_ASAP7_75t_SL g1039 ( .A(n_141), .B(n_650), .Y(n_1039) );
AOI22xp33_ASAP7_75t_SL g970 ( .A1(n_142), .A2(n_207), .B1(n_409), .B2(n_416), .Y(n_970) );
AO22x2_ASAP7_75t_L g380 ( .A1(n_143), .A2(n_223), .B1(n_373), .B2(n_377), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g996 ( .A(n_143), .B(n_997), .Y(n_996) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_144), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g981 ( .A(n_145), .Y(n_981) );
AOI22xp33_ASAP7_75t_SL g951 ( .A1(n_146), .A2(n_263), .B1(n_441), .B2(n_721), .Y(n_951) );
AOI221xp5_ASAP7_75t_L g575 ( .A1(n_147), .A2(n_174), .B1(n_461), .B2(n_550), .C(n_576), .Y(n_575) );
AOI22xp33_ASAP7_75t_SL g1046 ( .A1(n_148), .A2(n_238), .B1(n_468), .B2(n_717), .Y(n_1046) );
AOI22xp33_ASAP7_75t_SL g708 ( .A1(n_149), .A2(n_160), .B1(n_561), .B2(n_709), .Y(n_708) );
AOI22xp33_ASAP7_75t_SL g972 ( .A1(n_150), .A2(n_239), .B1(n_421), .B2(n_973), .Y(n_972) );
CKINVDCx20_ASAP7_75t_R g906 ( .A(n_152), .Y(n_906) );
AOI22xp33_ASAP7_75t_SL g1036 ( .A1(n_153), .A2(n_244), .B1(n_628), .B2(n_923), .Y(n_1036) );
CKINVDCx20_ASAP7_75t_R g624 ( .A(n_156), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_159), .A2(n_232), .B1(n_507), .B2(n_657), .Y(n_880) );
AOI22xp33_ASAP7_75t_SL g710 ( .A1(n_161), .A2(n_296), .B1(n_711), .B2(n_714), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g631 ( .A(n_163), .Y(n_631) );
AOI22xp33_ASAP7_75t_SL g1045 ( .A1(n_166), .A2(n_176), .B1(n_424), .B2(n_469), .Y(n_1045) );
CKINVDCx20_ASAP7_75t_R g849 ( .A(n_169), .Y(n_849) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_170), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g966 ( .A(n_172), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_173), .A2(n_271), .B1(n_450), .B2(n_658), .Y(n_862) );
AOI22xp33_ASAP7_75t_SL g1042 ( .A1(n_177), .A2(n_328), .B1(n_461), .B2(n_553), .Y(n_1042) );
XNOR2xp5_ASAP7_75t_L g962 ( .A(n_183), .B(n_963), .Y(n_962) );
AOI22xp33_ASAP7_75t_SL g682 ( .A1(n_185), .A2(n_213), .B1(n_446), .B2(n_655), .Y(n_682) );
AOI22xp33_ASAP7_75t_SL g683 ( .A1(n_187), .A2(n_205), .B1(n_465), .B2(n_512), .Y(n_683) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_189), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_191), .A2(n_210), .B1(n_450), .B2(n_472), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_192), .A2(n_311), .B1(n_615), .B2(n_616), .Y(n_614) );
NAND2xp5_ASAP7_75t_SL g1012 ( .A(n_194), .B(n_650), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_195), .A2(n_327), .B1(n_385), .B2(n_496), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g580 ( .A(n_196), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_197), .A2(n_235), .B1(n_514), .B2(n_515), .Y(n_941) );
AOI22xp33_ASAP7_75t_SL g836 ( .A1(n_200), .A2(n_277), .B1(n_796), .B2(n_837), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g979 ( .A(n_201), .B(n_714), .Y(n_979) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_202), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_203), .A2(n_333), .B1(n_461), .B2(n_743), .Y(n_742) );
OA22x2_ASAP7_75t_L g667 ( .A1(n_204), .A2(n_668), .B1(n_669), .B2(n_670), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_204), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_208), .A2(n_225), .B1(n_505), .B2(n_645), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_209), .A2(n_299), .B1(n_550), .B2(n_643), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_215), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_216), .B(n_416), .Y(n_1038) );
CKINVDCx20_ASAP7_75t_R g1007 ( .A(n_217), .Y(n_1007) );
AOI22xp33_ASAP7_75t_SL g866 ( .A1(n_218), .A2(n_266), .B1(n_505), .B2(n_515), .Y(n_866) );
INVx2_ASAP7_75t_L g359 ( .A(n_219), .Y(n_359) );
CKINVDCx20_ASAP7_75t_R g674 ( .A(n_228), .Y(n_674) );
XNOR2x1_ASAP7_75t_L g917 ( .A(n_229), .B(n_918), .Y(n_917) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_233), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g846 ( .A(n_234), .Y(n_846) );
CKINVDCx20_ASAP7_75t_R g831 ( .A(n_237), .Y(n_831) );
AOI22xp33_ASAP7_75t_SL g716 ( .A1(n_245), .A2(n_265), .B1(n_508), .B2(n_717), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g915 ( .A(n_246), .Y(n_915) );
CKINVDCx20_ASAP7_75t_R g893 ( .A(n_247), .Y(n_893) );
CKINVDCx20_ASAP7_75t_R g870 ( .A(n_249), .Y(n_870) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_252), .Y(n_829) );
OA22x2_ASAP7_75t_L g885 ( .A1(n_253), .A2(n_886), .B1(n_887), .B2(n_888), .Y(n_885) );
CKINVDCx16_ASAP7_75t_R g886 ( .A(n_253), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_254), .B(n_650), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_255), .A2(n_324), .B1(n_464), .B2(n_465), .Y(n_463) );
INVx1_ASAP7_75t_L g373 ( .A(n_257), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_257), .Y(n_375) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_258), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g852 ( .A(n_259), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_261), .A2(n_308), .B1(n_658), .B2(n_837), .Y(n_904) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_262), .Y(n_383) );
AOI22xp33_ASAP7_75t_SL g510 ( .A1(n_264), .A2(n_300), .B1(n_511), .B2(n_512), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g913 ( .A(n_269), .Y(n_913) );
AOI211xp5_ASAP7_75t_L g350 ( .A1(n_272), .A2(n_351), .B(n_360), .C(n_1000), .Y(n_350) );
CKINVDCx20_ASAP7_75t_R g573 ( .A(n_273), .Y(n_573) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_276), .Y(n_619) );
CKINVDCx20_ASAP7_75t_R g896 ( .A(n_278), .Y(n_896) );
CKINVDCx20_ASAP7_75t_R g899 ( .A(n_279), .Y(n_899) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_280), .A2(n_762), .B1(n_763), .B2(n_789), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_280), .Y(n_762) );
XNOR2x1_ASAP7_75t_L g842 ( .A(n_281), .B(n_843), .Y(n_842) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_282), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g900 ( .A(n_283), .Y(n_900) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_284), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_285), .A2(n_331), .B1(n_405), .B2(n_478), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g630 ( .A(n_286), .Y(n_630) );
CKINVDCx20_ASAP7_75t_R g881 ( .A(n_287), .Y(n_881) );
INVx1_ASAP7_75t_L g358 ( .A(n_289), .Y(n_358) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_290), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g1028 ( .A(n_291), .Y(n_1028) );
INVx1_ASAP7_75t_L g356 ( .A(n_292), .Y(n_356) );
CKINVDCx20_ASAP7_75t_R g894 ( .A(n_294), .Y(n_894) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_295), .Y(n_522) );
AOI22xp33_ASAP7_75t_SL g745 ( .A1(n_298), .A2(n_337), .B1(n_468), .B2(n_514), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_301), .A2(n_345), .B1(n_395), .B2(n_404), .Y(n_850) );
XOR2x2_ASAP7_75t_L g812 ( .A(n_303), .B(n_813), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_307), .B(n_475), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_312), .A2(n_343), .B1(n_394), .B2(n_652), .Y(n_871) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_313), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g921 ( .A(n_315), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_316), .B(n_499), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_317), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_318), .A2(n_348), .B1(n_475), .B2(n_476), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_319), .Y(n_570) );
AOI22xp5_ASAP7_75t_SL g1001 ( .A1(n_321), .A2(n_1002), .B1(n_1003), .B2(n_1022), .Y(n_1001) );
CKINVDCx20_ASAP7_75t_R g1022 ( .A(n_321), .Y(n_1022) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_323), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_325), .A2(n_335), .B1(n_572), .B2(n_788), .Y(n_799) );
XNOR2x1_ASAP7_75t_L g518 ( .A(n_326), .B(n_519), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g978 ( .A(n_329), .Y(n_978) );
CKINVDCx20_ASAP7_75t_R g680 ( .A(n_330), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_332), .B(n_417), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_340), .B(n_533), .Y(n_827) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_341), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g694 ( .A(n_342), .Y(n_694) );
CKINVDCx20_ASAP7_75t_R g664 ( .A(n_344), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_346), .B(n_1011), .Y(n_1010) );
CKINVDCx20_ASAP7_75t_R g351 ( .A(n_352), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_353), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_355), .B(n_357), .Y(n_354) );
HB1xp67_ASAP7_75t_L g991 ( .A(n_356), .Y(n_991) );
OAI21xp5_ASAP7_75t_L g1026 ( .A1(n_357), .A2(n_990), .B(n_1027), .Y(n_1026) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_755), .B1(n_985), .B2(n_986), .C(n_987), .Y(n_360) );
INVx1_ASAP7_75t_L g985 ( .A(n_361), .Y(n_985) );
XOR2xp5_ASAP7_75t_L g361 ( .A(n_362), .B(n_598), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_453), .B1(n_454), .B2(n_597), .Y(n_362) );
INVx1_ASAP7_75t_L g597 ( .A(n_363), .Y(n_597) );
INVx1_ASAP7_75t_L g452 ( .A(n_365), .Y(n_452) );
NAND3xp33_ASAP7_75t_L g365 ( .A(n_366), .B(n_419), .C(n_437), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_367), .B(n_398), .Y(n_366) );
OAI222xp33_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_383), .B1(n_384), .B2(n_391), .C1(n_392), .C2(n_397), .Y(n_367) );
OAI221xp5_ASAP7_75t_L g623 ( .A1(n_368), .A2(n_384), .B1(n_624), .B2(n_625), .C(n_626), .Y(n_623) );
BUFx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx4_ASAP7_75t_L g591 ( .A(n_369), .Y(n_591) );
OAI21xp5_ASAP7_75t_L g869 ( .A1(n_369), .A2(n_870), .B(n_871), .Y(n_869) );
OAI21xp5_ASAP7_75t_SL g920 ( .A1(n_369), .A2(n_921), .B(n_922), .Y(n_920) );
OAI21xp5_ASAP7_75t_L g943 ( .A1(n_369), .A2(n_944), .B(n_945), .Y(n_943) );
OAI21xp5_ASAP7_75t_SL g1006 ( .A1(n_369), .A2(n_1007), .B(n_1008), .Y(n_1006) );
INVx4_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx3_ASAP7_75t_L g481 ( .A(n_370), .Y(n_481) );
INVx2_ASAP7_75t_L g494 ( .A(n_370), .Y(n_494) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_370), .Y(n_660) );
INVx2_ASAP7_75t_SL g699 ( .A(n_370), .Y(n_699) );
AND2x6_ASAP7_75t_L g370 ( .A(n_371), .B(n_378), .Y(n_370) );
AND2x4_ASAP7_75t_L g405 ( .A(n_371), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g543 ( .A(n_371), .Y(n_543) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_376), .Y(n_371) );
AND2x2_ASAP7_75t_L g390 ( .A(n_372), .B(n_380), .Y(n_390) );
INVx2_ASAP7_75t_L g415 ( .A(n_372), .Y(n_415) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g377 ( .A(n_375), .Y(n_377) );
INVx2_ASAP7_75t_L g389 ( .A(n_376), .Y(n_389) );
INVx1_ASAP7_75t_L g403 ( .A(n_376), .Y(n_403) );
OR2x2_ASAP7_75t_L g414 ( .A(n_376), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g418 ( .A(n_376), .B(n_415), .Y(n_418) );
AND2x4_ASAP7_75t_L g422 ( .A(n_378), .B(n_418), .Y(n_422) );
AND2x6_ASAP7_75t_L g441 ( .A(n_378), .B(n_413), .Y(n_441) );
AND2x2_ASAP7_75t_L g448 ( .A(n_378), .B(n_427), .Y(n_448) );
AND2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_381), .Y(n_378) );
AND2x2_ASAP7_75t_L g412 ( .A(n_379), .B(n_382), .Y(n_412) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g426 ( .A(n_380), .B(n_407), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_380), .B(n_382), .Y(n_436) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g388 ( .A(n_382), .Y(n_388) );
INVx1_ASAP7_75t_L g407 ( .A(n_382), .Y(n_407) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_385), .Y(n_384) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_386), .Y(n_484) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_386), .Y(n_533) );
BUFx2_ASAP7_75t_L g807 ( .A(n_386), .Y(n_807) );
BUFx4f_ASAP7_75t_SL g876 ( .A(n_386), .Y(n_876) );
AND2x4_ASAP7_75t_L g386 ( .A(n_387), .B(n_390), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx1_ASAP7_75t_L g396 ( .A(n_388), .Y(n_396) );
AND2x2_ASAP7_75t_L g427 ( .A(n_389), .B(n_415), .Y(n_427) );
INVx1_ASAP7_75t_L g516 ( .A(n_389), .Y(n_516) );
AND2x4_ASAP7_75t_L g395 ( .A(n_390), .B(n_396), .Y(n_395) );
AND2x4_ASAP7_75t_L g401 ( .A(n_390), .B(n_402), .Y(n_401) );
NAND2x1p5_ASAP7_75t_L g538 ( .A(n_390), .B(n_516), .Y(n_538) );
OAI222xp33_ASAP7_75t_L g696 ( .A1(n_392), .A2(n_697), .B1(n_698), .B2(n_699), .C1(n_700), .C2(n_701), .Y(n_696) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx4f_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx12f_ASAP7_75t_L g496 ( .A(n_395), .Y(n_496) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_395), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_408), .Y(n_398) );
BUFx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx3_ASAP7_75t_L g478 ( .A(n_401), .Y(n_478) );
INVx1_ASAP7_75t_L g776 ( .A(n_401), .Y(n_776) );
BUFx2_ASAP7_75t_L g928 ( .A(n_401), .Y(n_928) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OR2x6_ASAP7_75t_L g435 ( .A(n_403), .B(n_436), .Y(n_435) );
BUFx3_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx6f_ASAP7_75t_L g652 ( .A(n_405), .Y(n_652) );
BUFx2_ASAP7_75t_SL g923 ( .A(n_405), .Y(n_923) );
BUFx2_ASAP7_75t_SL g1014 ( .A(n_405), .Y(n_1014) );
INVx1_ASAP7_75t_L g544 ( .A(n_406), .Y(n_544) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
BUFx6f_ASAP7_75t_L g650 ( .A(n_409), .Y(n_650) );
INVx5_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g475 ( .A(n_410), .Y(n_475) );
INVx2_ASAP7_75t_L g499 ( .A(n_410), .Y(n_499) );
INVx4_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x4_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
AND2x6_ASAP7_75t_L g417 ( .A(n_412), .B(n_418), .Y(n_417) );
AND2x4_ASAP7_75t_L g451 ( .A(n_412), .B(n_427), .Y(n_451) );
INVx1_ASAP7_75t_L g525 ( .A(n_412), .Y(n_525) );
NAND2x1p5_ASAP7_75t_L g529 ( .A(n_412), .B(n_418), .Y(n_529) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g524 ( .A(n_414), .B(n_525), .Y(n_524) );
BUFx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx4f_ASAP7_75t_L g476 ( .A(n_417), .Y(n_476) );
INVx1_ASAP7_75t_SL g803 ( .A(n_417), .Y(n_803) );
AND2x2_ASAP7_75t_L g432 ( .A(n_418), .B(n_426), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_418), .B(n_426), .Y(n_579) );
AND2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_428), .Y(n_419) );
BUFx3_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx6_ASAP7_75t_L g462 ( .A(n_422), .Y(n_462) );
BUFx3_ASAP7_75t_L g511 ( .A(n_422), .Y(n_511) );
BUFx3_ASAP7_75t_L g561 ( .A(n_422), .Y(n_561) );
BUFx3_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
BUFx3_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx3_ASAP7_75t_L g505 ( .A(n_425), .Y(n_505) );
BUFx3_ASAP7_75t_L g568 ( .A(n_425), .Y(n_568) );
BUFx3_ASAP7_75t_L g721 ( .A(n_425), .Y(n_721) );
AND2x2_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_426), .B(n_427), .Y(n_911) );
AND2x4_ASAP7_75t_L g443 ( .A(n_427), .B(n_444), .Y(n_443) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g464 ( .A(n_431), .Y(n_464) );
INVx5_ASAP7_75t_L g512 ( .A(n_431), .Y(n_512) );
BUFx3_ASAP7_75t_L g554 ( .A(n_431), .Y(n_554) );
INVx3_ASAP7_75t_L g657 ( .A(n_431), .Y(n_657) );
INVx4_ASAP7_75t_L g713 ( .A(n_431), .Y(n_713) );
INVx8_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx2_ASAP7_75t_L g465 ( .A(n_434), .Y(n_465) );
BUFx2_ASAP7_75t_L g582 ( .A(n_434), .Y(n_582) );
BUFx4f_ASAP7_75t_SL g616 ( .A(n_434), .Y(n_616) );
BUFx2_ASAP7_75t_L g658 ( .A(n_434), .Y(n_658) );
INVx6_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_SL g555 ( .A(n_435), .Y(n_555) );
INVx1_ASAP7_75t_SL g714 ( .A(n_435), .Y(n_714) );
INVx1_ASAP7_75t_L g796 ( .A(n_435), .Y(n_796) );
INVx1_ASAP7_75t_L g444 ( .A(n_436), .Y(n_444) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_445), .Y(n_437) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx5_ASAP7_75t_SL g508 ( .A(n_440), .Y(n_508) );
INVx4_ASAP7_75t_L g572 ( .A(n_440), .Y(n_572) );
INVx2_ASAP7_75t_L g642 ( .A(n_440), .Y(n_642) );
INVx2_ASAP7_75t_SL g879 ( .A(n_440), .Y(n_879) );
INVx11_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx11_ASAP7_75t_L g470 ( .A(n_441), .Y(n_470) );
BUFx3_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx3_ASAP7_75t_L g472 ( .A(n_443), .Y(n_472) );
INVx1_ASAP7_75t_L g559 ( .A(n_443), .Y(n_559) );
BUFx3_ASAP7_75t_L g643 ( .A(n_443), .Y(n_643) );
BUFx2_ASAP7_75t_SL g717 ( .A(n_443), .Y(n_717) );
BUFx2_ASAP7_75t_L g782 ( .A(n_443), .Y(n_782) );
BUFx2_ASAP7_75t_SL g835 ( .A(n_443), .Y(n_835) );
AND2x2_ASAP7_75t_L g515 ( .A(n_444), .B(n_516), .Y(n_515) );
INVx3_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx3_ASAP7_75t_L g645 ( .A(n_447), .Y(n_645) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx2_ASAP7_75t_SL g468 ( .A(n_448), .Y(n_468) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_448), .Y(n_507) );
BUFx2_ASAP7_75t_SL g976 ( .A(n_448), .Y(n_976) );
BUFx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
BUFx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_451), .Y(n_514) );
INVx2_ASAP7_75t_L g613 ( .A(n_451), .Y(n_613) );
BUFx3_ASAP7_75t_L g655 ( .A(n_451), .Y(n_655) );
BUFx3_ASAP7_75t_L g723 ( .A(n_451), .Y(n_723) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OAI22xp5_ASAP7_75t_SL g454 ( .A1(n_455), .A2(n_562), .B1(n_563), .B2(n_596), .Y(n_454) );
INVx1_ASAP7_75t_L g596 ( .A(n_455), .Y(n_596) );
AO22x1_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_457), .B1(n_485), .B2(n_486), .Y(n_455) );
INVx1_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
NOR4xp75_ASAP7_75t_L g458 ( .A(n_459), .B(n_466), .C(n_473), .D(n_479), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_460), .B(n_463), .Y(n_459) );
INVx2_ASAP7_75t_L g907 ( .A(n_461), .Y(n_907) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx3_ASAP7_75t_L g607 ( .A(n_462), .Y(n_607) );
INVx2_ASAP7_75t_L g788 ( .A(n_462), .Y(n_788) );
INVx2_ASAP7_75t_L g861 ( .A(n_462), .Y(n_861) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_467), .B(n_471), .Y(n_466) );
INVx4_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_SL g606 ( .A(n_470), .Y(n_606) );
INVx3_ASAP7_75t_L g743 ( .A(n_470), .Y(n_743) );
NOR2xp33_ASAP7_75t_L g980 ( .A(n_470), .B(n_981), .Y(n_980) );
INVx1_ASAP7_75t_L g574 ( .A(n_472), .Y(n_574) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_474), .B(n_477), .Y(n_473) );
BUFx2_ASAP7_75t_L g584 ( .A(n_475), .Y(n_584) );
OAI21xp5_ASAP7_75t_SL g479 ( .A1(n_480), .A2(n_482), .B(n_483), .Y(n_479) );
OAI21xp33_ASAP7_75t_L g848 ( .A1(n_480), .A2(n_849), .B(n_850), .Y(n_848) );
OAI21xp33_ASAP7_75t_SL g895 ( .A1(n_480), .A2(n_896), .B(n_897), .Y(n_895) );
INVx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
BUFx6f_ASAP7_75t_L g592 ( .A(n_484), .Y(n_592) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
XNOR2x1_ASAP7_75t_SL g486 ( .A(n_487), .B(n_518), .Y(n_486) );
INVx3_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
XOR2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_517), .Y(n_489) );
NAND2x1p5_ASAP7_75t_L g490 ( .A(n_491), .B(n_502), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_492), .B(n_497), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_494), .B(n_495), .Y(n_492) );
OAI21xp33_ASAP7_75t_SL g530 ( .A1(n_494), .A2(n_531), .B(n_532), .Y(n_530) );
OAI221xp5_ASAP7_75t_L g822 ( .A1(n_494), .A2(n_823), .B1(n_824), .B2(n_826), .C(n_827), .Y(n_822) );
OAI21xp5_ASAP7_75t_SL g1034 ( .A1(n_494), .A2(n_1035), .B(n_1036), .Y(n_1034) );
BUFx4f_ASAP7_75t_SL g593 ( .A(n_496), .Y(n_593) );
INVx2_ASAP7_75t_L g663 ( .A(n_496), .Y(n_663) );
NAND3xp33_ASAP7_75t_L g497 ( .A(n_498), .B(n_500), .C(n_501), .Y(n_497) );
NOR2x1_ASAP7_75t_L g502 ( .A(n_503), .B(n_509), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_506), .Y(n_503) );
INVx3_ASAP7_75t_L g549 ( .A(n_507), .Y(n_549) );
BUFx3_ASAP7_75t_L g609 ( .A(n_507), .Y(n_609) );
BUFx3_ASAP7_75t_L g709 ( .A(n_507), .Y(n_709) );
BUFx6f_ASAP7_75t_L g786 ( .A(n_507), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_513), .Y(n_509) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_512), .Y(n_615) );
INVx4_ASAP7_75t_L g551 ( .A(n_514), .Y(n_551) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_545), .Y(n_519) );
NOR3xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_530), .C(n_534), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B1(n_526), .B2(n_527), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_523), .A2(n_619), .B1(n_620), .B2(n_621), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_523), .A2(n_528), .B1(n_673), .B2(n_674), .Y(n_672) );
BUFx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_524), .Y(n_693) );
INVx2_ASAP7_75t_L g818 ( .A(n_524), .Y(n_818) );
OAI22xp5_ASAP7_75t_L g845 ( .A1(n_524), .A2(n_621), .B1(n_846), .B2(n_847), .Y(n_845) );
OAI22xp5_ASAP7_75t_SL g890 ( .A1(n_527), .A2(n_891), .B1(n_893), .B2(n_894), .Y(n_890) );
BUFx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OAI22xp5_ASAP7_75t_SL g692 ( .A1(n_528), .A2(n_693), .B1(n_694), .B2(n_695), .Y(n_692) );
INVx2_ASAP7_75t_L g821 ( .A(n_528), .Y(n_821) );
BUFx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g622 ( .A(n_529), .Y(n_622) );
BUFx2_ASAP7_75t_L g661 ( .A(n_533), .Y(n_661) );
INVx4_ASAP7_75t_L g770 ( .A(n_533), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_536), .B1(n_539), .B2(n_540), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_536), .A2(n_630), .B1(n_631), .B2(n_632), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_536), .A2(n_542), .B1(n_736), .B2(n_737), .Y(n_735) );
INVx3_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g587 ( .A(n_537), .Y(n_587) );
INVx4_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_538), .A2(n_542), .B1(n_679), .B2(n_680), .Y(n_678) );
BUFx3_ASAP7_75t_L g703 ( .A(n_538), .Y(n_703) );
HB1xp67_ASAP7_75t_L g830 ( .A(n_538), .Y(n_830) );
OAI22xp33_ASAP7_75t_SL g898 ( .A1(n_538), .A2(n_632), .B1(n_899), .B2(n_900), .Y(n_898) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g632 ( .A(n_541), .Y(n_632) );
CKINVDCx16_ASAP7_75t_R g541 ( .A(n_542), .Y(n_541) );
BUFx2_ASAP7_75t_L g589 ( .A(n_542), .Y(n_589) );
OR2x6_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_546), .B(n_556), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_552), .Y(n_546) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx4_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx3_ASAP7_75t_L g781 ( .A(n_551), .Y(n_781) );
INVx3_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_560), .Y(n_556) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g912 ( .A1(n_559), .A2(n_913), .B1(n_914), .B2(n_915), .Y(n_912) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g595 ( .A(n_564), .Y(n_595) );
AND4x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_575), .C(n_583), .D(n_590), .Y(n_564) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
BUFx2_ASAP7_75t_L g973 ( .A(n_568), .Y(n_973) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_571), .B1(n_573), .B2(n_574), .Y(n_569) );
INVx1_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_578), .B1(n_580), .B2(n_581), .Y(n_576) );
OAI21xp33_ASAP7_75t_L g977 ( .A1(n_578), .A2(n_978), .B(n_979), .Y(n_977) );
BUFx2_ASAP7_75t_R g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .B1(n_588), .B2(n_589), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g851 ( .A1(n_587), .A2(n_852), .B1(n_853), .B2(n_854), .Y(n_851) );
INVx2_ASAP7_75t_SL g697 ( .A(n_592), .Y(n_697) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_666), .B1(n_753), .B2(n_754), .Y(n_598) );
INVx1_ASAP7_75t_L g754 ( .A(n_599), .Y(n_754) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_635), .B1(n_636), .B2(n_665), .Y(n_600) );
INVx1_ASAP7_75t_L g665 ( .A(n_601), .Y(n_665) );
INVx1_ASAP7_75t_SL g634 ( .A(n_602), .Y(n_634) );
AND2x2_ASAP7_75t_SL g602 ( .A(n_603), .B(n_617), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_604), .B(n_610), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_608), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_614), .Y(n_610) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NOR3xp33_ASAP7_75t_L g617 ( .A(n_618), .B(n_623), .C(n_629), .Y(n_617) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g648 ( .A(n_622), .Y(n_648) );
BUFx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
BUFx3_ASAP7_75t_L g825 ( .A(n_628), .Y(n_825) );
OAI22xp5_ASAP7_75t_SL g702 ( .A1(n_632), .A2(n_703), .B1(n_704), .B2(n_705), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g828 ( .A1(n_632), .A2(n_829), .B1(n_830), .B2(n_831), .Y(n_828) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AO22x1_ASAP7_75t_L g725 ( .A1(n_637), .A2(n_638), .B1(n_726), .B2(n_749), .Y(n_725) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
XOR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_664), .Y(n_638) );
NAND4xp75_ASAP7_75t_L g639 ( .A(n_640), .B(n_646), .C(n_653), .D(n_659), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_644), .Y(n_640) );
OA211x2_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_648), .B(n_649), .C(n_651), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_648), .A2(n_693), .B1(n_730), .B2(n_731), .Y(n_729) );
INVx1_ASAP7_75t_SL g778 ( .A(n_652), .Y(n_778) );
AND2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_656), .Y(n_653) );
INVx1_ASAP7_75t_L g914 ( .A(n_655), .Y(n_914) );
INVx2_ASAP7_75t_L g766 ( .A(n_660), .Y(n_766) );
INVx3_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g753 ( .A(n_666), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_687), .B1(n_751), .B2(n_752), .Y(n_666) );
INVx2_ASAP7_75t_SL g751 ( .A(n_667), .Y(n_751) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AND3x1_ASAP7_75t_L g670 ( .A(n_671), .B(n_681), .C(n_684), .Y(n_670) );
NOR3xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_675), .C(n_678), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
AND2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
AND2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
INVx1_ASAP7_75t_L g752 ( .A(n_687), .Y(n_752) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_724), .B1(n_725), .B2(n_750), .Y(n_687) );
INVx2_ASAP7_75t_L g750 ( .A(n_688), .Y(n_750) );
XNOR2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
AND2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_706), .Y(n_690) );
NOR3xp33_ASAP7_75t_L g691 ( .A(n_692), .B(n_696), .C(n_702), .Y(n_691) );
INVx1_ASAP7_75t_L g892 ( .A(n_693), .Y(n_892) );
OAI21xp5_ASAP7_75t_SL g732 ( .A1(n_699), .A2(n_733), .B(n_734), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_707), .B(n_715), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_708), .B(n_710), .Y(n_707) );
INVx3_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
BUFx6f_ASAP7_75t_L g837 ( .A(n_713), .Y(n_837) );
BUFx2_ASAP7_75t_L g1018 ( .A(n_713), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_716), .B(n_718), .Y(n_715) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
BUFx4f_ASAP7_75t_SL g741 ( .A(n_721), .Y(n_741) );
BUFx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g749 ( .A(n_726), .Y(n_749) );
INVx2_ASAP7_75t_L g747 ( .A(n_727), .Y(n_747) );
AND2x2_ASAP7_75t_L g727 ( .A(n_728), .B(n_738), .Y(n_727) );
NOR3xp33_ASAP7_75t_L g728 ( .A(n_729), .B(n_732), .C(n_735), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_744), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_742), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
INVx1_ASAP7_75t_L g986 ( .A(n_755), .Y(n_986) );
XOR2xp5_ASAP7_75t_L g755 ( .A(n_756), .B(n_959), .Y(n_755) );
AOI22xp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_808), .B1(n_957), .B2(n_958), .Y(n_756) );
INVx1_ASAP7_75t_L g957 ( .A(n_757), .Y(n_957) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_759), .B1(n_790), .B2(n_791), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
BUFx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g789 ( .A(n_763), .Y(n_789) );
NAND3x1_ASAP7_75t_L g763 ( .A(n_764), .B(n_779), .C(n_784), .Y(n_763) );
NOR2x1_ASAP7_75t_L g764 ( .A(n_765), .B(n_771), .Y(n_764) );
OAI21xp5_ASAP7_75t_SL g765 ( .A1(n_766), .A2(n_767), .B(n_768), .Y(n_765) );
OAI21xp5_ASAP7_75t_SL g965 ( .A1(n_766), .A2(n_966), .B(n_967), .Y(n_965) );
INVx3_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
NAND3xp33_ASAP7_75t_L g771 ( .A(n_772), .B(n_773), .C(n_774), .Y(n_771) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g805 ( .A(n_776), .Y(n_805) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
AND2x2_ASAP7_75t_L g779 ( .A(n_780), .B(n_783), .Y(n_779) );
AND2x2_ASAP7_75t_L g784 ( .A(n_785), .B(n_787), .Y(n_784) );
INVx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
NAND4xp75_ASAP7_75t_L g792 ( .A(n_793), .B(n_797), .C(n_800), .D(n_806), .Y(n_792) );
AND2x2_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
AND2x2_ASAP7_75t_L g797 ( .A(n_798), .B(n_799), .Y(n_797) );
AND2x2_ASAP7_75t_SL g800 ( .A(n_801), .B(n_804), .Y(n_800) );
INVx1_ASAP7_75t_SL g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_SL g1011 ( .A(n_803), .Y(n_1011) );
INVx1_ASAP7_75t_L g853 ( .A(n_807), .Y(n_853) );
INVx1_ASAP7_75t_L g958 ( .A(n_808), .Y(n_958) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
AOI22xp5_ASAP7_75t_L g810 ( .A1(n_811), .A2(n_884), .B1(n_955), .B2(n_956), .Y(n_810) );
INVx2_ASAP7_75t_L g955 ( .A(n_811), .Y(n_955) );
OA22x2_ASAP7_75t_L g811 ( .A1(n_812), .A2(n_841), .B1(n_882), .B2(n_883), .Y(n_811) );
INVx2_ASAP7_75t_L g882 ( .A(n_812), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_814), .B(n_832), .Y(n_813) );
NOR3xp33_ASAP7_75t_L g814 ( .A(n_815), .B(n_822), .C(n_828), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_816), .A2(n_817), .B1(n_819), .B2(n_820), .Y(n_815) );
INVx2_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_833), .B(n_838), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_834), .B(n_836), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_839), .B(n_840), .Y(n_838) );
INVx2_ASAP7_75t_L g883 ( .A(n_841), .Y(n_883) );
XOR2x2_ASAP7_75t_L g841 ( .A(n_842), .B(n_863), .Y(n_841) );
AND2x2_ASAP7_75t_L g843 ( .A(n_844), .B(n_855), .Y(n_843) );
NOR3xp33_ASAP7_75t_L g844 ( .A(n_845), .B(n_848), .C(n_851), .Y(n_844) );
NOR2xp33_ASAP7_75t_L g855 ( .A(n_856), .B(n_859), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_857), .B(n_858), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_860), .B(n_862), .Y(n_859) );
INVx2_ASAP7_75t_L g982 ( .A(n_863), .Y(n_982) );
XOR2x2_ASAP7_75t_L g863 ( .A(n_864), .B(n_881), .Y(n_863) );
NAND3x1_ASAP7_75t_L g864 ( .A(n_865), .B(n_868), .C(n_877), .Y(n_864) );
AND2x2_ASAP7_75t_L g865 ( .A(n_866), .B(n_867), .Y(n_865) );
NOR2x1_ASAP7_75t_L g868 ( .A(n_869), .B(n_872), .Y(n_868) );
NAND3xp33_ASAP7_75t_L g872 ( .A(n_873), .B(n_874), .C(n_875), .Y(n_872) );
AND2x2_ASAP7_75t_L g877 ( .A(n_878), .B(n_880), .Y(n_877) );
INVx1_ASAP7_75t_L g956 ( .A(n_884), .Y(n_956) );
XNOR2x2_ASAP7_75t_L g884 ( .A(n_885), .B(n_916), .Y(n_884) );
INVx2_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
AND2x2_ASAP7_75t_L g888 ( .A(n_889), .B(n_901), .Y(n_888) );
NOR3xp33_ASAP7_75t_L g889 ( .A(n_890), .B(n_895), .C(n_898), .Y(n_889) );
INVx2_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
NOR3xp33_ASAP7_75t_L g901 ( .A(n_902), .B(n_905), .C(n_912), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_903), .B(n_904), .Y(n_902) );
OAI22xp5_ASAP7_75t_L g905 ( .A1(n_906), .A2(n_907), .B1(n_908), .B2(n_909), .Y(n_905) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
OAI22x1_ASAP7_75t_L g916 ( .A1(n_917), .A2(n_936), .B1(n_937), .B2(n_954), .Y(n_916) );
INVx2_ASAP7_75t_L g954 ( .A(n_917), .Y(n_954) );
AND2x4_ASAP7_75t_L g918 ( .A(n_919), .B(n_929), .Y(n_918) );
NOR2xp33_ASAP7_75t_L g919 ( .A(n_920), .B(n_924), .Y(n_919) );
NAND3xp33_ASAP7_75t_L g924 ( .A(n_925), .B(n_926), .C(n_927), .Y(n_924) );
NOR2x1_ASAP7_75t_L g929 ( .A(n_930), .B(n_933), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_931), .B(n_932), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_934), .B(n_935), .Y(n_933) );
INVx3_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
XOR2x2_ASAP7_75t_L g937 ( .A(n_938), .B(n_953), .Y(n_937) );
NAND3x1_ASAP7_75t_SL g938 ( .A(n_939), .B(n_942), .C(n_950), .Y(n_938) );
AND2x2_ASAP7_75t_L g939 ( .A(n_940), .B(n_941), .Y(n_939) );
NOR2x1_ASAP7_75t_L g942 ( .A(n_943), .B(n_946), .Y(n_942) );
NAND3xp33_ASAP7_75t_L g946 ( .A(n_947), .B(n_948), .C(n_949), .Y(n_946) );
AND2x2_ASAP7_75t_L g950 ( .A(n_951), .B(n_952), .Y(n_950) );
INVx1_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
INVx1_ASAP7_75t_SL g960 ( .A(n_961), .Y(n_960) );
OAI22x1_ASAP7_75t_L g961 ( .A1(n_962), .A2(n_982), .B1(n_983), .B2(n_984), .Y(n_961) );
INVx1_ASAP7_75t_L g983 ( .A(n_962), .Y(n_983) );
NAND3x1_ASAP7_75t_L g963 ( .A(n_964), .B(n_971), .C(n_975), .Y(n_963) );
NOR2xp33_ASAP7_75t_L g964 ( .A(n_965), .B(n_968), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g968 ( .A(n_969), .B(n_970), .Y(n_968) );
AND2x2_ASAP7_75t_L g971 ( .A(n_972), .B(n_974), .Y(n_971) );
INVx1_ASAP7_75t_L g984 ( .A(n_982), .Y(n_984) );
INVx1_ASAP7_75t_SL g987 ( .A(n_988), .Y(n_987) );
NOR2x1_ASAP7_75t_L g988 ( .A(n_989), .B(n_993), .Y(n_988) );
OR2x2_ASAP7_75t_SL g1049 ( .A(n_989), .B(n_994), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_990), .B(n_992), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
OAI322xp33_ASAP7_75t_L g1000 ( .A1(n_991), .A2(n_1001), .A3(n_1023), .B1(n_1025), .B2(n_1028), .C1(n_1029), .C2(n_1047), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_991), .B(n_1024), .Y(n_1027) );
CKINVDCx16_ASAP7_75t_R g1024 ( .A(n_992), .Y(n_1024) );
CKINVDCx20_ASAP7_75t_R g993 ( .A(n_994), .Y(n_993) );
NAND2xp5_ASAP7_75t_L g994 ( .A(n_995), .B(n_996), .Y(n_994) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_998), .B(n_999), .Y(n_997) );
CKINVDCx14_ASAP7_75t_R g1002 ( .A(n_1003), .Y(n_1002) );
HB1xp67_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
NAND3x1_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1015), .C(n_1019), .Y(n_1004) );
NOR2x1_ASAP7_75t_L g1005 ( .A(n_1006), .B(n_1009), .Y(n_1005) );
NAND3xp33_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1012), .C(n_1013), .Y(n_1009) );
AND2x2_ASAP7_75t_L g1015 ( .A(n_1016), .B(n_1017), .Y(n_1015) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_1020), .B(n_1021), .Y(n_1019) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
CKINVDCx16_ASAP7_75t_R g1025 ( .A(n_1026), .Y(n_1025) );
XOR2x2_ASAP7_75t_L g1031 ( .A(n_1028), .B(n_1032), .Y(n_1031) );
INVx1_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
NAND3x1_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1041), .C(n_1044), .Y(n_1032) );
NOR2xp33_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1037), .Y(n_1033) );
NAND3xp33_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1039), .C(n_1040), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1043), .Y(n_1041) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_1045), .B(n_1046), .Y(n_1044) );
CKINVDCx20_ASAP7_75t_R g1047 ( .A(n_1048), .Y(n_1047) );
CKINVDCx20_ASAP7_75t_R g1048 ( .A(n_1049), .Y(n_1048) );
endmodule