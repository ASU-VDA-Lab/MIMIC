module fake_netlist_6_4587_n_3374 (n_52, n_591, n_435, n_1, n_91, n_793, n_326, n_801, n_256, n_853, n_440, n_587, n_695, n_507, n_580, n_762, n_209, n_367, n_465, n_680, n_741, n_760, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_828, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_740, n_578, n_703, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_820, n_783, n_106, n_725, n_358, n_160, n_751, n_449, n_131, n_749, n_798, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_805, n_396, n_495, n_815, n_350, n_78, n_84, n_585, n_732, n_568, n_392, n_840, n_442, n_480, n_142, n_724, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_823, n_349, n_643, n_233, n_617, n_698, n_845, n_255, n_807, n_739, n_284, n_400, n_140, n_337, n_865, n_214, n_485, n_67, n_15, n_443, n_246, n_768, n_38, n_471, n_289, n_421, n_781, n_424, n_789, n_615, n_59, n_181, n_182, n_238, n_573, n_769, n_202, n_320, n_108, n_639, n_676, n_327, n_794, n_727, n_369, n_597, n_685, n_280, n_287, n_832, n_353, n_610, n_555, n_389, n_814, n_415, n_830, n_65, n_230, n_605, n_461, n_141, n_383, n_826, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_747, n_852, n_667, n_71, n_74, n_229, n_542, n_847, n_644, n_682, n_851, n_621, n_305, n_72, n_721, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_791, n_35, n_183, n_510, n_837, n_836, n_79, n_863, n_375, n_601, n_338, n_522, n_466, n_704, n_748, n_506, n_56, n_763, n_360, n_603, n_119, n_235, n_536, n_866, n_622, n_147, n_191, n_340, n_710, n_387, n_452, n_616, n_658, n_744, n_39, n_344, n_73, n_581, n_428, n_761, n_785, n_746, n_609, n_765, n_432, n_641, n_822, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_758, n_842, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_772, n_96, n_8, n_843, n_797, n_666, n_371, n_795, n_770, n_567, n_189, n_738, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_838, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_844, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_752, n_112, n_172, n_713, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_782, n_490, n_803, n_290, n_220, n_809, n_118, n_224, n_48, n_25, n_93, n_839, n_80, n_734, n_708, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_779, n_9, n_800, n_460, n_107, n_854, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_366, n_777, n_407, n_450, n_103, n_808, n_272, n_526, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_717, n_46, n_330, n_771, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_824, n_279, n_686, n_796, n_252, n_757, n_228, n_565, n_594, n_719, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_813, n_592, n_745, n_654, n_323, n_829, n_606, n_393, n_818, n_411, n_503, n_716, n_152, n_623, n_92, n_599, n_513, n_855, n_776, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_731, n_859, n_406, n_483, n_735, n_102, n_204, n_482, n_755, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_792, n_476, n_714, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_860, n_481, n_788, n_819, n_821, n_325, n_767, n_804, n_329, n_464, n_600, n_831, n_802, n_561, n_33, n_477, n_549, n_533, n_408, n_806, n_864, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_833, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_345, n_409, n_231, n_354, n_689, n_40, n_799, n_505, n_240, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_810, n_635, n_95, n_787, n_311, n_10, n_403, n_723, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_764, n_556, n_159, n_157, n_162, n_692, n_733, n_754, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_849, n_560, n_753, n_642, n_276, n_569, n_441, n_221, n_811, n_444, n_586, n_423, n_146, n_737, n_318, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_790, n_582, n_4, n_199, n_138, n_266, n_296, n_861, n_674, n_857, n_775, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_759, n_355, n_426, n_317, n_149, n_632, n_702, n_431, n_90, n_347, n_812, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_780, n_773, n_675, n_85, n_99, n_257, n_730, n_655, n_13, n_706, n_786, n_670, n_203, n_286, n_254, n_207, n_834, n_242, n_835, n_19, n_47, n_690, n_29, n_850, n_75, n_401, n_324, n_743, n_766, n_816, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_848, n_120, n_251, n_301, n_274, n_636, n_825, n_728, n_681, n_729, n_110, n_151, n_774, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_784, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_688, n_722, n_862, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_637, n_295, n_385, n_701, n_817, n_629, n_388, n_190, n_858, n_262, n_484, n_613, n_736, n_187, n_846, n_501, n_841, n_531, n_827, n_60, n_361, n_508, n_663, n_856, n_379, n_170, n_778, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_3374);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_793;
input n_326;
input n_801;
input n_256;
input n_853;
input n_440;
input n_587;
input n_695;
input n_507;
input n_580;
input n_762;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_760;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_828;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_740;
input n_578;
input n_703;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_820;
input n_783;
input n_106;
input n_725;
input n_358;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_798;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_805;
input n_396;
input n_495;
input n_815;
input n_350;
input n_78;
input n_84;
input n_585;
input n_732;
input n_568;
input n_392;
input n_840;
input n_442;
input n_480;
input n_142;
input n_724;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_823;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_845;
input n_255;
input n_807;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_865;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_768;
input n_38;
input n_471;
input n_289;
input n_421;
input n_781;
input n_424;
input n_789;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_769;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_794;
input n_727;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_832;
input n_353;
input n_610;
input n_555;
input n_389;
input n_814;
input n_415;
input n_830;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_826;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_747;
input n_852;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_621;
input n_305;
input n_72;
input n_721;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_791;
input n_35;
input n_183;
input n_510;
input n_837;
input n_836;
input n_79;
input n_863;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_704;
input n_748;
input n_506;
input n_56;
input n_763;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_866;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_387;
input n_452;
input n_616;
input n_658;
input n_744;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_761;
input n_785;
input n_746;
input n_609;
input n_765;
input n_432;
input n_641;
input n_822;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_758;
input n_842;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_772;
input n_96;
input n_8;
input n_843;
input n_797;
input n_666;
input n_371;
input n_795;
input n_770;
input n_567;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_838;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_844;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_752;
input n_112;
input n_172;
input n_713;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_782;
input n_490;
input n_803;
input n_290;
input n_220;
input n_809;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_839;
input n_80;
input n_734;
input n_708;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_779;
input n_9;
input n_800;
input n_460;
input n_107;
input n_854;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_366;
input n_777;
input n_407;
input n_450;
input n_103;
input n_808;
input n_272;
input n_526;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_717;
input n_46;
input n_330;
input n_771;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_824;
input n_279;
input n_686;
input n_796;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_813;
input n_592;
input n_745;
input n_654;
input n_323;
input n_829;
input n_606;
input n_393;
input n_818;
input n_411;
input n_503;
input n_716;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_855;
input n_776;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_731;
input n_859;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_755;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_792;
input n_476;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_860;
input n_481;
input n_788;
input n_819;
input n_821;
input n_325;
input n_767;
input n_804;
input n_329;
input n_464;
input n_600;
input n_831;
input n_802;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_806;
input n_864;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_833;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_799;
input n_505;
input n_240;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_810;
input n_635;
input n_95;
input n_787;
input n_311;
input n_10;
input n_403;
input n_723;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_764;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_733;
input n_754;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_849;
input n_560;
input n_753;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_811;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_790;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_861;
input n_674;
input n_857;
input n_775;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_759;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_812;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_780;
input n_773;
input n_675;
input n_85;
input n_99;
input n_257;
input n_730;
input n_655;
input n_13;
input n_706;
input n_786;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_834;
input n_242;
input n_835;
input n_19;
input n_47;
input n_690;
input n_29;
input n_850;
input n_75;
input n_401;
input n_324;
input n_743;
input n_766;
input n_816;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_848;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_825;
input n_728;
input n_681;
input n_729;
input n_110;
input n_151;
input n_774;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_784;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_688;
input n_722;
input n_862;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_637;
input n_295;
input n_385;
input n_701;
input n_817;
input n_629;
input n_388;
input n_190;
input n_858;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_846;
input n_501;
input n_841;
input n_531;
input n_827;
input n_60;
input n_361;
input n_508;
input n_663;
input n_856;
input n_379;
input n_170;
input n_778;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_3374;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_1613;
wire n_1458;
wire n_1234;
wire n_2576;
wire n_3254;
wire n_1674;
wire n_1199;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_1189;
wire n_3152;
wire n_1212;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_1357;
wire n_1853;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_3088;
wire n_1923;
wire n_3257;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_1708;
wire n_1151;
wire n_2977;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_3332;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_3030;
wire n_2291;
wire n_2299;
wire n_3340;
wire n_873;
wire n_1371;
wire n_1285;
wire n_2886;
wire n_2974;
wire n_1985;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_1172;
wire n_2509;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_3345;
wire n_2074;
wire n_2447;
wire n_2919;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1772;
wire n_1232;
wire n_1572;
wire n_1874;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_2480;
wire n_2739;
wire n_3023;
wire n_3232;
wire n_1313;
wire n_2791;
wire n_3251;
wire n_1056;
wire n_3316;
wire n_2212;
wire n_3063;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3048;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_940;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_3028;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3077;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3107;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_2836;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_1467;
wire n_3297;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_2085;
wire n_3368;
wire n_917;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_913;
wire n_1658;
wire n_2593;
wire n_867;
wire n_3269;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_1986;
wire n_2397;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2907;
wire n_2735;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_2850;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_3373;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_1381;
wire n_2961;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_2669;
wire n_2925;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_2522;
wire n_2792;
wire n_1328;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_3118;
wire n_3315;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_1530;
wire n_939;
wire n_1543;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1599;
wire n_1068;
wire n_982;
wire n_2674;
wire n_2832;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_2831;
wire n_2998;
wire n_3317;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_2455;
wire n_2876;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_2355;
wire n_966;
wire n_2908;
wire n_3168;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_1793;
wire n_2922;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_3092;
wire n_3055;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_3294;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_2459;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_3369;
wire n_1982;
wire n_2878;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3247;
wire n_871;
wire n_3069;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_1165;
wire n_2749;
wire n_2008;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_2254;
wire n_3346;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_928;
wire n_1801;
wire n_1214;
wire n_2347;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_1157;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3153;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_2916;
wire n_1063;
wire n_1588;
wire n_2963;
wire n_2947;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_2980;
wire n_1965;
wire n_2476;
wire n_3280;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_890;
wire n_2377;
wire n_3271;
wire n_2178;
wire n_950;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_2887;
wire n_2075;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_2431;
wire n_3073;
wire n_2987;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_2078;
wire n_1634;
wire n_3252;
wire n_2932;
wire n_1767;
wire n_3253;
wire n_1779;
wire n_1465;
wire n_3337;
wire n_3209;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_2893;
wire n_1627;
wire n_1164;
wire n_1295;
wire n_2954;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_2913;
wire n_874;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_3366;
wire n_2631;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_963;
wire n_2767;
wire n_894;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_2707;
wire n_3240;
wire n_1514;
wire n_1863;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_872;
wire n_1139;
wire n_1714;
wire n_3179;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_2537;
wire n_2897;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_3171;
wire n_1913;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_3158;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_2590;
wire n_2643;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_1492;
wire n_987;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_3104;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_1432;
wire n_2208;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_1809;
wire n_3119;
wire n_2958;
wire n_1577;
wire n_2948;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_2936;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1448;
wire n_1087;
wire n_3173;
wire n_1992;
wire n_1049;
wire n_3223;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_3129;
wire n_1849;
wire n_2848;
wire n_919;
wire n_2868;
wire n_1698;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_1299;
wire n_2896;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_998;
wire n_3200;
wire n_1665;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_2338;
wire n_1424;
wire n_3324;
wire n_3341;
wire n_1073;
wire n_1000;
wire n_1195;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_1507;
wire n_2482;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3006;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_3201;
wire n_1142;
wire n_2849;
wire n_1475;
wire n_1048;
wire n_1398;
wire n_1774;
wire n_884;
wire n_1201;
wire n_2354;
wire n_2682;
wire n_3032;
wire n_3103;
wire n_2589;
wire n_1395;
wire n_2199;
wire n_2110;
wire n_2661;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_1021;
wire n_931;
wire n_1207;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_3331;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3087;
wire n_3072;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_889;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_1310;
wire n_3142;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_1837;
wire n_964;
wire n_1314;
wire n_2218;
wire n_2788;
wire n_3196;
wire n_2435;
wire n_954;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_3327;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_1877;
wire n_3144;
wire n_3211;
wire n_3244;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2784;
wire n_2301;
wire n_2209;
wire n_3287;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_970;
wire n_3306;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_3033;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_1223;
wire n_2990;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3226;
wire n_3323;
wire n_3364;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_914;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_2920;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_3188;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_3243;
wire n_1617;
wire n_3260;
wire n_3370;
wire n_1470;
wire n_2550;
wire n_3093;
wire n_3175;
wire n_3214;
wire n_1243;
wire n_2732;
wire n_2928;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_3284;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_1390;
wire n_906;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_2863;
wire n_3299;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_3360;
wire n_2135;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_2049;
wire n_1331;
wire n_2627;
wire n_956;
wire n_960;
wire n_2276;
wire n_3234;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3016;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_2993;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_1129;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_1869;
wire n_2911;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_1593;
wire n_1202;
wire n_1030;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_2942;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_2555;
wire n_3338;
wire n_2219;
wire n_1203;
wire n_2851;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_999;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_2984;
wire n_994;
wire n_2263;
wire n_3291;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3194;
wire n_3250;
wire n_1934;
wire n_3276;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_1871;
wire n_2924;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_1510;
wire n_892;
wire n_3120;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_2302;
wire n_1667;
wire n_1206;
wire n_3230;
wire n_1037;
wire n_1397;
wire n_3268;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_901;
wire n_1499;
wire n_2755;
wire n_3141;
wire n_923;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_3131;
wire n_2439;
wire n_1108;
wire n_1818;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_2740;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_3213;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3010;
wire n_2499;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_2486;
wire n_3132;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3238;
wire n_2235;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_1043;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_2964;
wire n_1692;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_1840;
wire n_1152;
wire n_1705;
wire n_3262;
wire n_2904;
wire n_2244;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_1405;
wire n_972;
wire n_2376;
wire n_1406;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_962;
wire n_1041;
wire n_2346;
wire n_3134;
wire n_1569;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_1288;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_2882;
wire n_3320;
wire n_2541;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2871;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_1846;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_2390;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_2986;
wire n_1900;
wire n_3246;
wire n_1548;
wire n_3044;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_2172;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2154;
wire n_2727;
wire n_2962;
wire n_2939;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_2533;
wire n_3157;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2945;
wire n_3061;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_2427;
wire n_3151;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_1706;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3156;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_2668;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_1650;
wire n_1794;
wire n_1045;
wire n_1962;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_3091;
wire n_2695;
wire n_3124;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_2671;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2923;
wire n_1804;
wire n_2888;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_2054;
wire n_876;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_3308;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_1098;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_1150;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1076;
wire n_1118;
wire n_2949;
wire n_1807;
wire n_1007;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_875;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_1953;
wire n_933;
wire n_3343;
wire n_3303;
wire n_978;
wire n_2752;
wire n_3135;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3034;
wire n_1132;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2969;
wire n_1338;
wire n_1097;
wire n_2787;
wire n_2395;
wire n_935;
wire n_3027;
wire n_1554;
wire n_3231;
wire n_1130;
wire n_3083;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_2380;
wire n_1120;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_1461;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_2935;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_918;
wire n_1848;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_971;
wire n_2702;
wire n_3241;
wire n_946;
wire n_2906;
wire n_1303;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_1689;
wire n_2180;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_1501;
wire n_1221;
wire n_3334;
wire n_1245;
wire n_3215;
wire n_3336;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_1561;
wire n_2741;
wire n_3114;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_2437;
wire n_2743;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3035;
wire n_990;
wire n_1500;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_3204;
wire n_1104;
wire n_1058;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_2242;
wire n_3362;
wire n_1509;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3290;
wire n_1109;
wire n_2222;
wire n_3256;
wire n_1276;
wire n_3176;
wire n_3309;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_2999;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_1584;
wire n_2425;
wire n_924;
wire n_1582;
wire n_2318;
wire n_3286;
wire n_2408;
wire n_1149;
wire n_3170;
wire n_1184;
wire n_2483;
wire n_2950;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_2592;
wire n_1525;
wire n_3098;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_1362;
wire n_1156;
wire n_3123;
wire n_2600;
wire n_984;
wire n_1829;
wire n_2035;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_868;
wire n_3038;
wire n_3086;
wire n_2033;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_3285;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_3361;
wire n_981;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_3344;
wire n_2334;
wire n_3295;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_1133;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_1996;
wire n_2367;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_941;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_2662;
wire n_3147;
wire n_3116;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3359;
wire n_2795;
wire n_2471;
wire n_3187;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_2065;
wire n_2879;
wire n_967;
wire n_2461;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_2968;
wire n_1170;
wire n_1629;
wire n_2221;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3001;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2185;
wire n_2086;
wire n_2927;
wire n_1836;
wire n_2774;
wire n_3039;
wire n_1226;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3274;
wire n_3333;
wire n_3186;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_2579;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_3085;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_3070;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_2991;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_1742;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g867 ( 
.A(n_131),
.Y(n_867)
);

CKINVDCx20_ASAP7_75t_R g868 ( 
.A(n_25),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_706),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_718),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_166),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_502),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_804),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_613),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_657),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_468),
.Y(n_876)
);

CKINVDCx20_ASAP7_75t_R g877 ( 
.A(n_396),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_499),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_713),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_22),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_293),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_664),
.Y(n_882)
);

BUFx2_ASAP7_75t_L g883 ( 
.A(n_161),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_290),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_790),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_8),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_16),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_709),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_119),
.Y(n_889)
);

BUFx2_ASAP7_75t_L g890 ( 
.A(n_478),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_731),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_582),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_407),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_548),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_365),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_769),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_271),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_801),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_811),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_684),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_32),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_845),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_64),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_747),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_467),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_863),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_854),
.Y(n_907)
);

INVx1_ASAP7_75t_SL g908 ( 
.A(n_308),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_626),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_735),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_749),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_252),
.Y(n_912)
);

BUFx10_ASAP7_75t_L g913 ( 
.A(n_802),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_662),
.Y(n_914)
);

INVx1_ASAP7_75t_SL g915 ( 
.A(n_281),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_671),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_610),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_645),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_734),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_711),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_565),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_682),
.Y(n_922)
);

BUFx10_ASAP7_75t_L g923 ( 
.A(n_755),
.Y(n_923)
);

BUFx6f_ASAP7_75t_L g924 ( 
.A(n_720),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_779),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_783),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_634),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_770),
.Y(n_928)
);

INVx1_ASAP7_75t_SL g929 ( 
.A(n_581),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_598),
.Y(n_930)
);

BUFx10_ASAP7_75t_L g931 ( 
.A(n_531),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_647),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_252),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_39),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_700),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_746),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_737),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_202),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_781),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_289),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_377),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_419),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_754),
.Y(n_943)
);

INVxp67_ASAP7_75t_L g944 ( 
.A(n_778),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_475),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_750),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_712),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_589),
.Y(n_948)
);

CKINVDCx20_ASAP7_75t_R g949 ( 
.A(n_786),
.Y(n_949)
);

INVx2_ASAP7_75t_SL g950 ( 
.A(n_696),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_674),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_439),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_837),
.Y(n_953)
);

INVx2_ASAP7_75t_SL g954 ( 
.A(n_6),
.Y(n_954)
);

CKINVDCx20_ASAP7_75t_R g955 ( 
.A(n_727),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_794),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_176),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_814),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_470),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_81),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_477),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_833),
.Y(n_962)
);

INVx2_ASAP7_75t_SL g963 ( 
.A(n_406),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_694),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_846),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_198),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_86),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_839),
.Y(n_968)
);

INVx1_ASAP7_75t_SL g969 ( 
.A(n_793),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_602),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_319),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_453),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_788),
.Y(n_973)
);

BUFx10_ASAP7_75t_L g974 ( 
.A(n_50),
.Y(n_974)
);

CKINVDCx20_ASAP7_75t_R g975 ( 
.A(n_250),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_704),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_194),
.Y(n_977)
);

INVxp67_ASAP7_75t_L g978 ( 
.A(n_740),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_276),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_623),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_400),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_812),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_745),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_726),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_772),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_821),
.Y(n_986)
);

CKINVDCx16_ASAP7_75t_R g987 ( 
.A(n_29),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_305),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_417),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_795),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_497),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_367),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_459),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_798),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_228),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_293),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_660),
.Y(n_997)
);

CKINVDCx20_ASAP7_75t_R g998 ( 
.A(n_784),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_653),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_789),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_153),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_338),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_30),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_341),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_632),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_659),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_600),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_842),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_715),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_64),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_447),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_77),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_114),
.Y(n_1013)
);

INVx1_ASAP7_75t_SL g1014 ( 
.A(n_10),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_752),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_445),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_337),
.Y(n_1017)
);

CKINVDCx20_ASAP7_75t_R g1018 ( 
.A(n_725),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_775),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_708),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_188),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_809),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_69),
.Y(n_1023)
);

BUFx2_ASAP7_75t_L g1024 ( 
.A(n_434),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_312),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_486),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_655),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_590),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_285),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_817),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_862),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_763),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_774),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_583),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_678),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_188),
.Y(n_1036)
);

CKINVDCx20_ASAP7_75t_R g1037 ( 
.A(n_855),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_768),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_787),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_354),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_776),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_572),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_270),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_803),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_608),
.Y(n_1045)
);

HB1xp67_ASAP7_75t_L g1046 ( 
.A(n_587),
.Y(n_1046)
);

BUFx3_ASAP7_75t_L g1047 ( 
.A(n_314),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_239),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_847),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_744),
.Y(n_1050)
);

BUFx5_ASAP7_75t_L g1051 ( 
.A(n_675),
.Y(n_1051)
);

CKINVDCx20_ASAP7_75t_R g1052 ( 
.A(n_157),
.Y(n_1052)
);

INVxp67_ASAP7_75t_L g1053 ( 
.A(n_515),
.Y(n_1053)
);

CKINVDCx20_ASAP7_75t_R g1054 ( 
.A(n_630),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_17),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_651),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_37),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_586),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_688),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_368),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_665),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_810),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_361),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_513),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_765),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_685),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_120),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_618),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_386),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_705),
.Y(n_1070)
);

INVx1_ASAP7_75t_SL g1071 ( 
.A(n_180),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_160),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_308),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_454),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_93),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_523),
.Y(n_1076)
);

CKINVDCx20_ASAP7_75t_R g1077 ( 
.A(n_807),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_306),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_3),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_2),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_510),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_411),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_416),
.Y(n_1083)
);

CKINVDCx20_ASAP7_75t_R g1084 ( 
.A(n_648),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_301),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_782),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_697),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_819),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_346),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_140),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_683),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_656),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_743),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_730),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_851),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_271),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_840),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_693),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_691),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_796),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_155),
.Y(n_1101)
);

BUFx10_ASAP7_75t_L g1102 ( 
.A(n_800),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_161),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_4),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_46),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_208),
.Y(n_1106)
);

BUFx2_ASAP7_75t_SL g1107 ( 
.A(n_434),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_442),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_805),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_835),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_409),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_654),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_698),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_738),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_741),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_736),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_733),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_505),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_672),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_264),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_336),
.Y(n_1121)
);

CKINVDCx20_ASAP7_75t_R g1122 ( 
.A(n_561),
.Y(n_1122)
);

CKINVDCx20_ASAP7_75t_R g1123 ( 
.A(n_238),
.Y(n_1123)
);

INVx1_ASAP7_75t_SL g1124 ( 
.A(n_268),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_767),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_680),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_29),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_751),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_822),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_661),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_392),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_834),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_780),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_826),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_667),
.Y(n_1135)
);

CKINVDCx14_ASAP7_75t_R g1136 ( 
.A(n_838),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_274),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_666),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_76),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_853),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_646),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_732),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_32),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_412),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_841),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_719),
.Y(n_1146)
);

CKINVDCx20_ASAP7_75t_R g1147 ( 
.A(n_454),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_729),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_758),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_761),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_714),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_836),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_507),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_686),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_384),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_766),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_205),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_431),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_325),
.Y(n_1159)
);

INVx1_ASAP7_75t_SL g1160 ( 
.A(n_823),
.Y(n_1160)
);

INVx1_ASAP7_75t_SL g1161 ( 
.A(n_728),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_690),
.Y(n_1162)
);

CKINVDCx20_ASAP7_75t_R g1163 ( 
.A(n_773),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_866),
.Y(n_1164)
);

INVx1_ASAP7_75t_SL g1165 ( 
.A(n_861),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_559),
.Y(n_1166)
);

CKINVDCx20_ASAP7_75t_R g1167 ( 
.A(n_627),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_22),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_156),
.Y(n_1169)
);

CKINVDCx16_ASAP7_75t_R g1170 ( 
.A(n_830),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_721),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_816),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_707),
.Y(n_1173)
);

CKINVDCx16_ASAP7_75t_R g1174 ( 
.A(n_172),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_673),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_844),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_771),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_423),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_827),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_92),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_85),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_831),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_100),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_44),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_6),
.Y(n_1185)
);

INVx1_ASAP7_75t_SL g1186 ( 
.A(n_628),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_860),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_756),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_485),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_815),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_663),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_133),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_143),
.Y(n_1193)
);

CKINVDCx20_ASAP7_75t_R g1194 ( 
.A(n_791),
.Y(n_1194)
);

CKINVDCx20_ASAP7_75t_R g1195 ( 
.A(n_37),
.Y(n_1195)
);

BUFx10_ASAP7_75t_L g1196 ( 
.A(n_402),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_649),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_759),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_650),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_437),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_820),
.Y(n_1201)
);

HB1xp67_ASAP7_75t_L g1202 ( 
.A(n_326),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_273),
.Y(n_1203)
);

CKINVDCx20_ASAP7_75t_R g1204 ( 
.A(n_702),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_445),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_615),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_824),
.Y(n_1207)
);

INVx1_ASAP7_75t_SL g1208 ( 
.A(n_554),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_21),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_383),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_762),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_677),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_742),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_597),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_303),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_10),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_593),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_692),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_174),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_624),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_828),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_757),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_825),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_80),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_524),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_658),
.Y(n_1226)
);

INVxp67_ASAP7_75t_L g1227 ( 
.A(n_202),
.Y(n_1227)
);

BUFx10_ASAP7_75t_L g1228 ( 
.A(n_147),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_724),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_563),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_123),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_575),
.Y(n_1232)
);

CKINVDCx20_ASAP7_75t_R g1233 ( 
.A(n_799),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_430),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_813),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_695),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_777),
.Y(n_1237)
);

INVx1_ASAP7_75t_SL g1238 ( 
.A(n_722),
.Y(n_1238)
);

BUFx3_ASAP7_75t_L g1239 ( 
.A(n_377),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_392),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_348),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_723),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_703),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_641),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_263),
.Y(n_1245)
);

BUFx3_ASAP7_75t_L g1246 ( 
.A(n_278),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_16),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_187),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_760),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_351),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_710),
.Y(n_1251)
);

INVx4_ASAP7_75t_R g1252 ( 
.A(n_681),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_509),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_319),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_288),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_519),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_385),
.Y(n_1257)
);

BUFx10_ASAP7_75t_L g1258 ( 
.A(n_164),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_806),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_858),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_140),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_195),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_138),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_764),
.Y(n_1264)
);

CKINVDCx16_ASAP7_75t_R g1265 ( 
.A(n_429),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_251),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_829),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_70),
.Y(n_1268)
);

CKINVDCx14_ASAP7_75t_R g1269 ( 
.A(n_114),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_184),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_194),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_850),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_376),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_687),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_636),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_832),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_8),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_748),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_325),
.Y(n_1279)
);

BUFx8_ASAP7_75t_SL g1280 ( 
.A(n_753),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_859),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_379),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_180),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_135),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_346),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_716),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_701),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_849),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_689),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_852),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_401),
.Y(n_1291)
);

CKINVDCx20_ASAP7_75t_R g1292 ( 
.A(n_739),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_808),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_635),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_13),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_797),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_676),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_848),
.Y(n_1298)
);

INVx2_ASAP7_75t_SL g1299 ( 
.A(n_395),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_668),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_87),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_355),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_294),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_479),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_843),
.Y(n_1305)
);

BUFx8_ASAP7_75t_SL g1306 ( 
.A(n_669),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_679),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_181),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_670),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_699),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_785),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_652),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_374),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_717),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_792),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_580),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_127),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_360),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_338),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_818),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_535),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_145),
.Y(n_1322)
);

BUFx10_ASAP7_75t_L g1323 ( 
.A(n_316),
.Y(n_1323)
);

INVxp67_ASAP7_75t_SL g1324 ( 
.A(n_980),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1284),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1284),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1074),
.Y(n_1327)
);

BUFx2_ASAP7_75t_L g1328 ( 
.A(n_883),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1280),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1074),
.Y(n_1330)
);

INVxp67_ASAP7_75t_L g1331 ( 
.A(n_1024),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1306),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1074),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1090),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1090),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1090),
.Y(n_1336)
);

INVxp33_ASAP7_75t_SL g1337 ( 
.A(n_1202),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1271),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_870),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_900),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1271),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_913),
.Y(n_1342)
);

CKINVDCx14_ASAP7_75t_R g1343 ( 
.A(n_1269),
.Y(n_1343)
);

INVxp67_ASAP7_75t_SL g1344 ( 
.A(n_1033),
.Y(n_1344)
);

CKINVDCx20_ASAP7_75t_R g1345 ( 
.A(n_949),
.Y(n_1345)
);

BUFx3_ASAP7_75t_L g1346 ( 
.A(n_913),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1271),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_873),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_933),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_988),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_874),
.Y(n_1351)
);

INVx1_ASAP7_75t_SL g1352 ( 
.A(n_1078),
.Y(n_1352)
);

CKINVDCx16_ASAP7_75t_R g1353 ( 
.A(n_987),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1047),
.Y(n_1354)
);

CKINVDCx20_ASAP7_75t_R g1355 ( 
.A(n_955),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_876),
.Y(n_1356)
);

INVxp33_ASAP7_75t_L g1357 ( 
.A(n_1200),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1067),
.Y(n_1358)
);

CKINVDCx20_ASAP7_75t_R g1359 ( 
.A(n_998),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1089),
.Y(n_1360)
);

CKINVDCx16_ASAP7_75t_R g1361 ( 
.A(n_1174),
.Y(n_1361)
);

INVxp33_ASAP7_75t_SL g1362 ( 
.A(n_880),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1131),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1239),
.Y(n_1364)
);

INVxp67_ASAP7_75t_SL g1365 ( 
.A(n_1046),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_878),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1246),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1279),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_867),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_871),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_884),
.Y(n_1371)
);

CKINVDCx20_ASAP7_75t_R g1372 ( 
.A(n_1018),
.Y(n_1372)
);

CKINVDCx20_ASAP7_75t_R g1373 ( 
.A(n_1037),
.Y(n_1373)
);

INVxp67_ASAP7_75t_L g1374 ( 
.A(n_974),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_887),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1051),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_897),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_912),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_934),
.Y(n_1379)
);

INVxp67_ASAP7_75t_SL g1380 ( 
.A(n_1211),
.Y(n_1380)
);

CKINVDCx20_ASAP7_75t_R g1381 ( 
.A(n_1054),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_940),
.Y(n_1382)
);

INVxp67_ASAP7_75t_SL g1383 ( 
.A(n_890),
.Y(n_1383)
);

CKINVDCx16_ASAP7_75t_R g1384 ( 
.A(n_1265),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_941),
.Y(n_1385)
);

BUFx10_ASAP7_75t_L g1386 ( 
.A(n_881),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_957),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_923),
.Y(n_1388)
);

INVxp33_ASAP7_75t_SL g1389 ( 
.A(n_886),
.Y(n_1389)
);

CKINVDCx20_ASAP7_75t_R g1390 ( 
.A(n_1077),
.Y(n_1390)
);

INVxp33_ASAP7_75t_SL g1391 ( 
.A(n_889),
.Y(n_1391)
);

CKINVDCx20_ASAP7_75t_R g1392 ( 
.A(n_1084),
.Y(n_1392)
);

INVxp67_ASAP7_75t_SL g1393 ( 
.A(n_920),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_979),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_879),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_882),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_995),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_885),
.Y(n_1398)
);

CKINVDCx20_ASAP7_75t_R g1399 ( 
.A(n_1122),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1002),
.Y(n_1400)
);

INVxp67_ASAP7_75t_SL g1401 ( 
.A(n_945),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1012),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1013),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1036),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_894),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1353),
.Y(n_1406)
);

CKINVDCx20_ASAP7_75t_R g1407 ( 
.A(n_1345),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1334),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1336),
.Y(n_1409)
);

INVx4_ASAP7_75t_L g1410 ( 
.A(n_1339),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1340),
.Y(n_1411)
);

BUFx6f_ASAP7_75t_L g1412 ( 
.A(n_1340),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1348),
.B(n_1136),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1351),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_1356),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_SL g1416 ( 
.A(n_1352),
.B(n_1170),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1343),
.B(n_926),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1327),
.Y(n_1418)
);

AOI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1337),
.A2(n_1167),
.B1(n_1189),
.B2(n_1163),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1383),
.B(n_968),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1330),
.Y(n_1421)
);

INVx5_ASAP7_75t_L g1422 ( 
.A(n_1340),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_1333),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1349),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1366),
.B(n_872),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_1335),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1338),
.Y(n_1427)
);

CKINVDCx11_ASAP7_75t_R g1428 ( 
.A(n_1386),
.Y(n_1428)
);

INVx3_ASAP7_75t_L g1429 ( 
.A(n_1341),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_L g1430 ( 
.A(n_1347),
.Y(n_1430)
);

BUFx6f_ASAP7_75t_L g1431 ( 
.A(n_1369),
.Y(n_1431)
);

BUFx2_ASAP7_75t_L g1432 ( 
.A(n_1342),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1370),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1325),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_1395),
.Y(n_1435)
);

BUFx6f_ASAP7_75t_L g1436 ( 
.A(n_1371),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1375),
.Y(n_1437)
);

CKINVDCx20_ASAP7_75t_R g1438 ( 
.A(n_1355),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1326),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1396),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1377),
.Y(n_1441)
);

AND2x6_ASAP7_75t_L g1442 ( 
.A(n_1346),
.B(n_943),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1378),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1379),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1361),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1382),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1385),
.Y(n_1447)
);

CKINVDCx8_ASAP7_75t_R g1448 ( 
.A(n_1384),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1387),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_SL g1450 ( 
.A1(n_1359),
.A2(n_877),
.B1(n_975),
.B2(n_868),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1394),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1393),
.B(n_1125),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1397),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1400),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1402),
.Y(n_1455)
);

CKINVDCx20_ASAP7_75t_R g1456 ( 
.A(n_1372),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1401),
.A2(n_1227),
.B1(n_895),
.B2(n_901),
.Y(n_1457)
);

BUFx6f_ASAP7_75t_L g1458 ( 
.A(n_1403),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_1398),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1404),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1405),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1350),
.Y(n_1462)
);

AND2x4_ASAP7_75t_L g1463 ( 
.A(n_1388),
.B(n_1220),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1376),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1354),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_L g1466 ( 
.A(n_1358),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1360),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1329),
.Y(n_1468)
);

INVx3_ASAP7_75t_L g1469 ( 
.A(n_1363),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1364),
.Y(n_1470)
);

AND2x6_ASAP7_75t_L g1471 ( 
.A(n_1367),
.B(n_943),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1368),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1331),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1324),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1328),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1411),
.Y(n_1476)
);

INVx3_ASAP7_75t_L g1477 ( 
.A(n_1412),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_1454),
.Y(n_1478)
);

NAND3xp33_ASAP7_75t_L g1479 ( 
.A(n_1474),
.B(n_1473),
.C(n_1416),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_1414),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1427),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1464),
.Y(n_1482)
);

INVx4_ASAP7_75t_L g1483 ( 
.A(n_1415),
.Y(n_1483)
);

NAND3xp33_ASAP7_75t_L g1484 ( 
.A(n_1457),
.B(n_1365),
.C(n_1344),
.Y(n_1484)
);

AOI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1425),
.A2(n_891),
.B(n_869),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1443),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1446),
.Y(n_1487)
);

INVxp33_ASAP7_75t_L g1488 ( 
.A(n_1450),
.Y(n_1488)
);

INVx5_ASAP7_75t_L g1489 ( 
.A(n_1466),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1420),
.B(n_1357),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1447),
.Y(n_1491)
);

INVx3_ASAP7_75t_L g1492 ( 
.A(n_1431),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1418),
.Y(n_1493)
);

INVx3_ASAP7_75t_L g1494 ( 
.A(n_1436),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1449),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1413),
.B(n_1362),
.Y(n_1496)
);

NAND2xp33_ASAP7_75t_L g1497 ( 
.A(n_1442),
.B(n_924),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1451),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1424),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1421),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1437),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1444),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1426),
.Y(n_1503)
);

AND3x2_ASAP7_75t_L g1504 ( 
.A(n_1406),
.B(n_978),
.C(n_944),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_L g1505 ( 
.A(n_1410),
.B(n_1389),
.Y(n_1505)
);

BUFx10_ASAP7_75t_L g1506 ( 
.A(n_1468),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1452),
.B(n_1391),
.Y(n_1507)
);

AND2x6_ASAP7_75t_L g1508 ( 
.A(n_1417),
.B(n_1462),
.Y(n_1508)
);

NAND3xp33_ASAP7_75t_L g1509 ( 
.A(n_1475),
.B(n_1380),
.C(n_1374),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1471),
.B(n_1442),
.Y(n_1510)
);

BUFx3_ASAP7_75t_L g1511 ( 
.A(n_1432),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1471),
.B(n_875),
.Y(n_1512)
);

INVx3_ASAP7_75t_L g1513 ( 
.A(n_1458),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1460),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_SL g1515 ( 
.A(n_1435),
.B(n_1332),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1466),
.Y(n_1516)
);

OAI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1419),
.A2(n_915),
.B1(n_1014),
.B2(n_908),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1440),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_R g1519 ( 
.A(n_1459),
.B(n_1373),
.Y(n_1519)
);

BUFx2_ASAP7_75t_L g1520 ( 
.A(n_1445),
.Y(n_1520)
);

XNOR2xp5_ASAP7_75t_L g1521 ( 
.A(n_1407),
.B(n_1381),
.Y(n_1521)
);

NAND3xp33_ASAP7_75t_L g1522 ( 
.A(n_1434),
.B(n_903),
.C(n_893),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1430),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_SL g1524 ( 
.A(n_1461),
.B(n_1386),
.Y(n_1524)
);

INVxp67_ASAP7_75t_SL g1525 ( 
.A(n_1454),
.Y(n_1525)
);

INVx2_ASAP7_75t_SL g1526 ( 
.A(n_1463),
.Y(n_1526)
);

INVx2_ASAP7_75t_SL g1527 ( 
.A(n_1469),
.Y(n_1527)
);

NAND3xp33_ASAP7_75t_SL g1528 ( 
.A(n_1448),
.B(n_1021),
.C(n_989),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1433),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1465),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1441),
.Y(n_1531)
);

BUFx6f_ASAP7_75t_SL g1532 ( 
.A(n_1439),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1467),
.Y(n_1533)
);

OR2x6_ASAP7_75t_L g1534 ( 
.A(n_1470),
.B(n_1107),
.Y(n_1534)
);

INVx4_ASAP7_75t_L g1535 ( 
.A(n_1422),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1472),
.Y(n_1536)
);

BUFx10_ASAP7_75t_L g1537 ( 
.A(n_1428),
.Y(n_1537)
);

BUFx6f_ASAP7_75t_L g1538 ( 
.A(n_1422),
.Y(n_1538)
);

INVxp67_ASAP7_75t_SL g1539 ( 
.A(n_1453),
.Y(n_1539)
);

BUFx6f_ASAP7_75t_L g1540 ( 
.A(n_1455),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1423),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1429),
.B(n_1390),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1408),
.B(n_939),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1409),
.B(n_1392),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1438),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1456),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1413),
.B(n_950),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1425),
.B(n_1399),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1411),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1411),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_SL g1551 ( 
.A(n_1416),
.B(n_923),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1443),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1412),
.Y(n_1553)
);

AOI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1464),
.A2(n_906),
.B(n_904),
.Y(n_1554)
);

OAI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1416),
.A2(n_1083),
.B1(n_1124),
.B2(n_1071),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1486),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1520),
.Y(n_1557)
);

BUFx3_ASAP7_75t_L g1558 ( 
.A(n_1514),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1507),
.B(n_1194),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1490),
.B(n_974),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_L g1561 ( 
.A(n_1478),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1487),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1496),
.B(n_1204),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1547),
.B(n_973),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1491),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1482),
.B(n_1006),
.Y(n_1566)
);

OA22x2_ASAP7_75t_L g1567 ( 
.A1(n_1551),
.A2(n_963),
.B1(n_1299),
.B2(n_954),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1511),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1529),
.Y(n_1569)
);

BUFx6f_ASAP7_75t_L g1570 ( 
.A(n_1478),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1495),
.B(n_1320),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1498),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1552),
.B(n_910),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1531),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_SL g1575 ( 
.A1(n_1548),
.A2(n_1123),
.B1(n_1147),
.B2(n_1052),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1499),
.B(n_1048),
.Y(n_1576)
);

BUFx6f_ASAP7_75t_L g1577 ( 
.A(n_1540),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1481),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1530),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1480),
.Y(n_1580)
);

NAND2x1p5_ASAP7_75t_L g1581 ( 
.A(n_1489),
.B(n_914),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1533),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1542),
.B(n_1196),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1536),
.Y(n_1584)
);

BUFx2_ASAP7_75t_L g1585 ( 
.A(n_1519),
.Y(n_1585)
);

NAND3xp33_ASAP7_75t_L g1586 ( 
.A(n_1484),
.B(n_952),
.C(n_942),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1493),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1500),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1492),
.B(n_1072),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1476),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1549),
.Y(n_1591)
);

NAND2x1p5_ASAP7_75t_L g1592 ( 
.A(n_1489),
.B(n_929),
.Y(n_1592)
);

CKINVDCx8_ASAP7_75t_R g1593 ( 
.A(n_1518),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1494),
.B(n_1073),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1550),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1539),
.B(n_911),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1513),
.B(n_1106),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1534),
.B(n_1196),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1526),
.B(n_1121),
.Y(n_1599)
);

INVxp33_ASAP7_75t_L g1600 ( 
.A(n_1521),
.Y(n_1600)
);

AO22x2_ASAP7_75t_L g1601 ( 
.A1(n_1528),
.A2(n_1137),
.B1(n_1318),
.B2(n_1127),
.Y(n_1601)
);

INVx6_ASAP7_75t_L g1602 ( 
.A(n_1537),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1503),
.B(n_1139),
.Y(n_1603)
);

BUFx6f_ASAP7_75t_L g1604 ( 
.A(n_1540),
.Y(n_1604)
);

BUFx2_ASAP7_75t_L g1605 ( 
.A(n_1534),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1505),
.B(n_916),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1541),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1516),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1523),
.B(n_1143),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1544),
.B(n_1233),
.Y(n_1610)
);

OA22x2_ASAP7_75t_L g1611 ( 
.A1(n_1504),
.A2(n_960),
.B1(n_971),
.B2(n_967),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1525),
.B(n_917),
.Y(n_1612)
);

INVxp67_ASAP7_75t_L g1613 ( 
.A(n_1509),
.Y(n_1613)
);

INVx4_ASAP7_75t_L g1614 ( 
.A(n_1538),
.Y(n_1614)
);

INVx3_ASAP7_75t_L g1615 ( 
.A(n_1477),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1554),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1501),
.Y(n_1617)
);

INVx5_ASAP7_75t_L g1618 ( 
.A(n_1538),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1502),
.Y(n_1619)
);

INVx1_ASAP7_75t_SL g1620 ( 
.A(n_1545),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1527),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1553),
.B(n_1155),
.Y(n_1622)
);

AND3x4_ASAP7_75t_L g1623 ( 
.A(n_1488),
.B(n_966),
.C(n_938),
.Y(n_1623)
);

AND3x1_ASAP7_75t_L g1624 ( 
.A(n_1546),
.B(n_1180),
.C(n_1178),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1543),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1485),
.Y(n_1626)
);

AND2x6_ASAP7_75t_L g1627 ( 
.A(n_1510),
.B(n_1184),
.Y(n_1627)
);

INVx1_ASAP7_75t_SL g1628 ( 
.A(n_1506),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1483),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1479),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1522),
.Y(n_1631)
);

NOR2xp33_ASAP7_75t_L g1632 ( 
.A(n_1517),
.B(n_1515),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1535),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1512),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1508),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1508),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1508),
.B(n_918),
.Y(n_1637)
);

NOR3xp33_ASAP7_75t_L g1638 ( 
.A(n_1555),
.B(n_1053),
.C(n_969),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1524),
.B(n_1185),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1532),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_SL g1641 ( 
.A(n_1497),
.B(n_1256),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1482),
.Y(n_1642)
);

BUFx6f_ASAP7_75t_L g1643 ( 
.A(n_1478),
.Y(n_1643)
);

XOR2x2_ASAP7_75t_L g1644 ( 
.A(n_1551),
.B(n_1),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1482),
.Y(n_1645)
);

AO22x2_ASAP7_75t_L g1646 ( 
.A1(n_1551),
.A2(n_1319),
.B1(n_1283),
.B2(n_1209),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_SL g1647 ( 
.A1(n_1488),
.A2(n_1282),
.B1(n_1023),
.B2(n_1245),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1486),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1490),
.B(n_1228),
.Y(n_1649)
);

INVx6_ASAP7_75t_L g1650 ( 
.A(n_1537),
.Y(n_1650)
);

BUFx3_ASAP7_75t_L g1651 ( 
.A(n_1514),
.Y(n_1651)
);

BUFx2_ASAP7_75t_L g1652 ( 
.A(n_1520),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1490),
.B(n_1228),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1514),
.B(n_1193),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1507),
.B(n_1292),
.Y(n_1655)
);

INVx3_ASAP7_75t_L g1656 ( 
.A(n_1478),
.Y(n_1656)
);

NAND2x1p5_ASAP7_75t_L g1657 ( 
.A(n_1499),
.B(n_1160),
.Y(n_1657)
);

BUFx3_ASAP7_75t_L g1658 ( 
.A(n_1514),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1486),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1547),
.B(n_922),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_SL g1661 ( 
.A(n_1507),
.B(n_1161),
.Y(n_1661)
);

BUFx6f_ASAP7_75t_L g1662 ( 
.A(n_1478),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1486),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1514),
.B(n_1247),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1547),
.B(n_928),
.Y(n_1665)
);

AND2x4_ASAP7_75t_L g1666 ( 
.A(n_1514),
.B(n_1255),
.Y(n_1666)
);

BUFx2_ASAP7_75t_L g1667 ( 
.A(n_1520),
.Y(n_1667)
);

CKINVDCx16_ASAP7_75t_R g1668 ( 
.A(n_1519),
.Y(n_1668)
);

AOI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1486),
.A2(n_892),
.B1(n_936),
.B2(n_888),
.Y(n_1669)
);

INVx1_ASAP7_75t_SL g1670 ( 
.A(n_1490),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1486),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_SL g1672 ( 
.A(n_1507),
.B(n_1165),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1486),
.Y(n_1673)
);

BUFx6f_ASAP7_75t_L g1674 ( 
.A(n_1478),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_1480),
.Y(n_1675)
);

AOI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1507),
.A2(n_1208),
.B1(n_1238),
.B2(n_1186),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1486),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1482),
.Y(n_1678)
);

INVx1_ASAP7_75t_SL g1679 ( 
.A(n_1490),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1486),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1486),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1486),
.Y(n_1682)
);

AO22x2_ASAP7_75t_L g1683 ( 
.A1(n_1551),
.A2(n_1308),
.B1(n_1270),
.B2(n_1261),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1547),
.B(n_948),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1507),
.B(n_972),
.Y(n_1685)
);

NAND3xp33_ASAP7_75t_L g1686 ( 
.A(n_1484),
.B(n_981),
.C(n_977),
.Y(n_1686)
);

BUFx6f_ASAP7_75t_L g1687 ( 
.A(n_1478),
.Y(n_1687)
);

NAND2x1p5_ASAP7_75t_L g1688 ( 
.A(n_1499),
.B(n_951),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1547),
.B(n_953),
.Y(n_1689)
);

AO22x2_ASAP7_75t_L g1690 ( 
.A1(n_1551),
.A2(n_1231),
.B1(n_1257),
.B2(n_1192),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_1480),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1514),
.B(n_1011),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1482),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1486),
.Y(n_1694)
);

BUFx3_ASAP7_75t_L g1695 ( 
.A(n_1514),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1482),
.Y(n_1696)
);

AO22x2_ASAP7_75t_L g1697 ( 
.A1(n_1551),
.A2(n_1120),
.B1(n_965),
.B2(n_993),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1490),
.B(n_1258),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1490),
.B(n_1258),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1490),
.B(n_1323),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1514),
.B(n_956),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1482),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1670),
.B(n_1323),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1610),
.A2(n_1027),
.B1(n_1034),
.B2(n_1022),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1563),
.B(n_1195),
.Y(n_1705)
);

INVx2_ASAP7_75t_SL g1706 ( 
.A(n_1652),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1556),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1625),
.B(n_1049),
.Y(n_1708)
);

AOI21xp5_ASAP7_75t_L g1709 ( 
.A1(n_1634),
.A2(n_1005),
.B(n_976),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1630),
.B(n_1058),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1685),
.B(n_1070),
.Y(n_1711)
);

INVx3_ASAP7_75t_L g1712 ( 
.A(n_1561),
.Y(n_1712)
);

INVxp67_ASAP7_75t_L g1713 ( 
.A(n_1560),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1606),
.B(n_1092),
.Y(n_1714)
);

INVx5_ASAP7_75t_L g1715 ( 
.A(n_1602),
.Y(n_1715)
);

BUFx4f_ASAP7_75t_SL g1716 ( 
.A(n_1628),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1562),
.Y(n_1717)
);

INVx3_ASAP7_75t_L g1718 ( 
.A(n_1561),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_SL g1719 ( 
.A(n_1632),
.B(n_896),
.Y(n_1719)
);

INVx2_ASAP7_75t_SL g1720 ( 
.A(n_1667),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1565),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_SL g1722 ( 
.A(n_1679),
.B(n_898),
.Y(n_1722)
);

OR2x6_ASAP7_75t_L g1723 ( 
.A(n_1568),
.B(n_1094),
.Y(n_1723)
);

INVx2_ASAP7_75t_SL g1724 ( 
.A(n_1557),
.Y(n_1724)
);

OR2x2_ASAP7_75t_SL g1725 ( 
.A(n_1668),
.B(n_1113),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1642),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1559),
.B(n_1100),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_1580),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_SL g1729 ( 
.A(n_1655),
.B(n_899),
.Y(n_1729)
);

INVx3_ASAP7_75t_L g1730 ( 
.A(n_1570),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1649),
.B(n_992),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1572),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1648),
.Y(n_1733)
);

OAI22xp5_ASAP7_75t_L g1734 ( 
.A1(n_1635),
.A2(n_1134),
.B1(n_1187),
.B2(n_1133),
.Y(n_1734)
);

NOR3xp33_ASAP7_75t_SL g1735 ( 
.A(n_1647),
.B(n_1001),
.C(n_996),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1645),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1678),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1693),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1638),
.A2(n_1217),
.B1(n_1300),
.B2(n_1206),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1659),
.Y(n_1740)
);

INVx2_ASAP7_75t_SL g1741 ( 
.A(n_1570),
.Y(n_1741)
);

OR2x6_ASAP7_75t_L g1742 ( 
.A(n_1650),
.B(n_1109),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1663),
.B(n_1114),
.Y(n_1743)
);

NAND3xp33_ASAP7_75t_SL g1744 ( 
.A(n_1575),
.B(n_1004),
.C(n_1003),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1671),
.Y(n_1745)
);

OAI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1626),
.A2(n_1129),
.B(n_1128),
.Y(n_1746)
);

BUFx3_ASAP7_75t_L g1747 ( 
.A(n_1643),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1673),
.Y(n_1748)
);

INVx4_ASAP7_75t_L g1749 ( 
.A(n_1618),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1677),
.B(n_1135),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1696),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1680),
.B(n_1141),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1681),
.B(n_1146),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1631),
.A2(n_1149),
.B1(n_1153),
.B2(n_1151),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_L g1755 ( 
.A(n_1620),
.B(n_1010),
.Y(n_1755)
);

AOI22xp33_ASAP7_75t_L g1756 ( 
.A1(n_1623),
.A2(n_1154),
.B1(n_1171),
.B2(n_1156),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1682),
.Y(n_1757)
);

INVx2_ASAP7_75t_SL g1758 ( 
.A(n_1643),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1694),
.B(n_1176),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1660),
.B(n_1665),
.Y(n_1760)
);

OAI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1616),
.A2(n_1197),
.B(n_1190),
.Y(n_1761)
);

AND2x6_ASAP7_75t_L g1762 ( 
.A(n_1636),
.B(n_1207),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_L g1763 ( 
.A(n_1583),
.B(n_1016),
.Y(n_1763)
);

BUFx3_ASAP7_75t_L g1764 ( 
.A(n_1662),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1653),
.B(n_1017),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1579),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1702),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1684),
.B(n_1218),
.Y(n_1768)
);

INVx1_ASAP7_75t_SL g1769 ( 
.A(n_1698),
.Y(n_1769)
);

AOI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1637),
.A2(n_1242),
.B(n_1230),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1582),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1584),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_SL g1773 ( 
.A(n_1629),
.B(n_902),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1689),
.B(n_1244),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1564),
.B(n_1699),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1574),
.Y(n_1776)
);

NAND2x1_ASAP7_75t_L g1777 ( 
.A(n_1577),
.B(n_1252),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1700),
.B(n_1260),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1627),
.A2(n_1274),
.B1(n_1293),
.B2(n_1286),
.Y(n_1779)
);

INVx5_ASAP7_75t_L g1780 ( 
.A(n_1627),
.Y(n_1780)
);

INVx2_ASAP7_75t_SL g1781 ( 
.A(n_1662),
.Y(n_1781)
);

AND2x4_ASAP7_75t_L g1782 ( 
.A(n_1558),
.B(n_1309),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1569),
.B(n_1312),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1578),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_SL g1785 ( 
.A(n_1577),
.B(n_905),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_1604),
.B(n_907),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_L g1787 ( 
.A(n_1613),
.B(n_1025),
.Y(n_1787)
);

BUFx3_ASAP7_75t_L g1788 ( 
.A(n_1674),
.Y(n_1788)
);

BUFx2_ASAP7_75t_L g1789 ( 
.A(n_1605),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1590),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1587),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1591),
.Y(n_1792)
);

OR2x6_ASAP7_75t_L g1793 ( 
.A(n_1585),
.B(n_1316),
.Y(n_1793)
);

BUFx6f_ASAP7_75t_L g1794 ( 
.A(n_1674),
.Y(n_1794)
);

BUFx12f_ASAP7_75t_L g1795 ( 
.A(n_1675),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1588),
.Y(n_1796)
);

O2A1O1Ixp5_ASAP7_75t_L g1797 ( 
.A1(n_1596),
.A2(n_1051),
.B(n_1102),
.C(n_931),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1595),
.Y(n_1798)
);

NOR2x1p5_ASAP7_75t_L g1799 ( 
.A(n_1691),
.B(n_1029),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1607),
.Y(n_1800)
);

AOI21x1_ASAP7_75t_L g1801 ( 
.A1(n_1571),
.A2(n_1051),
.B(n_919),
.Y(n_1801)
);

BUFx6f_ASAP7_75t_L g1802 ( 
.A(n_1687),
.Y(n_1802)
);

BUFx2_ASAP7_75t_L g1803 ( 
.A(n_1687),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1608),
.Y(n_1804)
);

AOI22xp33_ASAP7_75t_L g1805 ( 
.A1(n_1586),
.A2(n_1051),
.B1(n_924),
.B2(n_900),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1603),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1609),
.Y(n_1807)
);

INVx2_ASAP7_75t_SL g1808 ( 
.A(n_1692),
.Y(n_1808)
);

BUFx6f_ASAP7_75t_L g1809 ( 
.A(n_1604),
.Y(n_1809)
);

BUFx10_ASAP7_75t_L g1810 ( 
.A(n_1639),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_SL g1811 ( 
.A(n_1676),
.B(n_909),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1621),
.Y(n_1812)
);

BUFx2_ASAP7_75t_L g1813 ( 
.A(n_1601),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1617),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1619),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1599),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1573),
.Y(n_1817)
);

CKINVDCx20_ASAP7_75t_R g1818 ( 
.A(n_1593),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1566),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_SL g1820 ( 
.A(n_1686),
.B(n_921),
.Y(n_1820)
);

INVx1_ASAP7_75t_SL g1821 ( 
.A(n_1651),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1657),
.B(n_1040),
.Y(n_1822)
);

XOR2x2_ASAP7_75t_L g1823 ( 
.A(n_1644),
.B(n_1),
.Y(n_1823)
);

NOR3xp33_ASAP7_75t_SL g1824 ( 
.A(n_1661),
.B(n_1055),
.C(n_1043),
.Y(n_1824)
);

INVx1_ASAP7_75t_SL g1825 ( 
.A(n_1658),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1622),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1612),
.B(n_925),
.Y(n_1827)
);

BUFx3_ASAP7_75t_L g1828 ( 
.A(n_1695),
.Y(n_1828)
);

OR2x2_ASAP7_75t_SL g1829 ( 
.A(n_1640),
.B(n_900),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1589),
.Y(n_1830)
);

INVx2_ASAP7_75t_SL g1831 ( 
.A(n_1576),
.Y(n_1831)
);

NAND2x1_ASAP7_75t_L g1832 ( 
.A(n_1656),
.B(n_924),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_SL g1833 ( 
.A(n_1672),
.B(n_927),
.Y(n_1833)
);

INVx1_ASAP7_75t_SL g1834 ( 
.A(n_1598),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1594),
.Y(n_1835)
);

INVx2_ASAP7_75t_SL g1836 ( 
.A(n_1654),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1597),
.Y(n_1837)
);

BUFx3_ASAP7_75t_L g1838 ( 
.A(n_1618),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1615),
.Y(n_1839)
);

BUFx2_ASAP7_75t_L g1840 ( 
.A(n_1646),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1664),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1666),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1669),
.B(n_1690),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1633),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1581),
.B(n_1057),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1701),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1567),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1600),
.B(n_1060),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1683),
.Y(n_1849)
);

AOI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1641),
.A2(n_1099),
.B(n_1064),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1697),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1624),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1611),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1688),
.Y(n_1854)
);

NOR2xp67_ASAP7_75t_L g1855 ( 
.A(n_1614),
.B(n_930),
.Y(n_1855)
);

CKINVDCx5p33_ASAP7_75t_R g1856 ( 
.A(n_1592),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_SL g1857 ( 
.A(n_1606),
.B(n_932),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1642),
.Y(n_1858)
);

OR2x6_ASAP7_75t_L g1859 ( 
.A(n_1652),
.B(n_1064),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1556),
.Y(n_1860)
);

BUFx2_ASAP7_75t_L g1861 ( 
.A(n_1652),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1625),
.B(n_935),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1625),
.B(n_937),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1642),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1625),
.B(n_946),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1625),
.B(n_947),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1638),
.A2(n_1051),
.B1(n_1099),
.B2(n_1064),
.Y(n_1867)
);

INVx3_ASAP7_75t_L g1868 ( 
.A(n_1561),
.Y(n_1868)
);

BUFx6f_ASAP7_75t_L g1869 ( 
.A(n_1561),
.Y(n_1869)
);

BUFx6f_ASAP7_75t_L g1870 ( 
.A(n_1561),
.Y(n_1870)
);

AND2x4_ASAP7_75t_L g1871 ( 
.A(n_1558),
.B(n_1063),
.Y(n_1871)
);

NOR3xp33_ASAP7_75t_SL g1872 ( 
.A(n_1647),
.B(n_1075),
.C(n_1069),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1642),
.Y(n_1873)
);

AOI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1610),
.A2(n_958),
.B1(n_961),
.B2(n_959),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_L g1875 ( 
.A(n_1610),
.B(n_1079),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1556),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1625),
.B(n_962),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_SL g1878 ( 
.A(n_1606),
.B(n_964),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1556),
.Y(n_1879)
);

CKINVDCx5p33_ASAP7_75t_R g1880 ( 
.A(n_1580),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1556),
.Y(n_1881)
);

INVx2_ASAP7_75t_SL g1882 ( 
.A(n_1652),
.Y(n_1882)
);

AOI21xp5_ASAP7_75t_L g1883 ( 
.A1(n_1625),
.A2(n_1112),
.B(n_1099),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1625),
.B(n_970),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_SL g1885 ( 
.A(n_1606),
.B(n_982),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_SL g1886 ( 
.A(n_1606),
.B(n_983),
.Y(n_1886)
);

INVx2_ASAP7_75t_SL g1887 ( 
.A(n_1652),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_SL g1888 ( 
.A(n_1606),
.B(n_984),
.Y(n_1888)
);

BUFx3_ASAP7_75t_L g1889 ( 
.A(n_1561),
.Y(n_1889)
);

AND2x6_ASAP7_75t_L g1890 ( 
.A(n_1635),
.B(n_1112),
.Y(n_1890)
);

NOR3xp33_ASAP7_75t_SL g1891 ( 
.A(n_1647),
.B(n_1082),
.C(n_1080),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1556),
.Y(n_1892)
);

INVx4_ASAP7_75t_L g1893 ( 
.A(n_1618),
.Y(n_1893)
);

INVx4_ASAP7_75t_L g1894 ( 
.A(n_1618),
.Y(n_1894)
);

AOI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1610),
.A2(n_985),
.B1(n_990),
.B2(n_986),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_1610),
.B(n_1085),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1642),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_SL g1898 ( 
.A(n_1606),
.B(n_991),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1625),
.B(n_994),
.Y(n_1899)
);

BUFx4f_ASAP7_75t_L g1900 ( 
.A(n_1602),
.Y(n_1900)
);

INVxp67_ASAP7_75t_L g1901 ( 
.A(n_1560),
.Y(n_1901)
);

INVx2_ASAP7_75t_SL g1902 ( 
.A(n_1652),
.Y(n_1902)
);

CKINVDCx5p33_ASAP7_75t_R g1903 ( 
.A(n_1580),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1625),
.B(n_997),
.Y(n_1904)
);

O2A1O1Ixp33_ASAP7_75t_L g1905 ( 
.A1(n_1705),
.A2(n_1102),
.B(n_931),
.C(n_1101),
.Y(n_1905)
);

BUFx6f_ASAP7_75t_L g1906 ( 
.A(n_1794),
.Y(n_1906)
);

AOI221xp5_ASAP7_75t_L g1907 ( 
.A1(n_1744),
.A2(n_1104),
.B1(n_1105),
.B2(n_1103),
.C(n_1096),
.Y(n_1907)
);

HB1xp67_ASAP7_75t_L g1908 ( 
.A(n_1861),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_SL g1909 ( 
.A(n_1769),
.B(n_999),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1760),
.B(n_1000),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1726),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_SL g1912 ( 
.A(n_1728),
.B(n_1007),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1875),
.B(n_1008),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1896),
.B(n_1009),
.Y(n_1914)
);

BUFx3_ASAP7_75t_L g1915 ( 
.A(n_1715),
.Y(n_1915)
);

NAND2x1p5_ASAP7_75t_L g1916 ( 
.A(n_1715),
.B(n_1112),
.Y(n_1916)
);

OAI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1711),
.A2(n_1019),
.B1(n_1020),
.B2(n_1015),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_SL g1918 ( 
.A(n_1775),
.B(n_1713),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1707),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_SL g1920 ( 
.A(n_1901),
.B(n_1817),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1727),
.B(n_1026),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1717),
.Y(n_1922)
);

BUFx2_ASAP7_75t_L g1923 ( 
.A(n_1706),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1736),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1721),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1732),
.Y(n_1926)
);

INVx4_ASAP7_75t_L g1927 ( 
.A(n_1900),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1733),
.Y(n_1928)
);

NOR2xp67_ASAP7_75t_L g1929 ( 
.A(n_1880),
.B(n_1028),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1740),
.Y(n_1930)
);

OR2x2_ASAP7_75t_L g1931 ( 
.A(n_1720),
.B(n_1882),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1737),
.Y(n_1932)
);

BUFx6f_ASAP7_75t_L g1933 ( 
.A(n_1794),
.Y(n_1933)
);

BUFx2_ASAP7_75t_L g1934 ( 
.A(n_1887),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1763),
.B(n_1030),
.Y(n_1935)
);

BUFx2_ASAP7_75t_L g1936 ( 
.A(n_1902),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1819),
.B(n_1031),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1745),
.B(n_1032),
.Y(n_1938)
);

AND3x1_ASAP7_75t_SL g1939 ( 
.A(n_1852),
.B(n_1111),
.C(n_1108),
.Y(n_1939)
);

AOI21xp5_ASAP7_75t_L g1940 ( 
.A1(n_1761),
.A2(n_1243),
.B(n_1237),
.Y(n_1940)
);

OAI22xp5_ASAP7_75t_L g1941 ( 
.A1(n_1746),
.A2(n_1038),
.B1(n_1039),
.B2(n_1035),
.Y(n_1941)
);

AOI22xp33_ASAP7_75t_SL g1942 ( 
.A1(n_1787),
.A2(n_1322),
.B1(n_1317),
.B2(n_1157),
.Y(n_1942)
);

INVx3_ASAP7_75t_L g1943 ( 
.A(n_1749),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1724),
.B(n_1144),
.Y(n_1944)
);

BUFx3_ASAP7_75t_L g1945 ( 
.A(n_1747),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1738),
.Y(n_1946)
);

INVx5_ASAP7_75t_L g1947 ( 
.A(n_1795),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1748),
.Y(n_1948)
);

BUFx2_ASAP7_75t_SL g1949 ( 
.A(n_1818),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1731),
.B(n_1158),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1757),
.B(n_1041),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1860),
.B(n_1042),
.Y(n_1952)
);

NAND2x1p5_ASAP7_75t_L g1953 ( 
.A(n_1821),
.B(n_1237),
.Y(n_1953)
);

BUFx6f_ASAP7_75t_L g1954 ( 
.A(n_1802),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1876),
.Y(n_1955)
);

AND3x1_ASAP7_75t_SL g1956 ( 
.A(n_1823),
.B(n_1168),
.C(n_1159),
.Y(n_1956)
);

AND2x6_ASAP7_75t_L g1957 ( 
.A(n_1849),
.B(n_1237),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1879),
.B(n_1044),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1765),
.B(n_1169),
.Y(n_1959)
);

INVx3_ASAP7_75t_L g1960 ( 
.A(n_1893),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1703),
.B(n_1181),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1881),
.B(n_1045),
.Y(n_1962)
);

INVx5_ASAP7_75t_L g1963 ( 
.A(n_1802),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1892),
.Y(n_1964)
);

AOI22xp33_ASAP7_75t_L g1965 ( 
.A1(n_1719),
.A2(n_1243),
.B1(n_1056),
.B2(n_1059),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1766),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1755),
.B(n_1183),
.Y(n_1967)
);

INVx3_ASAP7_75t_L g1968 ( 
.A(n_1894),
.Y(n_1968)
);

INVx3_ASAP7_75t_L g1969 ( 
.A(n_1828),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1710),
.B(n_1050),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1708),
.B(n_1061),
.Y(n_1971)
);

BUFx3_ASAP7_75t_L g1972 ( 
.A(n_1764),
.Y(n_1972)
);

HB1xp67_ASAP7_75t_L g1973 ( 
.A(n_1789),
.Y(n_1973)
);

BUFx6f_ASAP7_75t_L g1974 ( 
.A(n_1869),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1751),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1771),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1772),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1816),
.B(n_1203),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1815),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1862),
.B(n_1062),
.Y(n_1980)
);

INVx5_ASAP7_75t_L g1981 ( 
.A(n_1869),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1776),
.Y(n_1982)
);

CKINVDCx5p33_ASAP7_75t_R g1983 ( 
.A(n_1903),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1863),
.B(n_1065),
.Y(n_1984)
);

NAND2xp33_ASAP7_75t_L g1985 ( 
.A(n_1704),
.B(n_1762),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1870),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1865),
.B(n_1066),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1866),
.B(n_1068),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1791),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1822),
.B(n_1205),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1877),
.B(n_1076),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1767),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_SL g1993 ( 
.A(n_1884),
.B(n_1081),
.Y(n_1993)
);

NOR2xp33_ASAP7_75t_L g1994 ( 
.A(n_1848),
.B(n_1210),
.Y(n_1994)
);

AND2x6_ASAP7_75t_L g1995 ( 
.A(n_1809),
.B(n_1870),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1796),
.Y(n_1996)
);

INVxp67_ASAP7_75t_L g1997 ( 
.A(n_1803),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1899),
.B(n_1086),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1800),
.Y(n_1999)
);

BUFx4f_ASAP7_75t_L g2000 ( 
.A(n_1809),
.Y(n_2000)
);

AOI21xp33_ASAP7_75t_L g2001 ( 
.A1(n_1904),
.A2(n_1729),
.B(n_1778),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1804),
.Y(n_2002)
);

NOR2xp33_ASAP7_75t_L g2003 ( 
.A(n_1834),
.B(n_1215),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1714),
.B(n_1087),
.Y(n_2004)
);

CKINVDCx11_ASAP7_75t_R g2005 ( 
.A(n_1742),
.Y(n_2005)
);

NOR2xp33_ASAP7_75t_L g2006 ( 
.A(n_1825),
.B(n_1216),
.Y(n_2006)
);

BUFx6f_ASAP7_75t_L g2007 ( 
.A(n_1838),
.Y(n_2007)
);

BUFx2_ASAP7_75t_L g2008 ( 
.A(n_1788),
.Y(n_2008)
);

NOR2xp33_ASAP7_75t_L g2009 ( 
.A(n_1840),
.B(n_1219),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1792),
.B(n_1088),
.Y(n_2010)
);

HB1xp67_ASAP7_75t_L g2011 ( 
.A(n_1889),
.Y(n_2011)
);

BUFx6f_ASAP7_75t_L g2012 ( 
.A(n_1741),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1814),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1798),
.B(n_1091),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_SL g2015 ( 
.A(n_1844),
.B(n_1093),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1784),
.Y(n_2016)
);

BUFx6f_ASAP7_75t_L g2017 ( 
.A(n_1758),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1790),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1858),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1864),
.Y(n_2020)
);

BUFx3_ASAP7_75t_L g2021 ( 
.A(n_1716),
.Y(n_2021)
);

OR2x6_ASAP7_75t_L g2022 ( 
.A(n_1831),
.B(n_1243),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1873),
.Y(n_2023)
);

AOI22xp5_ASAP7_75t_L g2024 ( 
.A1(n_1853),
.A2(n_1097),
.B1(n_1098),
.B2(n_1095),
.Y(n_2024)
);

BUFx6f_ASAP7_75t_L g2025 ( 
.A(n_1781),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1897),
.B(n_1110),
.Y(n_2026)
);

BUFx3_ASAP7_75t_L g2027 ( 
.A(n_1712),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1827),
.B(n_1115),
.Y(n_2028)
);

NOR2xp33_ASAP7_75t_L g2029 ( 
.A(n_1813),
.B(n_1224),
.Y(n_2029)
);

BUFx2_ASAP7_75t_L g2030 ( 
.A(n_1718),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1743),
.B(n_1116),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1845),
.B(n_1234),
.Y(n_2032)
);

OR2x2_ASAP7_75t_L g2033 ( 
.A(n_1808),
.B(n_1240),
.Y(n_2033)
);

CKINVDCx20_ASAP7_75t_R g2034 ( 
.A(n_1725),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1783),
.Y(n_2035)
);

INVxp67_ASAP7_75t_SL g2036 ( 
.A(n_1730),
.Y(n_2036)
);

AND2x4_ASAP7_75t_L g2037 ( 
.A(n_1836),
.B(n_456),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1812),
.Y(n_2038)
);

BUFx6f_ASAP7_75t_L g2039 ( 
.A(n_1868),
.Y(n_2039)
);

HB1xp67_ASAP7_75t_L g2040 ( 
.A(n_1851),
.Y(n_2040)
);

INVx3_ASAP7_75t_L g2041 ( 
.A(n_1810),
.Y(n_2041)
);

NOR2xp33_ASAP7_75t_L g2042 ( 
.A(n_1856),
.B(n_1722),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1750),
.Y(n_2043)
);

INVxp67_ASAP7_75t_SL g2044 ( 
.A(n_1841),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1752),
.Y(n_2045)
);

BUFx2_ASAP7_75t_L g2046 ( 
.A(n_1871),
.Y(n_2046)
);

OAI22xp5_ASAP7_75t_L g2047 ( 
.A1(n_1843),
.A2(n_1118),
.B1(n_1119),
.B2(n_1117),
.Y(n_2047)
);

INVx6_ASAP7_75t_L g2048 ( 
.A(n_1742),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_SL g2049 ( 
.A(n_1854),
.B(n_1126),
.Y(n_2049)
);

INVx6_ASAP7_75t_L g2050 ( 
.A(n_1780),
.Y(n_2050)
);

BUFx6f_ASAP7_75t_L g2051 ( 
.A(n_1846),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1799),
.B(n_1241),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1839),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_2043),
.B(n_1756),
.Y(n_2054)
);

AOI22xp33_ASAP7_75t_L g2055 ( 
.A1(n_1994),
.A2(n_1811),
.B1(n_1847),
.B2(n_1754),
.Y(n_2055)
);

BUFx3_ASAP7_75t_L g2056 ( 
.A(n_1915),
.Y(n_2056)
);

BUFx12f_ASAP7_75t_L g2057 ( 
.A(n_1927),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1919),
.Y(n_2058)
);

AOI21xp5_ASAP7_75t_L g2059 ( 
.A1(n_2001),
.A2(n_1850),
.B(n_1898),
.Y(n_2059)
);

BUFx2_ASAP7_75t_L g2060 ( 
.A(n_1908),
.Y(n_2060)
);

BUFx3_ASAP7_75t_L g2061 ( 
.A(n_2000),
.Y(n_2061)
);

INVxp67_ASAP7_75t_L g2062 ( 
.A(n_1973),
.Y(n_2062)
);

NOR2xp33_ASAP7_75t_L g2063 ( 
.A(n_1967),
.B(n_1773),
.Y(n_2063)
);

AOI22xp5_ASAP7_75t_L g2064 ( 
.A1(n_2042),
.A2(n_1895),
.B1(n_1874),
.B2(n_1842),
.Y(n_2064)
);

NOR2x1_ASAP7_75t_SL g2065 ( 
.A(n_2045),
.B(n_1801),
.Y(n_2065)
);

INVx3_ASAP7_75t_L g2066 ( 
.A(n_1945),
.Y(n_2066)
);

INVx4_ASAP7_75t_L g2067 ( 
.A(n_1963),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1922),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1910),
.B(n_1753),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1925),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1926),
.Y(n_2071)
);

BUFx8_ASAP7_75t_L g2072 ( 
.A(n_2008),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_2035),
.B(n_1759),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1928),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1930),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1948),
.Y(n_2076)
);

NOR2xp33_ASAP7_75t_L g2077 ( 
.A(n_1935),
.B(n_1793),
.Y(n_2077)
);

BUFx2_ASAP7_75t_L g2078 ( 
.A(n_1923),
.Y(n_2078)
);

BUFx2_ASAP7_75t_L g2079 ( 
.A(n_1934),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1955),
.Y(n_2080)
);

INVx4_ASAP7_75t_L g2081 ( 
.A(n_1963),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1913),
.B(n_1914),
.Y(n_2082)
);

INVx2_ASAP7_75t_L g2083 ( 
.A(n_1964),
.Y(n_2083)
);

OAI22xp33_ASAP7_75t_L g2084 ( 
.A1(n_1912),
.A2(n_1793),
.B1(n_1859),
.B2(n_1723),
.Y(n_2084)
);

OAI22xp5_ASAP7_75t_L g2085 ( 
.A1(n_1966),
.A2(n_1878),
.B1(n_1885),
.B2(n_1857),
.Y(n_2085)
);

INVx4_ASAP7_75t_L g2086 ( 
.A(n_1981),
.Y(n_2086)
);

INVx6_ASAP7_75t_L g2087 ( 
.A(n_1981),
.Y(n_2087)
);

AOI22xp5_ASAP7_75t_L g2088 ( 
.A1(n_2034),
.A2(n_1855),
.B1(n_1735),
.B2(n_1872),
.Y(n_2088)
);

OAI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_1976),
.A2(n_1886),
.B1(n_1888),
.B2(n_1739),
.Y(n_2089)
);

AOI22xp5_ASAP7_75t_L g2090 ( 
.A1(n_2006),
.A2(n_1891),
.B1(n_1833),
.B2(n_1835),
.Y(n_2090)
);

CKINVDCx5p33_ASAP7_75t_R g2091 ( 
.A(n_1983),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1977),
.Y(n_2092)
);

BUFx8_ASAP7_75t_L g2093 ( 
.A(n_1936),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1979),
.Y(n_2094)
);

BUFx2_ASAP7_75t_L g2095 ( 
.A(n_1995),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_SL g2096 ( 
.A(n_2051),
.B(n_1780),
.Y(n_2096)
);

BUFx6f_ASAP7_75t_L g2097 ( 
.A(n_1906),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1982),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1918),
.B(n_1768),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1989),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1937),
.B(n_1774),
.Y(n_2101)
);

INVx1_ASAP7_75t_SL g2102 ( 
.A(n_1931),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_SL g2103 ( 
.A(n_2051),
.B(n_1824),
.Y(n_2103)
);

AOI221xp5_ASAP7_75t_L g2104 ( 
.A1(n_2009),
.A2(n_1867),
.B1(n_1779),
.B2(n_1806),
.C(n_1807),
.Y(n_2104)
);

AND2x4_ASAP7_75t_L g2105 ( 
.A(n_1972),
.B(n_1969),
.Y(n_2105)
);

BUFx6f_ASAP7_75t_L g2106 ( 
.A(n_1906),
.Y(n_2106)
);

NOR2xp33_ASAP7_75t_L g2107 ( 
.A(n_1920),
.B(n_1723),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1996),
.Y(n_2108)
);

BUFx6f_ASAP7_75t_L g2109 ( 
.A(n_1933),
.Y(n_2109)
);

OAI22xp33_ASAP7_75t_L g2110 ( 
.A1(n_2044),
.A2(n_1859),
.B1(n_1826),
.B2(n_1830),
.Y(n_2110)
);

INVxp67_ASAP7_75t_SL g2111 ( 
.A(n_1997),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1999),
.Y(n_2112)
);

INVxp67_ASAP7_75t_SL g2113 ( 
.A(n_2011),
.Y(n_2113)
);

OR2x6_ASAP7_75t_SL g2114 ( 
.A(n_2047),
.B(n_1837),
.Y(n_2114)
);

AND2x4_ASAP7_75t_L g2115 ( 
.A(n_2027),
.B(n_1782),
.Y(n_2115)
);

HB1xp67_ASAP7_75t_L g2116 ( 
.A(n_1933),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_1921),
.B(n_2002),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2013),
.Y(n_2118)
);

AOI22xp33_ASAP7_75t_L g2119 ( 
.A1(n_1985),
.A2(n_1762),
.B1(n_1820),
.B2(n_1786),
.Y(n_2119)
);

INVx1_ASAP7_75t_SL g2120 ( 
.A(n_2021),
.Y(n_2120)
);

OAI22xp5_ASAP7_75t_L g2121 ( 
.A1(n_1980),
.A2(n_1829),
.B1(n_1777),
.B2(n_1805),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2018),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2019),
.Y(n_2123)
);

OAI22xp5_ASAP7_75t_SL g2124 ( 
.A1(n_1942),
.A2(n_1250),
.B1(n_1254),
.B2(n_1248),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2020),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2023),
.Y(n_2126)
);

BUFx12f_ASAP7_75t_L g2127 ( 
.A(n_2005),
.Y(n_2127)
);

AOI21xp5_ASAP7_75t_L g2128 ( 
.A1(n_1940),
.A2(n_1709),
.B(n_1785),
.Y(n_2128)
);

INVx1_ASAP7_75t_SL g2129 ( 
.A(n_1949),
.Y(n_2129)
);

OAI22xp5_ASAP7_75t_L g2130 ( 
.A1(n_1984),
.A2(n_1734),
.B1(n_1770),
.B2(n_1883),
.Y(n_2130)
);

AOI22xp33_ASAP7_75t_L g2131 ( 
.A1(n_1907),
.A2(n_1762),
.B1(n_1890),
.B2(n_1132),
.Y(n_2131)
);

NAND2xp33_ASAP7_75t_L g2132 ( 
.A(n_1995),
.B(n_1890),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_1970),
.B(n_1890),
.Y(n_2133)
);

NAND3xp33_ASAP7_75t_L g2134 ( 
.A(n_1905),
.B(n_1797),
.C(n_1263),
.Y(n_2134)
);

OAI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_1987),
.A2(n_1832),
.B1(n_1138),
.B2(n_1140),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1911),
.Y(n_2136)
);

HB1xp67_ASAP7_75t_L g2137 ( 
.A(n_1954),
.Y(n_2137)
);

AOI22xp33_ASAP7_75t_L g2138 ( 
.A1(n_1950),
.A2(n_1142),
.B1(n_1145),
.B2(n_1130),
.Y(n_2138)
);

BUFx3_ASAP7_75t_L g2139 ( 
.A(n_1954),
.Y(n_2139)
);

AND2x4_ASAP7_75t_L g2140 ( 
.A(n_2041),
.B(n_457),
.Y(n_2140)
);

INVx3_ASAP7_75t_L g2141 ( 
.A(n_2007),
.Y(n_2141)
);

AND2x4_ASAP7_75t_L g2142 ( 
.A(n_2046),
.B(n_2030),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_1961),
.B(n_1262),
.Y(n_2143)
);

INVx2_ASAP7_75t_SL g2144 ( 
.A(n_2007),
.Y(n_2144)
);

HB1xp67_ASAP7_75t_L g2145 ( 
.A(n_1974),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1924),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_1932),
.Y(n_2147)
);

AOI22xp5_ASAP7_75t_L g2148 ( 
.A1(n_1990),
.A2(n_1314),
.B1(n_1315),
.B2(n_1311),
.Y(n_2148)
);

BUFx2_ASAP7_75t_L g2149 ( 
.A(n_1974),
.Y(n_2149)
);

HB1xp67_ASAP7_75t_L g2150 ( 
.A(n_1986),
.Y(n_2150)
);

INVx3_ASAP7_75t_L g2151 ( 
.A(n_1986),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_1959),
.B(n_1266),
.Y(n_2152)
);

AND2x4_ASAP7_75t_L g2153 ( 
.A(n_1943),
.B(n_1960),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1946),
.Y(n_2154)
);

BUFx2_ASAP7_75t_SL g2155 ( 
.A(n_1947),
.Y(n_2155)
);

NAND2x1p5_ASAP7_75t_L g2156 ( 
.A(n_1947),
.B(n_465),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2032),
.B(n_1268),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1975),
.Y(n_2158)
);

AOI21xp33_ASAP7_75t_L g2159 ( 
.A1(n_2003),
.A2(n_1277),
.B(n_1273),
.Y(n_2159)
);

INVx2_ASAP7_75t_SL g2160 ( 
.A(n_2050),
.Y(n_2160)
);

HB1xp67_ASAP7_75t_L g2161 ( 
.A(n_2012),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_1992),
.Y(n_2162)
);

INVx5_ASAP7_75t_L g2163 ( 
.A(n_2012),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_2016),
.Y(n_2164)
);

BUFx6f_ASAP7_75t_L g2165 ( 
.A(n_2017),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2038),
.Y(n_2166)
);

BUFx6f_ASAP7_75t_L g2167 ( 
.A(n_2017),
.Y(n_2167)
);

AND3x2_ASAP7_75t_L g2168 ( 
.A(n_2040),
.B(n_0),
.C(n_2),
.Y(n_2168)
);

AND2x6_ASAP7_75t_L g2169 ( 
.A(n_2037),
.B(n_458),
.Y(n_2169)
);

AOI21xp5_ASAP7_75t_L g2170 ( 
.A1(n_2028),
.A2(n_1971),
.B(n_1988),
.Y(n_2170)
);

A2O1A1Ixp33_ASAP7_75t_L g2171 ( 
.A1(n_1991),
.A2(n_1150),
.B(n_1152),
.C(n_1148),
.Y(n_2171)
);

BUFx6f_ASAP7_75t_L g2172 ( 
.A(n_2025),
.Y(n_2172)
);

INVx3_ASAP7_75t_L g2173 ( 
.A(n_2039),
.Y(n_2173)
);

A2O1A1Ixp33_ASAP7_75t_L g2174 ( 
.A1(n_1998),
.A2(n_1164),
.B(n_1166),
.C(n_1162),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_2053),
.Y(n_2175)
);

AOI21xp5_ASAP7_75t_L g2176 ( 
.A1(n_1993),
.A2(n_1175),
.B(n_1172),
.Y(n_2176)
);

AOI22xp33_ASAP7_75t_L g2177 ( 
.A1(n_1965),
.A2(n_1917),
.B1(n_1941),
.B2(n_2029),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2026),
.Y(n_2178)
);

BUFx6f_ASAP7_75t_L g2179 ( 
.A(n_2025),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2010),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_2004),
.B(n_1173),
.Y(n_2181)
);

BUFx6f_ASAP7_75t_L g2182 ( 
.A(n_2039),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2014),
.Y(n_2183)
);

BUFx6f_ASAP7_75t_L g2184 ( 
.A(n_2048),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_1938),
.Y(n_2185)
);

AND2x6_ASAP7_75t_L g2186 ( 
.A(n_2052),
.B(n_460),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_1951),
.B(n_1177),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_1978),
.B(n_1285),
.Y(n_2188)
);

BUFx2_ASAP7_75t_L g2189 ( 
.A(n_2036),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_1944),
.B(n_1291),
.Y(n_2190)
);

BUFx2_ASAP7_75t_L g2191 ( 
.A(n_2022),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_1952),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_1958),
.Y(n_2193)
);

NOR2x1_ASAP7_75t_SL g2194 ( 
.A(n_2015),
.B(n_461),
.Y(n_2194)
);

AOI221xp5_ASAP7_75t_L g2195 ( 
.A1(n_1909),
.A2(n_1302),
.B1(n_1303),
.B2(n_1301),
.C(n_1295),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_1962),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1957),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1957),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2031),
.Y(n_2199)
);

AOI21xp33_ASAP7_75t_L g2200 ( 
.A1(n_2033),
.A2(n_1313),
.B(n_1182),
.Y(n_2200)
);

NOR2xp33_ASAP7_75t_L g2201 ( 
.A(n_1968),
.B(n_1179),
.Y(n_2201)
);

BUFx10_ASAP7_75t_L g2202 ( 
.A(n_1939),
.Y(n_2202)
);

AOI222xp33_ASAP7_75t_L g2203 ( 
.A1(n_1956),
.A2(n_1199),
.B1(n_1191),
.B2(n_1201),
.C1(n_1198),
.C2(n_1188),
.Y(n_2203)
);

NOR2xp33_ASAP7_75t_L g2204 ( 
.A(n_2049),
.B(n_1212),
.Y(n_2204)
);

BUFx6f_ASAP7_75t_L g2205 ( 
.A(n_1916),
.Y(n_2205)
);

A2O1A1Ixp33_ASAP7_75t_L g2206 ( 
.A1(n_2177),
.A2(n_2024),
.B(n_1929),
.C(n_1214),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2199),
.B(n_1953),
.Y(n_2207)
);

OAI21x1_ASAP7_75t_L g2208 ( 
.A1(n_2128),
.A2(n_463),
.B(n_462),
.Y(n_2208)
);

INVx2_ASAP7_75t_SL g2209 ( 
.A(n_2163),
.Y(n_2209)
);

AO31x2_ASAP7_75t_L g2210 ( 
.A1(n_2065),
.A2(n_466),
.A3(n_469),
.B(n_464),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_2188),
.B(n_1213),
.Y(n_2211)
);

INVx3_ASAP7_75t_SL g2212 ( 
.A(n_2091),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_2068),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_2076),
.Y(n_2214)
);

OAI21x1_ASAP7_75t_L g2215 ( 
.A1(n_2059),
.A2(n_472),
.B(n_471),
.Y(n_2215)
);

AO21x2_ASAP7_75t_L g2216 ( 
.A1(n_2134),
.A2(n_1222),
.B(n_1221),
.Y(n_2216)
);

INVxp67_ASAP7_75t_L g2217 ( 
.A(n_2060),
.Y(n_2217)
);

O2A1O1Ixp5_ASAP7_75t_L g2218 ( 
.A1(n_2103),
.A2(n_1225),
.B(n_1226),
.C(n_1223),
.Y(n_2218)
);

NOR2xp33_ASAP7_75t_L g2219 ( 
.A(n_2185),
.B(n_1229),
.Y(n_2219)
);

OAI21x1_ASAP7_75t_L g2220 ( 
.A1(n_2130),
.A2(n_2170),
.B(n_2119),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2083),
.Y(n_2221)
);

OAI21x1_ASAP7_75t_L g2222 ( 
.A1(n_2121),
.A2(n_474),
.B(n_473),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2152),
.B(n_1232),
.Y(n_2223)
);

INVx6_ASAP7_75t_L g2224 ( 
.A(n_2072),
.Y(n_2224)
);

OAI22xp5_ASAP7_75t_L g2225 ( 
.A1(n_2064),
.A2(n_1236),
.B1(n_1249),
.B2(n_1235),
.Y(n_2225)
);

OAI21x1_ASAP7_75t_L g2226 ( 
.A1(n_2089),
.A2(n_480),
.B(n_476),
.Y(n_2226)
);

NAND2x1p5_ASAP7_75t_L g2227 ( 
.A(n_2163),
.B(n_481),
.Y(n_2227)
);

OA21x2_ASAP7_75t_L g2228 ( 
.A1(n_2133),
.A2(n_2099),
.B(n_2117),
.Y(n_2228)
);

AND2x4_ASAP7_75t_L g2229 ( 
.A(n_2105),
.B(n_482),
.Y(n_2229)
);

AOI22xp33_ASAP7_75t_SL g2230 ( 
.A1(n_2063),
.A2(n_1253),
.B1(n_1259),
.B2(n_1251),
.Y(n_2230)
);

AND2x2_ASAP7_75t_L g2231 ( 
.A(n_2143),
.B(n_1264),
.Y(n_2231)
);

AO21x2_ASAP7_75t_L g2232 ( 
.A1(n_2082),
.A2(n_1272),
.B(n_1267),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2092),
.Y(n_2233)
);

AOI22xp33_ASAP7_75t_L g2234 ( 
.A1(n_2159),
.A2(n_1321),
.B1(n_1276),
.B2(n_1278),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2192),
.B(n_1275),
.Y(n_2235)
);

A2O1A1Ixp33_ASAP7_75t_L g2236 ( 
.A1(n_2055),
.A2(n_1287),
.B(n_1288),
.C(n_1281),
.Y(n_2236)
);

NOR2xp33_ASAP7_75t_R g2237 ( 
.A(n_2061),
.B(n_1289),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2098),
.Y(n_2238)
);

AOI22xp33_ASAP7_75t_L g2239 ( 
.A1(n_2124),
.A2(n_1310),
.B1(n_1290),
.B2(n_1296),
.Y(n_2239)
);

OAI21x1_ASAP7_75t_L g2240 ( 
.A1(n_2085),
.A2(n_484),
.B(n_483),
.Y(n_2240)
);

OA21x2_ASAP7_75t_L g2241 ( 
.A1(n_2069),
.A2(n_1297),
.B(n_1294),
.Y(n_2241)
);

INVx2_ASAP7_75t_SL g2242 ( 
.A(n_2087),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2058),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2070),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2071),
.Y(n_2245)
);

OAI21xp5_ASAP7_75t_L g2246 ( 
.A1(n_2101),
.A2(n_1304),
.B(n_1298),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2074),
.Y(n_2247)
);

BUFx3_ASAP7_75t_L g2248 ( 
.A(n_2165),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_2112),
.Y(n_2249)
);

OAI21x1_ASAP7_75t_L g2250 ( 
.A1(n_2122),
.A2(n_488),
.B(n_487),
.Y(n_2250)
);

INVx2_ASAP7_75t_L g2251 ( 
.A(n_2146),
.Y(n_2251)
);

BUFx3_ASAP7_75t_L g2252 ( 
.A(n_2165),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2075),
.Y(n_2253)
);

OAI21x1_ASAP7_75t_L g2254 ( 
.A1(n_2123),
.A2(n_490),
.B(n_489),
.Y(n_2254)
);

OAI21xp33_ASAP7_75t_SL g2255 ( 
.A1(n_2054),
.A2(n_492),
.B(n_491),
.Y(n_2255)
);

NOR2xp33_ASAP7_75t_L g2256 ( 
.A(n_2193),
.B(n_1305),
.Y(n_2256)
);

OAI21x1_ASAP7_75t_L g2257 ( 
.A1(n_2125),
.A2(n_494),
.B(n_493),
.Y(n_2257)
);

INVxp67_ASAP7_75t_L g2258 ( 
.A(n_2078),
.Y(n_2258)
);

INVx1_ASAP7_75t_SL g2259 ( 
.A(n_2102),
.Y(n_2259)
);

OAI21x1_ASAP7_75t_L g2260 ( 
.A1(n_2126),
.A2(n_496),
.B(n_495),
.Y(n_2260)
);

O2A1O1Ixp33_ASAP7_75t_L g2261 ( 
.A1(n_2110),
.A2(n_4),
.B(n_0),
.C(n_3),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2080),
.Y(n_2262)
);

OAI21xp5_ASAP7_75t_L g2263 ( 
.A1(n_2180),
.A2(n_1307),
.B(n_5),
.Y(n_2263)
);

AND2x4_ASAP7_75t_SL g2264 ( 
.A(n_2067),
.B(n_498),
.Y(n_2264)
);

OAI22xp5_ASAP7_75t_L g2265 ( 
.A1(n_2077),
.A2(n_9),
.B1(n_5),
.B2(n_7),
.Y(n_2265)
);

OAI21x1_ASAP7_75t_L g2266 ( 
.A1(n_2166),
.A2(n_501),
.B(n_500),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_2157),
.B(n_7),
.Y(n_2267)
);

OR2x6_ASAP7_75t_L g2268 ( 
.A(n_2155),
.B(n_503),
.Y(n_2268)
);

NOR3xp33_ASAP7_75t_L g2269 ( 
.A(n_2084),
.B(n_9),
.C(n_11),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_2147),
.Y(n_2270)
);

INVxp67_ASAP7_75t_L g2271 ( 
.A(n_2079),
.Y(n_2271)
);

OAI21x1_ASAP7_75t_L g2272 ( 
.A1(n_2118),
.A2(n_506),
.B(n_504),
.Y(n_2272)
);

A2O1A1Ixp33_ASAP7_75t_L g2273 ( 
.A1(n_2183),
.A2(n_13),
.B(n_11),
.C(n_12),
.Y(n_2273)
);

OAI21x1_ASAP7_75t_L g2274 ( 
.A1(n_2094),
.A2(n_511),
.B(n_508),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2100),
.Y(n_2275)
);

AO31x2_ASAP7_75t_L g2276 ( 
.A1(n_2194),
.A2(n_2171),
.A3(n_2174),
.B(n_2135),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2108),
.Y(n_2277)
);

AND2x4_ASAP7_75t_L g2278 ( 
.A(n_2160),
.B(n_512),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2154),
.Y(n_2279)
);

AO21x2_ASAP7_75t_L g2280 ( 
.A1(n_2181),
.A2(n_516),
.B(n_514),
.Y(n_2280)
);

AOI22xp33_ASAP7_75t_L g2281 ( 
.A1(n_2196),
.A2(n_15),
.B1(n_12),
.B2(n_14),
.Y(n_2281)
);

OAI21x1_ASAP7_75t_L g2282 ( 
.A1(n_2136),
.A2(n_518),
.B(n_517),
.Y(n_2282)
);

OR2x6_ASAP7_75t_L g2283 ( 
.A(n_2057),
.B(n_520),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_2190),
.B(n_14),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2158),
.Y(n_2285)
);

AO21x2_ASAP7_75t_L g2286 ( 
.A1(n_2090),
.A2(n_522),
.B(n_521),
.Y(n_2286)
);

NOR2xp33_ASAP7_75t_SL g2287 ( 
.A(n_2081),
.B(n_525),
.Y(n_2287)
);

OAI21x1_ASAP7_75t_L g2288 ( 
.A1(n_2162),
.A2(n_527),
.B(n_526),
.Y(n_2288)
);

OR2x6_ASAP7_75t_L g2289 ( 
.A(n_2086),
.B(n_528),
.Y(n_2289)
);

OAI22xp5_ASAP7_75t_L g2290 ( 
.A1(n_2073),
.A2(n_2138),
.B1(n_2107),
.B2(n_2178),
.Y(n_2290)
);

OAI21x1_ASAP7_75t_L g2291 ( 
.A1(n_2164),
.A2(n_530),
.B(n_529),
.Y(n_2291)
);

AO21x2_ASAP7_75t_L g2292 ( 
.A1(n_2187),
.A2(n_533),
.B(n_532),
.Y(n_2292)
);

NAND2x1p5_ASAP7_75t_L g2293 ( 
.A(n_2167),
.B(n_534),
.Y(n_2293)
);

OAI22xp5_ASAP7_75t_L g2294 ( 
.A1(n_2111),
.A2(n_18),
.B1(n_15),
.B2(n_17),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_2104),
.B(n_18),
.Y(n_2295)
);

AOI22xp33_ASAP7_75t_L g2296 ( 
.A1(n_2200),
.A2(n_2204),
.B1(n_2186),
.B2(n_2202),
.Y(n_2296)
);

AO21x2_ASAP7_75t_L g2297 ( 
.A1(n_2176),
.A2(n_537),
.B(n_536),
.Y(n_2297)
);

OAI22xp33_ASAP7_75t_L g2298 ( 
.A1(n_2088),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2175),
.Y(n_2299)
);

AOI21x1_ASAP7_75t_L g2300 ( 
.A1(n_2197),
.A2(n_539),
.B(n_538),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2189),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2113),
.Y(n_2302)
);

BUFx3_ASAP7_75t_L g2303 ( 
.A(n_2167),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_2182),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_2182),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2198),
.Y(n_2306)
);

CKINVDCx11_ASAP7_75t_R g2307 ( 
.A(n_2127),
.Y(n_2307)
);

AOI21xp5_ASAP7_75t_L g2308 ( 
.A1(n_2201),
.A2(n_857),
.B(n_856),
.Y(n_2308)
);

AOI21x1_ASAP7_75t_L g2309 ( 
.A1(n_2096),
.A2(n_541),
.B(n_540),
.Y(n_2309)
);

BUFx6f_ASAP7_75t_L g2310 ( 
.A(n_2248),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2243),
.Y(n_2311)
);

AOI22xp33_ASAP7_75t_L g2312 ( 
.A1(n_2269),
.A2(n_2186),
.B1(n_2169),
.B2(n_2131),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2228),
.B(n_2114),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_2213),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_2214),
.Y(n_2315)
);

AND2x4_ASAP7_75t_L g2316 ( 
.A(n_2258),
.B(n_2142),
.Y(n_2316)
);

AND2x2_ASAP7_75t_L g2317 ( 
.A(n_2284),
.B(n_2129),
.Y(n_2317)
);

OAI22xp33_ASAP7_75t_L g2318 ( 
.A1(n_2263),
.A2(n_2156),
.B1(n_2148),
.B2(n_2191),
.Y(n_2318)
);

AOI21xp5_ASAP7_75t_L g2319 ( 
.A1(n_2220),
.A2(n_2308),
.B(n_2206),
.Y(n_2319)
);

NAND2x1p5_ASAP7_75t_L g2320 ( 
.A(n_2259),
.B(n_2095),
.Y(n_2320)
);

OAI22xp5_ASAP7_75t_L g2321 ( 
.A1(n_2296),
.A2(n_2239),
.B1(n_2295),
.B2(n_2290),
.Y(n_2321)
);

CKINVDCx20_ASAP7_75t_R g2322 ( 
.A(n_2307),
.Y(n_2322)
);

CKINVDCx5p33_ASAP7_75t_R g2323 ( 
.A(n_2212),
.Y(n_2323)
);

OAI222xp33_ASAP7_75t_L g2324 ( 
.A1(n_2298),
.A2(n_2062),
.B1(n_2120),
.B2(n_2168),
.C1(n_2140),
.C2(n_2161),
.Y(n_2324)
);

INVx6_ASAP7_75t_L g2325 ( 
.A(n_2252),
.Y(n_2325)
);

OAI21xp5_ASAP7_75t_L g2326 ( 
.A1(n_2236),
.A2(n_2203),
.B(n_2195),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2244),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2245),
.Y(n_2328)
);

INVx2_ASAP7_75t_SL g2329 ( 
.A(n_2303),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2247),
.Y(n_2330)
);

OR2x6_ASAP7_75t_L g2331 ( 
.A(n_2268),
.B(n_2184),
.Y(n_2331)
);

AOI221xp5_ASAP7_75t_L g2332 ( 
.A1(n_2265),
.A2(n_2145),
.B1(n_2150),
.B2(n_2137),
.C(n_2116),
.Y(n_2332)
);

AOI22xp33_ASAP7_75t_L g2333 ( 
.A1(n_2267),
.A2(n_2186),
.B1(n_2169),
.B2(n_2093),
.Y(n_2333)
);

INVx3_ASAP7_75t_L g2334 ( 
.A(n_2304),
.Y(n_2334)
);

BUFx2_ASAP7_75t_L g2335 ( 
.A(n_2217),
.Y(n_2335)
);

AOI211xp5_ASAP7_75t_L g2336 ( 
.A1(n_2294),
.A2(n_2132),
.B(n_2115),
.C(n_2205),
.Y(n_2336)
);

NOR2xp33_ASAP7_75t_L g2337 ( 
.A(n_2271),
.B(n_2066),
.Y(n_2337)
);

AOI22xp33_ASAP7_75t_L g2338 ( 
.A1(n_2225),
.A2(n_2169),
.B1(n_2205),
.B2(n_2184),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2253),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2262),
.Y(n_2340)
);

OAI22xp33_ASAP7_75t_L g2341 ( 
.A1(n_2287),
.A2(n_2056),
.B1(n_2179),
.B2(n_2172),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_2249),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_2251),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2299),
.B(n_2149),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2275),
.Y(n_2345)
);

AOI221xp5_ASAP7_75t_SL g2346 ( 
.A1(n_2261),
.A2(n_2273),
.B1(n_2281),
.B2(n_2246),
.C(n_2255),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_2270),
.Y(n_2347)
);

OAI22xp5_ASAP7_75t_L g2348 ( 
.A1(n_2230),
.A2(n_2179),
.B1(n_2172),
.B2(n_2153),
.Y(n_2348)
);

AOI22xp33_ASAP7_75t_L g2349 ( 
.A1(n_2219),
.A2(n_2141),
.B1(n_2139),
.B2(n_2151),
.Y(n_2349)
);

OAI21x1_ASAP7_75t_L g2350 ( 
.A1(n_2215),
.A2(n_2173),
.B(n_543),
.Y(n_2350)
);

AOI21xp5_ASAP7_75t_L g2351 ( 
.A1(n_2216),
.A2(n_2144),
.B(n_2106),
.Y(n_2351)
);

BUFx2_ASAP7_75t_L g2352 ( 
.A(n_2301),
.Y(n_2352)
);

AOI22xp33_ASAP7_75t_SL g2353 ( 
.A1(n_2286),
.A2(n_2106),
.B1(n_2109),
.B2(n_2097),
.Y(n_2353)
);

NAND2xp33_ASAP7_75t_SL g2354 ( 
.A(n_2237),
.B(n_2097),
.Y(n_2354)
);

INVx4_ASAP7_75t_L g2355 ( 
.A(n_2224),
.Y(n_2355)
);

OAI211xp5_ASAP7_75t_L g2356 ( 
.A1(n_2234),
.A2(n_2109),
.B(n_23),
.C(n_19),
.Y(n_2356)
);

AOI22xp5_ASAP7_75t_L g2357 ( 
.A1(n_2256),
.A2(n_24),
.B1(n_20),
.B2(n_23),
.Y(n_2357)
);

CKINVDCx11_ASAP7_75t_R g2358 ( 
.A(n_2305),
.Y(n_2358)
);

OAI22xp5_ASAP7_75t_L g2359 ( 
.A1(n_2207),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_2359)
);

AOI22xp33_ASAP7_75t_L g2360 ( 
.A1(n_2289),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2277),
.Y(n_2361)
);

AND2x2_ASAP7_75t_L g2362 ( 
.A(n_2279),
.B(n_542),
.Y(n_2362)
);

OAI221xp5_ASAP7_75t_L g2363 ( 
.A1(n_2235),
.A2(n_30),
.B1(n_27),
.B2(n_28),
.C(n_31),
.Y(n_2363)
);

INVx3_ASAP7_75t_L g2364 ( 
.A(n_2209),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2285),
.Y(n_2365)
);

AND2x4_ASAP7_75t_L g2366 ( 
.A(n_2352),
.B(n_2302),
.Y(n_2366)
);

AND2x2_ASAP7_75t_L g2367 ( 
.A(n_2313),
.B(n_2221),
.Y(n_2367)
);

AOI22xp33_ASAP7_75t_L g2368 ( 
.A1(n_2326),
.A2(n_2232),
.B1(n_2241),
.B2(n_2283),
.Y(n_2368)
);

INVx3_ASAP7_75t_SL g2369 ( 
.A(n_2323),
.Y(n_2369)
);

HB1xp67_ASAP7_75t_L g2370 ( 
.A(n_2365),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_2311),
.Y(n_2371)
);

OR2x6_ASAP7_75t_L g2372 ( 
.A(n_2331),
.B(n_2320),
.Y(n_2372)
);

BUFx6f_ASAP7_75t_L g2373 ( 
.A(n_2310),
.Y(n_2373)
);

NAND2xp33_ASAP7_75t_R g2374 ( 
.A(n_2331),
.B(n_2283),
.Y(n_2374)
);

CKINVDCx5p33_ASAP7_75t_R g2375 ( 
.A(n_2322),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2314),
.B(n_2233),
.Y(n_2376)
);

OAI21xp33_ASAP7_75t_L g2377 ( 
.A1(n_2357),
.A2(n_2211),
.B(n_2223),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2327),
.Y(n_2378)
);

AOI22xp33_ASAP7_75t_L g2379 ( 
.A1(n_2321),
.A2(n_2289),
.B1(n_2268),
.B2(n_2292),
.Y(n_2379)
);

AND2x2_ASAP7_75t_L g2380 ( 
.A(n_2317),
.B(n_2238),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2328),
.Y(n_2381)
);

AND2x2_ASAP7_75t_L g2382 ( 
.A(n_2330),
.B(n_2306),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2315),
.B(n_2231),
.Y(n_2383)
);

HB1xp67_ASAP7_75t_L g2384 ( 
.A(n_2339),
.Y(n_2384)
);

INVxp67_ASAP7_75t_L g2385 ( 
.A(n_2335),
.Y(n_2385)
);

AND2x2_ASAP7_75t_L g2386 ( 
.A(n_2340),
.B(n_2222),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2345),
.Y(n_2387)
);

CKINVDCx16_ASAP7_75t_R g2388 ( 
.A(n_2355),
.Y(n_2388)
);

OR2x2_ASAP7_75t_L g2389 ( 
.A(n_2361),
.B(n_2280),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2342),
.B(n_2229),
.Y(n_2390)
);

NOR2xp33_ASAP7_75t_L g2391 ( 
.A(n_2316),
.B(n_2278),
.Y(n_2391)
);

CKINVDCx5p33_ASAP7_75t_R g2392 ( 
.A(n_2358),
.Y(n_2392)
);

OR2x2_ASAP7_75t_L g2393 ( 
.A(n_2344),
.B(n_2226),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2343),
.Y(n_2394)
);

NOR3xp33_ASAP7_75t_SL g2395 ( 
.A(n_2363),
.B(n_2218),
.C(n_2264),
.Y(n_2395)
);

NAND2x1p5_ASAP7_75t_L g2396 ( 
.A(n_2364),
.B(n_2240),
.Y(n_2396)
);

AOI22xp33_ASAP7_75t_L g2397 ( 
.A1(n_2312),
.A2(n_2297),
.B1(n_2227),
.B2(n_2293),
.Y(n_2397)
);

NAND3xp33_ASAP7_75t_L g2398 ( 
.A(n_2346),
.B(n_2242),
.C(n_2276),
.Y(n_2398)
);

OR2x2_ASAP7_75t_L g2399 ( 
.A(n_2347),
.B(n_2210),
.Y(n_2399)
);

NAND2xp33_ASAP7_75t_SL g2400 ( 
.A(n_2360),
.B(n_2309),
.Y(n_2400)
);

HB1xp67_ASAP7_75t_L g2401 ( 
.A(n_2334),
.Y(n_2401)
);

INVxp67_ASAP7_75t_SL g2402 ( 
.A(n_2319),
.Y(n_2402)
);

AO31x2_ASAP7_75t_L g2403 ( 
.A1(n_2359),
.A2(n_2210),
.A3(n_2300),
.B(n_2208),
.Y(n_2403)
);

AOI22xp33_ASAP7_75t_L g2404 ( 
.A1(n_2318),
.A2(n_2274),
.B1(n_2254),
.B2(n_2257),
.Y(n_2404)
);

INVx1_ASAP7_75t_SL g2405 ( 
.A(n_2325),
.Y(n_2405)
);

NOR3xp33_ASAP7_75t_SL g2406 ( 
.A(n_2324),
.B(n_2276),
.C(n_2260),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2362),
.Y(n_2407)
);

OR2x6_ASAP7_75t_L g2408 ( 
.A(n_2351),
.B(n_2250),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2353),
.Y(n_2409)
);

OR2x2_ASAP7_75t_L g2410 ( 
.A(n_2337),
.B(n_2266),
.Y(n_2410)
);

NAND2xp33_ASAP7_75t_R g2411 ( 
.A(n_2354),
.B(n_2272),
.Y(n_2411)
);

CKINVDCx5p33_ASAP7_75t_R g2412 ( 
.A(n_2310),
.Y(n_2412)
);

OR2x6_ASAP7_75t_L g2413 ( 
.A(n_2329),
.B(n_2282),
.Y(n_2413)
);

AND2x2_ASAP7_75t_L g2414 ( 
.A(n_2333),
.B(n_2288),
.Y(n_2414)
);

AND2x4_ASAP7_75t_L g2415 ( 
.A(n_2349),
.B(n_2291),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_SL g2416 ( 
.A(n_2341),
.B(n_544),
.Y(n_2416)
);

AND2x4_ASAP7_75t_L g2417 ( 
.A(n_2338),
.B(n_545),
.Y(n_2417)
);

NAND2xp33_ASAP7_75t_R g2418 ( 
.A(n_2350),
.B(n_31),
.Y(n_2418)
);

CKINVDCx20_ASAP7_75t_R g2419 ( 
.A(n_2325),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2348),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2332),
.Y(n_2421)
);

INVx2_ASAP7_75t_L g2422 ( 
.A(n_2356),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2336),
.Y(n_2423)
);

NOR3xp33_ASAP7_75t_SL g2424 ( 
.A(n_2363),
.B(n_33),
.C(n_34),
.Y(n_2424)
);

NOR2xp33_ASAP7_75t_R g2425 ( 
.A(n_2322),
.B(n_546),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2370),
.Y(n_2426)
);

HB1xp67_ASAP7_75t_L g2427 ( 
.A(n_2384),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2378),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2381),
.Y(n_2429)
);

INVx2_ASAP7_75t_SL g2430 ( 
.A(n_2373),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2387),
.Y(n_2431)
);

BUFx3_ASAP7_75t_L g2432 ( 
.A(n_2419),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2371),
.Y(n_2433)
);

AND2x2_ASAP7_75t_L g2434 ( 
.A(n_2367),
.B(n_33),
.Y(n_2434)
);

INVxp67_ASAP7_75t_L g2435 ( 
.A(n_2401),
.Y(n_2435)
);

AND2x2_ASAP7_75t_L g2436 ( 
.A(n_2385),
.B(n_34),
.Y(n_2436)
);

AND2x2_ASAP7_75t_L g2437 ( 
.A(n_2366),
.B(n_35),
.Y(n_2437)
);

AND2x2_ASAP7_75t_L g2438 ( 
.A(n_2380),
.B(n_2382),
.Y(n_2438)
);

AND2x2_ASAP7_75t_L g2439 ( 
.A(n_2372),
.B(n_35),
.Y(n_2439)
);

AND2x2_ASAP7_75t_L g2440 ( 
.A(n_2372),
.B(n_36),
.Y(n_2440)
);

AND2x2_ASAP7_75t_L g2441 ( 
.A(n_2405),
.B(n_36),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2394),
.B(n_38),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2389),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2399),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2376),
.Y(n_2445)
);

BUFx6f_ASAP7_75t_L g2446 ( 
.A(n_2373),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_2386),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2393),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2410),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2409),
.Y(n_2450)
);

AO31x2_ASAP7_75t_L g2451 ( 
.A1(n_2421),
.A2(n_40),
.A3(n_38),
.B(n_39),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2407),
.Y(n_2452)
);

HB1xp67_ASAP7_75t_L g2453 ( 
.A(n_2408),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2388),
.B(n_40),
.Y(n_2454)
);

OAI21xp5_ASAP7_75t_SL g2455 ( 
.A1(n_2377),
.A2(n_43),
.B(n_42),
.Y(n_2455)
);

HB1xp67_ASAP7_75t_L g2456 ( 
.A(n_2408),
.Y(n_2456)
);

AND2x2_ASAP7_75t_L g2457 ( 
.A(n_2414),
.B(n_41),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_2383),
.Y(n_2458)
);

INVx2_ASAP7_75t_SL g2459 ( 
.A(n_2412),
.Y(n_2459)
);

OR2x2_ASAP7_75t_L g2460 ( 
.A(n_2402),
.B(n_41),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2398),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2413),
.Y(n_2462)
);

AND2x4_ASAP7_75t_L g2463 ( 
.A(n_2415),
.B(n_42),
.Y(n_2463)
);

AND2x2_ASAP7_75t_L g2464 ( 
.A(n_2369),
.B(n_43),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2420),
.Y(n_2465)
);

OR2x2_ASAP7_75t_L g2466 ( 
.A(n_2390),
.B(n_44),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_2413),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_2403),
.Y(n_2468)
);

INVx2_ASAP7_75t_L g2469 ( 
.A(n_2403),
.Y(n_2469)
);

BUFx3_ASAP7_75t_L g2470 ( 
.A(n_2392),
.Y(n_2470)
);

AND2x2_ASAP7_75t_L g2471 ( 
.A(n_2391),
.B(n_45),
.Y(n_2471)
);

AND2x2_ASAP7_75t_L g2472 ( 
.A(n_2423),
.B(n_45),
.Y(n_2472)
);

AOI22xp33_ASAP7_75t_L g2473 ( 
.A1(n_2400),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_2473)
);

HB1xp67_ASAP7_75t_L g2474 ( 
.A(n_2418),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2396),
.Y(n_2475)
);

AND2x2_ASAP7_75t_L g2476 ( 
.A(n_2422),
.B(n_47),
.Y(n_2476)
);

INVx1_ASAP7_75t_SL g2477 ( 
.A(n_2375),
.Y(n_2477)
);

AND2x2_ASAP7_75t_L g2478 ( 
.A(n_2379),
.B(n_48),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2417),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2406),
.Y(n_2480)
);

OR2x2_ASAP7_75t_L g2481 ( 
.A(n_2404),
.B(n_49),
.Y(n_2481)
);

INVx2_ASAP7_75t_L g2482 ( 
.A(n_2416),
.Y(n_2482)
);

INVx4_ASAP7_75t_L g2483 ( 
.A(n_2374),
.Y(n_2483)
);

HB1xp67_ASAP7_75t_L g2484 ( 
.A(n_2411),
.Y(n_2484)
);

INVx3_ASAP7_75t_L g2485 ( 
.A(n_2425),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_2424),
.B(n_49),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2368),
.Y(n_2487)
);

AND2x2_ASAP7_75t_L g2488 ( 
.A(n_2397),
.B(n_50),
.Y(n_2488)
);

AND2x2_ASAP7_75t_L g2489 ( 
.A(n_2395),
.B(n_51),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_2367),
.B(n_51),
.Y(n_2490)
);

INVxp67_ASAP7_75t_R g2491 ( 
.A(n_2367),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_2371),
.Y(n_2492)
);

OR2x2_ASAP7_75t_L g2493 ( 
.A(n_2370),
.B(n_52),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_2371),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2371),
.Y(n_2495)
);

AND2x2_ASAP7_75t_L g2496 ( 
.A(n_2367),
.B(n_52),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2371),
.Y(n_2497)
);

AND2x2_ASAP7_75t_L g2498 ( 
.A(n_2367),
.B(n_53),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2370),
.Y(n_2499)
);

INVx2_ASAP7_75t_L g2500 ( 
.A(n_2371),
.Y(n_2500)
);

OAI21xp5_ASAP7_75t_L g2501 ( 
.A1(n_2368),
.A2(n_53),
.B(n_54),
.Y(n_2501)
);

AND2x2_ASAP7_75t_L g2502 ( 
.A(n_2367),
.B(n_54),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2371),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2370),
.Y(n_2504)
);

BUFx3_ASAP7_75t_L g2505 ( 
.A(n_2419),
.Y(n_2505)
);

INVx2_ASAP7_75t_L g2506 ( 
.A(n_2371),
.Y(n_2506)
);

OR2x2_ASAP7_75t_L g2507 ( 
.A(n_2370),
.B(n_55),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2370),
.Y(n_2508)
);

OAI22xp5_ASAP7_75t_L g2509 ( 
.A1(n_2473),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_2509)
);

OAI221xp5_ASAP7_75t_L g2510 ( 
.A1(n_2501),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.C(n_59),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2450),
.B(n_58),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_2491),
.B(n_2438),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_L g2513 ( 
.A(n_2445),
.B(n_59),
.Y(n_2513)
);

AND2x2_ASAP7_75t_L g2514 ( 
.A(n_2491),
.B(n_2435),
.Y(n_2514)
);

OA211x2_ASAP7_75t_L g2515 ( 
.A1(n_2486),
.A2(n_62),
.B(n_60),
.C(n_61),
.Y(n_2515)
);

OAI22xp5_ASAP7_75t_L g2516 ( 
.A1(n_2474),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_2516)
);

NAND3xp33_ASAP7_75t_L g2517 ( 
.A(n_2461),
.B(n_63),
.C(n_65),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2448),
.B(n_63),
.Y(n_2518)
);

OAI22xp5_ASAP7_75t_L g2519 ( 
.A1(n_2455),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_2519)
);

OAI22xp5_ASAP7_75t_L g2520 ( 
.A1(n_2482),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_2520)
);

NOR3xp33_ASAP7_75t_L g2521 ( 
.A(n_2487),
.B(n_68),
.C(n_69),
.Y(n_2521)
);

OAI21xp33_ASAP7_75t_L g2522 ( 
.A1(n_2481),
.A2(n_70),
.B(n_71),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2458),
.B(n_71),
.Y(n_2523)
);

OAI221xp5_ASAP7_75t_SL g2524 ( 
.A1(n_2489),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.C(n_75),
.Y(n_2524)
);

AND2x2_ASAP7_75t_L g2525 ( 
.A(n_2483),
.B(n_72),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2428),
.Y(n_2526)
);

AOI221xp5_ASAP7_75t_L g2527 ( 
.A1(n_2478),
.A2(n_2488),
.B1(n_2480),
.B2(n_2476),
.C(n_2472),
.Y(n_2527)
);

AND2x2_ASAP7_75t_L g2528 ( 
.A(n_2427),
.B(n_73),
.Y(n_2528)
);

AND2x2_ASAP7_75t_L g2529 ( 
.A(n_2449),
.B(n_74),
.Y(n_2529)
);

OAI22xp5_ASAP7_75t_L g2530 ( 
.A1(n_2479),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2426),
.B(n_78),
.Y(n_2531)
);

OAI21xp33_ASAP7_75t_L g2532 ( 
.A1(n_2460),
.A2(n_78),
.B(n_79),
.Y(n_2532)
);

OAI21xp33_ASAP7_75t_L g2533 ( 
.A1(n_2457),
.A2(n_2484),
.B(n_2463),
.Y(n_2533)
);

AND2x2_ASAP7_75t_L g2534 ( 
.A(n_2467),
.B(n_79),
.Y(n_2534)
);

AND2x2_ASAP7_75t_L g2535 ( 
.A(n_2499),
.B(n_80),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2504),
.B(n_81),
.Y(n_2536)
);

NAND3xp33_ASAP7_75t_L g2537 ( 
.A(n_2453),
.B(n_82),
.C(n_83),
.Y(n_2537)
);

AOI221xp5_ASAP7_75t_L g2538 ( 
.A1(n_2442),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.C(n_85),
.Y(n_2538)
);

AOI22xp33_ASAP7_75t_L g2539 ( 
.A1(n_2463),
.A2(n_87),
.B1(n_84),
.B2(n_86),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_2508),
.B(n_88),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_2452),
.B(n_88),
.Y(n_2541)
);

AOI221xp5_ASAP7_75t_L g2542 ( 
.A1(n_2443),
.A2(n_2490),
.B1(n_2498),
.B2(n_2496),
.C(n_2434),
.Y(n_2542)
);

OAI21xp5_ASAP7_75t_L g2543 ( 
.A1(n_2456),
.A2(n_89),
.B(n_90),
.Y(n_2543)
);

NAND3xp33_ASAP7_75t_L g2544 ( 
.A(n_2462),
.B(n_89),
.C(n_90),
.Y(n_2544)
);

OAI22xp5_ASAP7_75t_L g2545 ( 
.A1(n_2465),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_2545)
);

AND2x2_ASAP7_75t_L g2546 ( 
.A(n_2447),
.B(n_91),
.Y(n_2546)
);

AND2x2_ASAP7_75t_L g2547 ( 
.A(n_2462),
.B(n_94),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_SL g2548 ( 
.A(n_2475),
.B(n_2470),
.Y(n_2548)
);

HB1xp67_ASAP7_75t_L g2549 ( 
.A(n_2444),
.Y(n_2549)
);

AND2x2_ASAP7_75t_L g2550 ( 
.A(n_2433),
.B(n_2492),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2494),
.B(n_94),
.Y(n_2551)
);

OAI22xp5_ASAP7_75t_L g2552 ( 
.A1(n_2430),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_2552)
);

OAI22xp5_ASAP7_75t_L g2553 ( 
.A1(n_2507),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_2553)
);

AND2x2_ASAP7_75t_L g2554 ( 
.A(n_2495),
.B(n_98),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_2497),
.B(n_98),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2500),
.B(n_99),
.Y(n_2556)
);

AOI221xp5_ASAP7_75t_L g2557 ( 
.A1(n_2502),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.C(n_102),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2428),
.Y(n_2558)
);

AND2x2_ASAP7_75t_L g2559 ( 
.A(n_2503),
.B(n_101),
.Y(n_2559)
);

OAI21xp33_ASAP7_75t_SL g2560 ( 
.A1(n_2493),
.A2(n_102),
.B(n_103),
.Y(n_2560)
);

NAND3xp33_ASAP7_75t_L g2561 ( 
.A(n_2468),
.B(n_103),
.C(n_104),
.Y(n_2561)
);

OAI22xp5_ASAP7_75t_L g2562 ( 
.A1(n_2466),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_2562)
);

AOI221xp5_ASAP7_75t_L g2563 ( 
.A1(n_2436),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.C(n_108),
.Y(n_2563)
);

NOR2xp33_ASAP7_75t_L g2564 ( 
.A(n_2477),
.B(n_107),
.Y(n_2564)
);

NOR2x1p5_ASAP7_75t_L g2565 ( 
.A(n_2485),
.B(n_2432),
.Y(n_2565)
);

OAI221xp5_ASAP7_75t_L g2566 ( 
.A1(n_2439),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.C(n_111),
.Y(n_2566)
);

AND2x2_ASAP7_75t_L g2567 ( 
.A(n_2506),
.B(n_2431),
.Y(n_2567)
);

OAI21xp33_ASAP7_75t_L g2568 ( 
.A1(n_2440),
.A2(n_109),
.B(n_110),
.Y(n_2568)
);

AND2x2_ASAP7_75t_L g2569 ( 
.A(n_2429),
.B(n_111),
.Y(n_2569)
);

AND2x2_ASAP7_75t_L g2570 ( 
.A(n_2429),
.B(n_112),
.Y(n_2570)
);

NAND4xp25_ASAP7_75t_SL g2571 ( 
.A(n_2454),
.B(n_115),
.C(n_112),
.D(n_113),
.Y(n_2571)
);

AOI221xp5_ASAP7_75t_L g2572 ( 
.A1(n_2441),
.A2(n_116),
.B1(n_113),
.B2(n_115),
.C(n_117),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_L g2573 ( 
.A(n_2437),
.B(n_116),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2469),
.B(n_2471),
.Y(n_2574)
);

AOI22xp33_ASAP7_75t_L g2575 ( 
.A1(n_2464),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_2451),
.B(n_118),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_L g2577 ( 
.A(n_2451),
.B(n_120),
.Y(n_2577)
);

AND2x2_ASAP7_75t_L g2578 ( 
.A(n_2505),
.B(n_121),
.Y(n_2578)
);

NOR3xp33_ASAP7_75t_L g2579 ( 
.A(n_2459),
.B(n_121),
.C(n_122),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_L g2580 ( 
.A(n_2446),
.B(n_122),
.Y(n_2580)
);

NAND3xp33_ASAP7_75t_L g2581 ( 
.A(n_2446),
.B(n_123),
.C(n_124),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_2450),
.B(n_124),
.Y(n_2582)
);

NAND3xp33_ASAP7_75t_L g2583 ( 
.A(n_2461),
.B(n_125),
.C(n_126),
.Y(n_2583)
);

AOI22xp33_ASAP7_75t_L g2584 ( 
.A1(n_2474),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_2584)
);

OAI22xp5_ASAP7_75t_L g2585 ( 
.A1(n_2473),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.Y(n_2585)
);

NAND3xp33_ASAP7_75t_L g2586 ( 
.A(n_2461),
.B(n_128),
.C(n_129),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_SL g2587 ( 
.A(n_2483),
.B(n_130),
.Y(n_2587)
);

NOR3xp33_ASAP7_75t_L g2588 ( 
.A(n_2501),
.B(n_131),
.C(n_132),
.Y(n_2588)
);

OAI22xp5_ASAP7_75t_L g2589 ( 
.A1(n_2473),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_L g2590 ( 
.A(n_2450),
.B(n_134),
.Y(n_2590)
);

AND2x2_ASAP7_75t_L g2591 ( 
.A(n_2491),
.B(n_135),
.Y(n_2591)
);

NAND4xp25_ASAP7_75t_L g2592 ( 
.A(n_2486),
.B(n_138),
.C(n_136),
.D(n_137),
.Y(n_2592)
);

OAI21xp5_ASAP7_75t_SL g2593 ( 
.A1(n_2455),
.A2(n_136),
.B(n_137),
.Y(n_2593)
);

AOI211xp5_ASAP7_75t_L g2594 ( 
.A1(n_2474),
.A2(n_142),
.B(n_139),
.C(n_141),
.Y(n_2594)
);

AND2x2_ASAP7_75t_L g2595 ( 
.A(n_2491),
.B(n_139),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2450),
.B(n_141),
.Y(n_2596)
);

AND2x2_ASAP7_75t_L g2597 ( 
.A(n_2491),
.B(n_142),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_L g2598 ( 
.A(n_2450),
.B(n_143),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_2450),
.B(n_144),
.Y(n_2599)
);

NAND3xp33_ASAP7_75t_L g2600 ( 
.A(n_2461),
.B(n_144),
.C(n_145),
.Y(n_2600)
);

OA211x2_ASAP7_75t_L g2601 ( 
.A1(n_2501),
.A2(n_148),
.B(n_146),
.C(n_147),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_L g2602 ( 
.A(n_2450),
.B(n_146),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2450),
.B(n_148),
.Y(n_2603)
);

AND2x2_ASAP7_75t_L g2604 ( 
.A(n_2491),
.B(n_149),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2491),
.B(n_149),
.Y(n_2605)
);

OAI21xp5_ASAP7_75t_SL g2606 ( 
.A1(n_2455),
.A2(n_150),
.B(n_151),
.Y(n_2606)
);

NOR2xp33_ASAP7_75t_L g2607 ( 
.A(n_2483),
.B(n_150),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_L g2608 ( 
.A(n_2450),
.B(n_151),
.Y(n_2608)
);

NAND3xp33_ASAP7_75t_L g2609 ( 
.A(n_2461),
.B(n_152),
.C(n_153),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_2450),
.B(n_152),
.Y(n_2610)
);

NAND4xp25_ASAP7_75t_L g2611 ( 
.A(n_2486),
.B(n_156),
.C(n_154),
.D(n_155),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2450),
.B(n_154),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2450),
.B(n_157),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_2450),
.B(n_158),
.Y(n_2614)
);

NAND3xp33_ASAP7_75t_L g2615 ( 
.A(n_2461),
.B(n_158),
.C(n_159),
.Y(n_2615)
);

NOR2xp33_ASAP7_75t_SL g2616 ( 
.A(n_2483),
.B(n_159),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2450),
.B(n_160),
.Y(n_2617)
);

OAI21xp33_ASAP7_75t_L g2618 ( 
.A1(n_2473),
.A2(n_162),
.B(n_163),
.Y(n_2618)
);

OAI221xp5_ASAP7_75t_L g2619 ( 
.A1(n_2501),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.C(n_165),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_L g2620 ( 
.A(n_2450),
.B(n_165),
.Y(n_2620)
);

AOI21xp33_ASAP7_75t_L g2621 ( 
.A1(n_2487),
.A2(n_166),
.B(n_167),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_SL g2622 ( 
.A(n_2483),
.B(n_167),
.Y(n_2622)
);

NAND3xp33_ASAP7_75t_L g2623 ( 
.A(n_2461),
.B(n_168),
.C(n_169),
.Y(n_2623)
);

AOI211xp5_ASAP7_75t_L g2624 ( 
.A1(n_2474),
.A2(n_170),
.B(n_168),
.C(n_169),
.Y(n_2624)
);

INVxp67_ASAP7_75t_L g2625 ( 
.A(n_2574),
.Y(n_2625)
);

HB1xp67_ASAP7_75t_L g2626 ( 
.A(n_2549),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_2526),
.Y(n_2627)
);

INVx2_ASAP7_75t_L g2628 ( 
.A(n_2558),
.Y(n_2628)
);

NAND3xp33_ASAP7_75t_L g2629 ( 
.A(n_2594),
.B(n_170),
.C(n_171),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2514),
.Y(n_2630)
);

AND2x2_ASAP7_75t_L g2631 ( 
.A(n_2512),
.B(n_171),
.Y(n_2631)
);

NAND2x1p5_ASAP7_75t_L g2632 ( 
.A(n_2548),
.B(n_172),
.Y(n_2632)
);

INVxp67_ASAP7_75t_L g2633 ( 
.A(n_2607),
.Y(n_2633)
);

AND2x4_ASAP7_75t_L g2634 ( 
.A(n_2565),
.B(n_2567),
.Y(n_2634)
);

AND2x2_ASAP7_75t_L g2635 ( 
.A(n_2550),
.B(n_2533),
.Y(n_2635)
);

AOI22xp33_ASAP7_75t_L g2636 ( 
.A1(n_2588),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2569),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2547),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2570),
.Y(n_2639)
);

INVx2_ASAP7_75t_L g2640 ( 
.A(n_2534),
.Y(n_2640)
);

OR2x2_ASAP7_75t_L g2641 ( 
.A(n_2518),
.B(n_173),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_SL g2642 ( 
.A(n_2527),
.B(n_175),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_L g2643 ( 
.A(n_2528),
.B(n_176),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2531),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2536),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2540),
.Y(n_2646)
);

AND2x2_ASAP7_75t_L g2647 ( 
.A(n_2591),
.B(n_177),
.Y(n_2647)
);

AND2x4_ASAP7_75t_SL g2648 ( 
.A(n_2595),
.B(n_177),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2551),
.Y(n_2649)
);

OR2x2_ASAP7_75t_L g2650 ( 
.A(n_2511),
.B(n_178),
.Y(n_2650)
);

AND2x2_ASAP7_75t_L g2651 ( 
.A(n_2597),
.B(n_178),
.Y(n_2651)
);

AND2x2_ASAP7_75t_L g2652 ( 
.A(n_2604),
.B(n_179),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2529),
.B(n_2535),
.Y(n_2653)
);

BUFx2_ASAP7_75t_L g2654 ( 
.A(n_2605),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2555),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2556),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2541),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2554),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2559),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2546),
.Y(n_2660)
);

OR2x2_ASAP7_75t_L g2661 ( 
.A(n_2582),
.B(n_179),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2513),
.Y(n_2662)
);

AND2x2_ASAP7_75t_L g2663 ( 
.A(n_2542),
.B(n_181),
.Y(n_2663)
);

AND2x2_ASAP7_75t_L g2664 ( 
.A(n_2525),
.B(n_2578),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_L g2665 ( 
.A(n_2523),
.B(n_182),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2590),
.Y(n_2666)
);

NOR2xp33_ASAP7_75t_L g2667 ( 
.A(n_2592),
.B(n_2611),
.Y(n_2667)
);

INVx1_ASAP7_75t_SL g2668 ( 
.A(n_2573),
.Y(n_2668)
);

INVxp67_ASAP7_75t_SL g2669 ( 
.A(n_2576),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2577),
.Y(n_2670)
);

NOR3xp33_ASAP7_75t_L g2671 ( 
.A(n_2510),
.B(n_182),
.C(n_183),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2596),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_2598),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_L g2674 ( 
.A(n_2599),
.B(n_183),
.Y(n_2674)
);

AND2x2_ASAP7_75t_L g2675 ( 
.A(n_2602),
.B(n_184),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2603),
.B(n_185),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2608),
.Y(n_2677)
);

AND2x4_ASAP7_75t_L g2678 ( 
.A(n_2610),
.B(n_185),
.Y(n_2678)
);

AND2x2_ASAP7_75t_L g2679 ( 
.A(n_2612),
.B(n_186),
.Y(n_2679)
);

OR2x2_ASAP7_75t_L g2680 ( 
.A(n_2613),
.B(n_186),
.Y(n_2680)
);

AND2x2_ASAP7_75t_L g2681 ( 
.A(n_2614),
.B(n_2617),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_L g2682 ( 
.A(n_2620),
.B(n_187),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2580),
.Y(n_2683)
);

INVx2_ASAP7_75t_L g2684 ( 
.A(n_2587),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2622),
.Y(n_2685)
);

HB1xp67_ASAP7_75t_L g2686 ( 
.A(n_2560),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_L g2687 ( 
.A(n_2521),
.B(n_189),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2561),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2517),
.Y(n_2689)
);

AND2x2_ASAP7_75t_L g2690 ( 
.A(n_2564),
.B(n_2543),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2532),
.B(n_189),
.Y(n_2691)
);

AND2x2_ASAP7_75t_L g2692 ( 
.A(n_2616),
.B(n_190),
.Y(n_2692)
);

AND2x2_ASAP7_75t_L g2693 ( 
.A(n_2579),
.B(n_190),
.Y(n_2693)
);

INVx2_ASAP7_75t_L g2694 ( 
.A(n_2537),
.Y(n_2694)
);

BUFx3_ASAP7_75t_L g2695 ( 
.A(n_2581),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2583),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2532),
.B(n_191),
.Y(n_2697)
);

AND2x4_ASAP7_75t_SL g2698 ( 
.A(n_2539),
.B(n_191),
.Y(n_2698)
);

OR2x2_ASAP7_75t_L g2699 ( 
.A(n_2544),
.B(n_2562),
.Y(n_2699)
);

OAI221xp5_ASAP7_75t_L g2700 ( 
.A1(n_2624),
.A2(n_195),
.B1(n_192),
.B2(n_193),
.C(n_196),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_L g2701 ( 
.A(n_2522),
.B(n_192),
.Y(n_2701)
);

HB1xp67_ASAP7_75t_L g2702 ( 
.A(n_2586),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2600),
.Y(n_2703)
);

INVx2_ASAP7_75t_L g2704 ( 
.A(n_2609),
.Y(n_2704)
);

INVx2_ASAP7_75t_L g2705 ( 
.A(n_2623),
.Y(n_2705)
);

OAI21xp5_ASAP7_75t_L g2706 ( 
.A1(n_2615),
.A2(n_193),
.B(n_196),
.Y(n_2706)
);

AND2x4_ASAP7_75t_SL g2707 ( 
.A(n_2575),
.B(n_197),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2553),
.Y(n_2708)
);

AOI221xp5_ASAP7_75t_L g2709 ( 
.A1(n_2524),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.C(n_200),
.Y(n_2709)
);

NOR2xp67_ASAP7_75t_L g2710 ( 
.A(n_2571),
.B(n_199),
.Y(n_2710)
);

AND2x2_ASAP7_75t_L g2711 ( 
.A(n_2568),
.B(n_200),
.Y(n_2711)
);

OR2x2_ASAP7_75t_L g2712 ( 
.A(n_2530),
.B(n_201),
.Y(n_2712)
);

NOR2xp33_ASAP7_75t_L g2713 ( 
.A(n_2566),
.B(n_2593),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2545),
.Y(n_2714)
);

AND2x2_ASAP7_75t_L g2715 ( 
.A(n_2516),
.B(n_201),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2515),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2520),
.Y(n_2717)
);

AND2x2_ASAP7_75t_L g2718 ( 
.A(n_2584),
.B(n_203),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2601),
.Y(n_2719)
);

INVx2_ASAP7_75t_L g2720 ( 
.A(n_2619),
.Y(n_2720)
);

AND2x2_ASAP7_75t_L g2721 ( 
.A(n_2606),
.B(n_203),
.Y(n_2721)
);

OR2x2_ASAP7_75t_L g2722 ( 
.A(n_2552),
.B(n_2519),
.Y(n_2722)
);

OR2x2_ASAP7_75t_L g2723 ( 
.A(n_2621),
.B(n_204),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2538),
.B(n_204),
.Y(n_2724)
);

AND2x2_ASAP7_75t_L g2725 ( 
.A(n_2572),
.B(n_205),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2563),
.Y(n_2726)
);

AND2x4_ASAP7_75t_L g2727 ( 
.A(n_2557),
.B(n_206),
.Y(n_2727)
);

AND2x2_ASAP7_75t_L g2728 ( 
.A(n_2618),
.B(n_2509),
.Y(n_2728)
);

AND2x2_ASAP7_75t_L g2729 ( 
.A(n_2585),
.B(n_206),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2589),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2526),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2567),
.B(n_207),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2526),
.Y(n_2733)
);

NOR2xp33_ASAP7_75t_L g2734 ( 
.A(n_2607),
.B(n_207),
.Y(n_2734)
);

INVx2_ASAP7_75t_L g2735 ( 
.A(n_2526),
.Y(n_2735)
);

AND2x4_ASAP7_75t_L g2736 ( 
.A(n_2514),
.B(n_208),
.Y(n_2736)
);

INVx2_ASAP7_75t_L g2737 ( 
.A(n_2526),
.Y(n_2737)
);

AND2x2_ASAP7_75t_L g2738 ( 
.A(n_2512),
.B(n_209),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_2526),
.Y(n_2739)
);

AOI22xp5_ASAP7_75t_L g2740 ( 
.A1(n_2588),
.A2(n_211),
.B1(n_209),
.B2(n_210),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2526),
.Y(n_2741)
);

BUFx2_ASAP7_75t_L g2742 ( 
.A(n_2549),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2526),
.Y(n_2743)
);

OAI221xp5_ASAP7_75t_SL g2744 ( 
.A1(n_2593),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.C(n_213),
.Y(n_2744)
);

AND2x2_ASAP7_75t_L g2745 ( 
.A(n_2512),
.B(n_212),
.Y(n_2745)
);

AND2x4_ASAP7_75t_L g2746 ( 
.A(n_2514),
.B(n_213),
.Y(n_2746)
);

AND2x2_ASAP7_75t_L g2747 ( 
.A(n_2512),
.B(n_214),
.Y(n_2747)
);

INVx2_ASAP7_75t_SL g2748 ( 
.A(n_2565),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2567),
.B(n_214),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2526),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2567),
.B(n_215),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2567),
.B(n_215),
.Y(n_2752)
);

BUFx2_ASAP7_75t_L g2753 ( 
.A(n_2514),
.Y(n_2753)
);

INVx2_ASAP7_75t_L g2754 ( 
.A(n_2526),
.Y(n_2754)
);

HB1xp67_ASAP7_75t_L g2755 ( 
.A(n_2549),
.Y(n_2755)
);

AND2x2_ASAP7_75t_L g2756 ( 
.A(n_2512),
.B(n_216),
.Y(n_2756)
);

INVx2_ASAP7_75t_L g2757 ( 
.A(n_2526),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2526),
.Y(n_2758)
);

HB1xp67_ASAP7_75t_L g2759 ( 
.A(n_2549),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2526),
.Y(n_2760)
);

INVx2_ASAP7_75t_L g2761 ( 
.A(n_2526),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2567),
.B(n_216),
.Y(n_2762)
);

AND2x2_ASAP7_75t_L g2763 ( 
.A(n_2753),
.B(n_217),
.Y(n_2763)
);

AND2x4_ASAP7_75t_L g2764 ( 
.A(n_2748),
.B(n_217),
.Y(n_2764)
);

AND2x2_ASAP7_75t_L g2765 ( 
.A(n_2654),
.B(n_218),
.Y(n_2765)
);

OR2x2_ASAP7_75t_L g2766 ( 
.A(n_2669),
.B(n_218),
.Y(n_2766)
);

OR2x2_ASAP7_75t_L g2767 ( 
.A(n_2670),
.B(n_219),
.Y(n_2767)
);

AND2x4_ASAP7_75t_L g2768 ( 
.A(n_2634),
.B(n_219),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2731),
.Y(n_2769)
);

AND2x2_ASAP7_75t_L g2770 ( 
.A(n_2654),
.B(n_220),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2630),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2733),
.Y(n_2772)
);

OR2x2_ASAP7_75t_L g2773 ( 
.A(n_2625),
.B(n_220),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2741),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2688),
.B(n_2702),
.Y(n_2775)
);

AND2x2_ASAP7_75t_L g2776 ( 
.A(n_2635),
.B(n_221),
.Y(n_2776)
);

AND2x2_ASAP7_75t_L g2777 ( 
.A(n_2681),
.B(n_221),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2742),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2743),
.Y(n_2779)
);

AND2x2_ASAP7_75t_L g2780 ( 
.A(n_2666),
.B(n_222),
.Y(n_2780)
);

INVxp67_ASAP7_75t_L g2781 ( 
.A(n_2686),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_L g2782 ( 
.A(n_2673),
.B(n_222),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2750),
.Y(n_2783)
);

INVxp67_ASAP7_75t_L g2784 ( 
.A(n_2689),
.Y(n_2784)
);

OR2x2_ASAP7_75t_L g2785 ( 
.A(n_2644),
.B(n_223),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2696),
.B(n_223),
.Y(n_2786)
);

AND2x4_ASAP7_75t_L g2787 ( 
.A(n_2683),
.B(n_224),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2760),
.Y(n_2788)
);

AND2x2_ASAP7_75t_L g2789 ( 
.A(n_2638),
.B(n_2668),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2742),
.Y(n_2790)
);

OAI21xp33_ASAP7_75t_L g2791 ( 
.A1(n_2671),
.A2(n_224),
.B(n_225),
.Y(n_2791)
);

AND2x2_ASAP7_75t_L g2792 ( 
.A(n_2637),
.B(n_225),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2703),
.B(n_226),
.Y(n_2793)
);

AND2x2_ASAP7_75t_SL g2794 ( 
.A(n_2690),
.B(n_226),
.Y(n_2794)
);

OR2x2_ASAP7_75t_L g2795 ( 
.A(n_2645),
.B(n_227),
.Y(n_2795)
);

INVx3_ASAP7_75t_L g2796 ( 
.A(n_2736),
.Y(n_2796)
);

INVx1_ASAP7_75t_SL g2797 ( 
.A(n_2664),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2704),
.B(n_227),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2705),
.B(n_228),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2627),
.Y(n_2800)
);

AND2x2_ASAP7_75t_L g2801 ( 
.A(n_2639),
.B(n_229),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2628),
.Y(n_2802)
);

AND2x4_ASAP7_75t_L g2803 ( 
.A(n_2640),
.B(n_2658),
.Y(n_2803)
);

AND2x4_ASAP7_75t_L g2804 ( 
.A(n_2659),
.B(n_229),
.Y(n_2804)
);

NOR2xp67_ASAP7_75t_L g2805 ( 
.A(n_2626),
.B(n_230),
.Y(n_2805)
);

AND2x4_ASAP7_75t_L g2806 ( 
.A(n_2660),
.B(n_230),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_2735),
.Y(n_2807)
);

AND2x2_ASAP7_75t_L g2808 ( 
.A(n_2646),
.B(n_231),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2737),
.Y(n_2809)
);

AND2x2_ASAP7_75t_L g2810 ( 
.A(n_2755),
.B(n_231),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2672),
.B(n_232),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2739),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_L g2813 ( 
.A(n_2677),
.B(n_2662),
.Y(n_2813)
);

AND2x4_ASAP7_75t_L g2814 ( 
.A(n_2649),
.B(n_232),
.Y(n_2814)
);

OR2x2_ASAP7_75t_L g2815 ( 
.A(n_2655),
.B(n_233),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_L g2816 ( 
.A(n_2656),
.B(n_233),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2754),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2757),
.Y(n_2818)
);

OR2x2_ASAP7_75t_L g2819 ( 
.A(n_2657),
.B(n_234),
.Y(n_2819)
);

INVx2_ASAP7_75t_L g2820 ( 
.A(n_2758),
.Y(n_2820)
);

NAND2xp5_ASAP7_75t_SL g2821 ( 
.A(n_2694),
.B(n_234),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2761),
.Y(n_2822)
);

INVx2_ASAP7_75t_L g2823 ( 
.A(n_2759),
.Y(n_2823)
);

INVxp67_ASAP7_75t_SL g2824 ( 
.A(n_2695),
.Y(n_2824)
);

OR2x2_ASAP7_75t_L g2825 ( 
.A(n_2714),
.B(n_2653),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2732),
.Y(n_2826)
);

OR2x2_ASAP7_75t_L g2827 ( 
.A(n_2749),
.B(n_235),
.Y(n_2827)
);

OR2x6_ASAP7_75t_L g2828 ( 
.A(n_2632),
.B(n_235),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2762),
.Y(n_2829)
);

AND2x2_ASAP7_75t_L g2830 ( 
.A(n_2631),
.B(n_236),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2751),
.Y(n_2831)
);

INVx2_ASAP7_75t_L g2832 ( 
.A(n_2684),
.Y(n_2832)
);

OR2x2_ASAP7_75t_L g2833 ( 
.A(n_2752),
.B(n_236),
.Y(n_2833)
);

INVx2_ASAP7_75t_L g2834 ( 
.A(n_2685),
.Y(n_2834)
);

AND2x2_ASAP7_75t_L g2835 ( 
.A(n_2738),
.B(n_237),
.Y(n_2835)
);

INVx2_ASAP7_75t_SL g2836 ( 
.A(n_2746),
.Y(n_2836)
);

NOR2xp33_ASAP7_75t_L g2837 ( 
.A(n_2633),
.B(n_237),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2708),
.Y(n_2838)
);

INVxp67_ASAP7_75t_L g2839 ( 
.A(n_2717),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2650),
.Y(n_2840)
);

INVxp67_ASAP7_75t_SL g2841 ( 
.A(n_2699),
.Y(n_2841)
);

OAI21xp5_ASAP7_75t_L g2842 ( 
.A1(n_2713),
.A2(n_238),
.B(n_239),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_2756),
.Y(n_2843)
);

AOI22xp5_ASAP7_75t_L g2844 ( 
.A1(n_2720),
.A2(n_242),
.B1(n_240),
.B2(n_241),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_2730),
.B(n_2678),
.Y(n_2845)
);

INVx2_ASAP7_75t_L g2846 ( 
.A(n_2747),
.Y(n_2846)
);

NAND2x1_ASAP7_75t_L g2847 ( 
.A(n_2745),
.B(n_241),
.Y(n_2847)
);

AND2x2_ASAP7_75t_L g2848 ( 
.A(n_2647),
.B(n_240),
.Y(n_2848)
);

AND2x2_ASAP7_75t_L g2849 ( 
.A(n_2651),
.B(n_242),
.Y(n_2849)
);

OR2x2_ASAP7_75t_L g2850 ( 
.A(n_2661),
.B(n_2680),
.Y(n_2850)
);

INVx1_ASAP7_75t_SL g2851 ( 
.A(n_2648),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2641),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_2675),
.B(n_243),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2674),
.Y(n_2854)
);

BUFx2_ASAP7_75t_L g2855 ( 
.A(n_2652),
.Y(n_2855)
);

OR2x2_ASAP7_75t_L g2856 ( 
.A(n_2643),
.B(n_243),
.Y(n_2856)
);

INVxp67_ASAP7_75t_L g2857 ( 
.A(n_2667),
.Y(n_2857)
);

AND2x2_ASAP7_75t_L g2858 ( 
.A(n_2679),
.B(n_244),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2676),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2682),
.Y(n_2860)
);

AND2x2_ASAP7_75t_L g2861 ( 
.A(n_2663),
.B(n_244),
.Y(n_2861)
);

AND2x2_ASAP7_75t_SL g2862 ( 
.A(n_2727),
.B(n_245),
.Y(n_2862)
);

AND2x2_ASAP7_75t_L g2863 ( 
.A(n_2734),
.B(n_245),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2665),
.Y(n_2864)
);

NAND2xp5_ASAP7_75t_L g2865 ( 
.A(n_2726),
.B(n_2693),
.Y(n_2865)
);

AND2x2_ASAP7_75t_L g2866 ( 
.A(n_2728),
.B(n_246),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2691),
.Y(n_2867)
);

INVx2_ASAP7_75t_SL g2868 ( 
.A(n_2692),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2697),
.Y(n_2869)
);

AND2x2_ASAP7_75t_L g2870 ( 
.A(n_2716),
.B(n_246),
.Y(n_2870)
);

INVx3_ASAP7_75t_L g2871 ( 
.A(n_2719),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2687),
.Y(n_2872)
);

AND2x2_ASAP7_75t_L g2873 ( 
.A(n_2642),
.B(n_2721),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2723),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2711),
.B(n_2722),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2701),
.Y(n_2876)
);

CKINVDCx16_ASAP7_75t_R g2877 ( 
.A(n_2725),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2712),
.Y(n_2878)
);

OR2x2_ASAP7_75t_L g2879 ( 
.A(n_2715),
.B(n_247),
.Y(n_2879)
);

NAND2x1_ASAP7_75t_SL g2880 ( 
.A(n_2710),
.B(n_247),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2729),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2740),
.B(n_248),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2724),
.Y(n_2883)
);

BUFx2_ASAP7_75t_L g2884 ( 
.A(n_2706),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2629),
.B(n_248),
.Y(n_2885)
);

OR2x2_ASAP7_75t_L g2886 ( 
.A(n_2744),
.B(n_249),
.Y(n_2886)
);

BUFx2_ASAP7_75t_L g2887 ( 
.A(n_2718),
.Y(n_2887)
);

AND2x2_ASAP7_75t_L g2888 ( 
.A(n_2707),
.B(n_249),
.Y(n_2888)
);

NAND2xp67_ASAP7_75t_L g2889 ( 
.A(n_2698),
.B(n_2700),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_2636),
.B(n_250),
.Y(n_2890)
);

INVx2_ASAP7_75t_L g2891 ( 
.A(n_2709),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_L g2892 ( 
.A(n_2669),
.B(n_251),
.Y(n_2892)
);

AND2x2_ASAP7_75t_L g2893 ( 
.A(n_2753),
.B(n_253),
.Y(n_2893)
);

AND2x4_ASAP7_75t_L g2894 ( 
.A(n_2748),
.B(n_253),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2731),
.Y(n_2895)
);

INVx2_ASAP7_75t_L g2896 ( 
.A(n_2753),
.Y(n_2896)
);

AND2x2_ASAP7_75t_L g2897 ( 
.A(n_2753),
.B(n_254),
.Y(n_2897)
);

AND2x2_ASAP7_75t_L g2898 ( 
.A(n_2753),
.B(n_254),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2731),
.Y(n_2899)
);

NOR2xp33_ASAP7_75t_L g2900 ( 
.A(n_2748),
.B(n_255),
.Y(n_2900)
);

AND2x2_ASAP7_75t_L g2901 ( 
.A(n_2753),
.B(n_255),
.Y(n_2901)
);

OR2x2_ASAP7_75t_L g2902 ( 
.A(n_2669),
.B(n_256),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2731),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2731),
.Y(n_2904)
);

INVx1_ASAP7_75t_SL g2905 ( 
.A(n_2664),
.Y(n_2905)
);

OR2x2_ASAP7_75t_L g2906 ( 
.A(n_2669),
.B(n_256),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2731),
.Y(n_2907)
);

AND2x2_ASAP7_75t_L g2908 ( 
.A(n_2753),
.B(n_257),
.Y(n_2908)
);

NOR2xp33_ASAP7_75t_L g2909 ( 
.A(n_2748),
.B(n_257),
.Y(n_2909)
);

INVx2_ASAP7_75t_L g2910 ( 
.A(n_2753),
.Y(n_2910)
);

OR2x2_ASAP7_75t_L g2911 ( 
.A(n_2669),
.B(n_258),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2731),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_L g2913 ( 
.A(n_2669),
.B(n_258),
.Y(n_2913)
);

NOR2x1_ASAP7_75t_L g2914 ( 
.A(n_2695),
.B(n_259),
.Y(n_2914)
);

NOR2xp33_ASAP7_75t_L g2915 ( 
.A(n_2748),
.B(n_259),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2731),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2753),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2731),
.Y(n_2918)
);

INVx2_ASAP7_75t_L g2919 ( 
.A(n_2753),
.Y(n_2919)
);

AND2x4_ASAP7_75t_L g2920 ( 
.A(n_2748),
.B(n_260),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2731),
.Y(n_2921)
);

BUFx2_ASAP7_75t_L g2922 ( 
.A(n_2748),
.Y(n_2922)
);

AND2x2_ASAP7_75t_L g2923 ( 
.A(n_2753),
.B(n_260),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2731),
.Y(n_2924)
);

INVx2_ASAP7_75t_L g2925 ( 
.A(n_2753),
.Y(n_2925)
);

AND2x2_ASAP7_75t_L g2926 ( 
.A(n_2753),
.B(n_261),
.Y(n_2926)
);

OR2x2_ASAP7_75t_L g2927 ( 
.A(n_2669),
.B(n_261),
.Y(n_2927)
);

OR2x2_ASAP7_75t_L g2928 ( 
.A(n_2669),
.B(n_262),
.Y(n_2928)
);

AND2x4_ASAP7_75t_L g2929 ( 
.A(n_2748),
.B(n_262),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_L g2930 ( 
.A(n_2669),
.B(n_263),
.Y(n_2930)
);

AND2x2_ASAP7_75t_L g2931 ( 
.A(n_2753),
.B(n_264),
.Y(n_2931)
);

AND2x2_ASAP7_75t_L g2932 ( 
.A(n_2753),
.B(n_265),
.Y(n_2932)
);

AND2x2_ASAP7_75t_L g2933 ( 
.A(n_2753),
.B(n_265),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2731),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2731),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_2669),
.B(n_266),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2669),
.B(n_266),
.Y(n_2937)
);

AOI21xp33_ASAP7_75t_L g2938 ( 
.A1(n_2713),
.A2(n_267),
.B(n_268),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_L g2939 ( 
.A(n_2669),
.B(n_267),
.Y(n_2939)
);

AND2x2_ASAP7_75t_L g2940 ( 
.A(n_2753),
.B(n_269),
.Y(n_2940)
);

NAND2x1p5_ASAP7_75t_L g2941 ( 
.A(n_2742),
.B(n_269),
.Y(n_2941)
);

INVx2_ASAP7_75t_SL g2942 ( 
.A(n_2634),
.Y(n_2942)
);

INVx2_ASAP7_75t_L g2943 ( 
.A(n_2753),
.Y(n_2943)
);

O2A1O1Ixp33_ASAP7_75t_L g2944 ( 
.A1(n_2642),
.A2(n_273),
.B(n_274),
.C(n_272),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2731),
.Y(n_2945)
);

OR2x2_ASAP7_75t_L g2946 ( 
.A(n_2669),
.B(n_270),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2731),
.Y(n_2947)
);

AND2x2_ASAP7_75t_L g2948 ( 
.A(n_2753),
.B(n_272),
.Y(n_2948)
);

AND2x2_ASAP7_75t_L g2949 ( 
.A(n_2753),
.B(n_275),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2731),
.Y(n_2950)
);

OR2x2_ASAP7_75t_L g2951 ( 
.A(n_2669),
.B(n_275),
.Y(n_2951)
);

INVx2_ASAP7_75t_L g2952 ( 
.A(n_2753),
.Y(n_2952)
);

AND2x4_ASAP7_75t_L g2953 ( 
.A(n_2748),
.B(n_276),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2731),
.Y(n_2954)
);

AND2x2_ASAP7_75t_L g2955 ( 
.A(n_2753),
.B(n_277),
.Y(n_2955)
);

AND2x2_ASAP7_75t_L g2956 ( 
.A(n_2753),
.B(n_277),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2769),
.Y(n_2957)
);

XOR2x2_ASAP7_75t_L g2958 ( 
.A(n_2880),
.B(n_278),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2772),
.Y(n_2959)
);

XOR2x2_ASAP7_75t_L g2960 ( 
.A(n_2862),
.B(n_279),
.Y(n_2960)
);

OR2x2_ASAP7_75t_L g2961 ( 
.A(n_2775),
.B(n_279),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_L g2962 ( 
.A(n_2824),
.B(n_280),
.Y(n_2962)
);

OAI32xp33_ASAP7_75t_L g2963 ( 
.A1(n_2781),
.A2(n_282),
.A3(n_280),
.B1(n_281),
.B2(n_283),
.Y(n_2963)
);

NAND4xp75_ASAP7_75t_L g2964 ( 
.A(n_2914),
.B(n_284),
.C(n_282),
.D(n_283),
.Y(n_2964)
);

AND2x2_ASAP7_75t_L g2965 ( 
.A(n_2922),
.B(n_284),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_2884),
.B(n_285),
.Y(n_2966)
);

OR2x2_ASAP7_75t_L g2967 ( 
.A(n_2825),
.B(n_286),
.Y(n_2967)
);

INVx2_ASAP7_75t_L g2968 ( 
.A(n_2942),
.Y(n_2968)
);

OR2x2_ASAP7_75t_L g2969 ( 
.A(n_2841),
.B(n_2823),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2774),
.Y(n_2970)
);

AOI22xp5_ASAP7_75t_L g2971 ( 
.A1(n_2791),
.A2(n_288),
.B1(n_286),
.B2(n_287),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2779),
.Y(n_2972)
);

INVx2_ASAP7_75t_L g2973 ( 
.A(n_2871),
.Y(n_2973)
);

OR2x2_ASAP7_75t_L g2974 ( 
.A(n_2874),
.B(n_287),
.Y(n_2974)
);

OAI22xp5_ASAP7_75t_L g2975 ( 
.A1(n_2805),
.A2(n_2877),
.B1(n_2784),
.B2(n_2891),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2783),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2788),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2895),
.Y(n_2978)
);

NAND2x1p5_ASAP7_75t_L g2979 ( 
.A(n_2847),
.B(n_289),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_SL g2980 ( 
.A(n_2797),
.B(n_290),
.Y(n_2980)
);

OR2x2_ASAP7_75t_L g2981 ( 
.A(n_2896),
.B(n_291),
.Y(n_2981)
);

AND2x2_ASAP7_75t_L g2982 ( 
.A(n_2905),
.B(n_291),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2899),
.Y(n_2983)
);

XOR2x2_ASAP7_75t_L g2984 ( 
.A(n_2794),
.B(n_292),
.Y(n_2984)
);

AND2x2_ASAP7_75t_L g2985 ( 
.A(n_2789),
.B(n_292),
.Y(n_2985)
);

NOR3xp33_ASAP7_75t_L g2986 ( 
.A(n_2842),
.B(n_294),
.C(n_295),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2910),
.Y(n_2987)
);

XNOR2xp5_ASAP7_75t_L g2988 ( 
.A(n_2851),
.B(n_295),
.Y(n_2988)
);

NAND4xp25_ASAP7_75t_L g2989 ( 
.A(n_2944),
.B(n_298),
.C(n_299),
.D(n_297),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2883),
.B(n_2840),
.Y(n_2990)
);

INVx3_ASAP7_75t_L g2991 ( 
.A(n_2796),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2903),
.Y(n_2992)
);

AND2x2_ASAP7_75t_L g2993 ( 
.A(n_2917),
.B(n_296),
.Y(n_2993)
);

AND2x4_ASAP7_75t_L g2994 ( 
.A(n_2868),
.B(n_296),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_SL g2995 ( 
.A(n_2919),
.B(n_297),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_2925),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2904),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2907),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2912),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2852),
.B(n_298),
.Y(n_3000)
);

NOR2xp67_ASAP7_75t_SL g3001 ( 
.A(n_2889),
.B(n_299),
.Y(n_3001)
);

AND2x2_ASAP7_75t_L g3002 ( 
.A(n_2943),
.B(n_300),
.Y(n_3002)
);

OAI22xp33_ASAP7_75t_L g3003 ( 
.A1(n_2828),
.A2(n_302),
.B1(n_300),
.B2(n_301),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2916),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2918),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2921),
.Y(n_3006)
);

INVx2_ASAP7_75t_SL g3007 ( 
.A(n_2768),
.Y(n_3007)
);

AOI22xp5_ASAP7_75t_L g3008 ( 
.A1(n_2952),
.A2(n_2839),
.B1(n_2873),
.B2(n_2838),
.Y(n_3008)
);

AND2x2_ASAP7_75t_L g3009 ( 
.A(n_2855),
.B(n_302),
.Y(n_3009)
);

INVx2_ASAP7_75t_L g3010 ( 
.A(n_2832),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2924),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2934),
.Y(n_3012)
);

AND2x4_ASAP7_75t_L g3013 ( 
.A(n_2778),
.B(n_303),
.Y(n_3013)
);

INVx3_ASAP7_75t_L g3014 ( 
.A(n_2836),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2935),
.Y(n_3015)
);

OAI32xp33_ASAP7_75t_L g3016 ( 
.A1(n_2886),
.A2(n_306),
.A3(n_304),
.B1(n_305),
.B2(n_307),
.Y(n_3016)
);

AND2x2_ASAP7_75t_L g3017 ( 
.A(n_2878),
.B(n_304),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_L g3018 ( 
.A(n_2872),
.B(n_307),
.Y(n_3018)
);

OAI22xp33_ASAP7_75t_L g3019 ( 
.A1(n_2828),
.A2(n_311),
.B1(n_309),
.B2(n_310),
.Y(n_3019)
);

INVx2_ASAP7_75t_SL g3020 ( 
.A(n_2790),
.Y(n_3020)
);

INVx2_ASAP7_75t_L g3021 ( 
.A(n_2834),
.Y(n_3021)
);

A2O1A1Ixp33_ASAP7_75t_L g3022 ( 
.A1(n_2938),
.A2(n_311),
.B(n_309),
.C(n_310),
.Y(n_3022)
);

AND2x4_ASAP7_75t_L g3023 ( 
.A(n_2771),
.B(n_312),
.Y(n_3023)
);

INVx1_ASAP7_75t_SL g3024 ( 
.A(n_2763),
.Y(n_3024)
);

AOI22xp5_ASAP7_75t_L g3025 ( 
.A1(n_2844),
.A2(n_315),
.B1(n_313),
.B2(n_314),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_L g3026 ( 
.A(n_2854),
.B(n_2859),
.Y(n_3026)
);

OAI32xp33_ASAP7_75t_L g3027 ( 
.A1(n_2941),
.A2(n_316),
.A3(n_313),
.B1(n_315),
.B2(n_317),
.Y(n_3027)
);

AOI22xp5_ASAP7_75t_L g3028 ( 
.A1(n_2867),
.A2(n_320),
.B1(n_317),
.B2(n_318),
.Y(n_3028)
);

BUFx3_ASAP7_75t_L g3029 ( 
.A(n_2764),
.Y(n_3029)
);

NOR2xp33_ASAP7_75t_SL g3030 ( 
.A(n_2893),
.B(n_318),
.Y(n_3030)
);

NAND2x1_ASAP7_75t_L g3031 ( 
.A(n_2807),
.B(n_320),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_2945),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2860),
.B(n_321),
.Y(n_3033)
);

OR2x2_ASAP7_75t_L g3034 ( 
.A(n_2850),
.B(n_321),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2869),
.B(n_322),
.Y(n_3035)
);

AND2x2_ASAP7_75t_L g3036 ( 
.A(n_2864),
.B(n_322),
.Y(n_3036)
);

AND2x2_ASAP7_75t_L g3037 ( 
.A(n_2803),
.B(n_323),
.Y(n_3037)
);

INVxp67_ASAP7_75t_SL g3038 ( 
.A(n_2887),
.Y(n_3038)
);

INVx2_ASAP7_75t_L g3039 ( 
.A(n_2843),
.Y(n_3039)
);

HB1xp67_ASAP7_75t_L g3040 ( 
.A(n_2820),
.Y(n_3040)
);

OR2x2_ASAP7_75t_L g3041 ( 
.A(n_2813),
.B(n_323),
.Y(n_3041)
);

OAI22xp33_ASAP7_75t_L g3042 ( 
.A1(n_2875),
.A2(n_327),
.B1(n_324),
.B2(n_326),
.Y(n_3042)
);

NOR4xp25_ASAP7_75t_L g3043 ( 
.A(n_2821),
.B(n_328),
.C(n_324),
.D(n_327),
.Y(n_3043)
);

AND2x2_ASAP7_75t_L g3044 ( 
.A(n_2826),
.B(n_328),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2947),
.Y(n_3045)
);

NOR2x1_ASAP7_75t_R g3046 ( 
.A(n_2894),
.B(n_329),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2950),
.Y(n_3047)
);

NOR2xp33_ASAP7_75t_L g3048 ( 
.A(n_2857),
.B(n_329),
.Y(n_3048)
);

AOI211x1_ASAP7_75t_L g3049 ( 
.A1(n_2882),
.A2(n_332),
.B(n_330),
.C(n_331),
.Y(n_3049)
);

AND2x2_ASAP7_75t_L g3050 ( 
.A(n_2829),
.B(n_330),
.Y(n_3050)
);

AOI22xp5_ASAP7_75t_L g3051 ( 
.A1(n_2876),
.A2(n_333),
.B1(n_331),
.B2(n_332),
.Y(n_3051)
);

INVxp33_ASAP7_75t_L g3052 ( 
.A(n_2865),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_L g3053 ( 
.A(n_2831),
.B(n_333),
.Y(n_3053)
);

AND2x2_ASAP7_75t_L g3054 ( 
.A(n_2881),
.B(n_334),
.Y(n_3054)
);

OAI22xp5_ASAP7_75t_L g3055 ( 
.A1(n_2845),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_3055)
);

NOR2xp33_ASAP7_75t_L g3056 ( 
.A(n_2786),
.B(n_2793),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2954),
.Y(n_3057)
);

INVx2_ASAP7_75t_L g3058 ( 
.A(n_2846),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2800),
.Y(n_3059)
);

INVxp33_ASAP7_75t_L g3060 ( 
.A(n_2900),
.Y(n_3060)
);

HB1xp67_ASAP7_75t_L g3061 ( 
.A(n_2765),
.Y(n_3061)
);

OA222x2_ASAP7_75t_L g3062 ( 
.A1(n_2766),
.A2(n_339),
.B1(n_341),
.B2(n_335),
.C1(n_337),
.C2(n_340),
.Y(n_3062)
);

INVxp67_ASAP7_75t_L g3063 ( 
.A(n_2770),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2802),
.Y(n_3064)
);

BUFx2_ASAP7_75t_L g3065 ( 
.A(n_2897),
.Y(n_3065)
);

NAND4xp25_ASAP7_75t_L g3066 ( 
.A(n_2885),
.B(n_342),
.C(n_343),
.D(n_340),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2809),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2812),
.Y(n_3068)
);

AND2x2_ASAP7_75t_L g3069 ( 
.A(n_2776),
.B(n_339),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2817),
.Y(n_3070)
);

OR2x6_ASAP7_75t_L g3071 ( 
.A(n_2898),
.B(n_342),
.Y(n_3071)
);

INVx2_ASAP7_75t_L g3072 ( 
.A(n_2818),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2822),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2773),
.Y(n_3074)
);

OR2x2_ASAP7_75t_L g3075 ( 
.A(n_2902),
.B(n_343),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_L g3076 ( 
.A(n_2808),
.B(n_344),
.Y(n_3076)
);

NAND4xp25_ASAP7_75t_L g3077 ( 
.A(n_2909),
.B(n_347),
.C(n_348),
.D(n_345),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2906),
.Y(n_3078)
);

NOR2x1p5_ASAP7_75t_SL g3079 ( 
.A(n_2911),
.B(n_344),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_2901),
.B(n_345),
.Y(n_3080)
);

AOI211xp5_ASAP7_75t_L g3081 ( 
.A1(n_2890),
.A2(n_350),
.B(n_347),
.C(n_349),
.Y(n_3081)
);

NOR2xp67_ASAP7_75t_L g3082 ( 
.A(n_2927),
.B(n_349),
.Y(n_3082)
);

NAND4xp25_ASAP7_75t_SL g3083 ( 
.A(n_2866),
.B(n_352),
.C(n_350),
.D(n_351),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2928),
.Y(n_3084)
);

AOI22xp5_ASAP7_75t_L g3085 ( 
.A1(n_2837),
.A2(n_354),
.B1(n_352),
.B2(n_353),
.Y(n_3085)
);

OR2x2_ASAP7_75t_L g3086 ( 
.A(n_2946),
.B(n_353),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2951),
.Y(n_3087)
);

OAI211xp5_ASAP7_75t_L g3088 ( 
.A1(n_2892),
.A2(n_357),
.B(n_355),
.C(n_356),
.Y(n_3088)
);

NAND4xp25_ASAP7_75t_L g3089 ( 
.A(n_2915),
.B(n_358),
.C(n_359),
.D(n_357),
.Y(n_3089)
);

INVx2_ASAP7_75t_L g3090 ( 
.A(n_2804),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_2815),
.Y(n_3091)
);

INVx2_ASAP7_75t_L g3092 ( 
.A(n_2819),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2785),
.Y(n_3093)
);

INVx1_ASAP7_75t_SL g3094 ( 
.A(n_2908),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2795),
.Y(n_3095)
);

OR2x2_ASAP7_75t_L g3096 ( 
.A(n_2782),
.B(n_356),
.Y(n_3096)
);

AOI33xp33_ASAP7_75t_L g3097 ( 
.A1(n_2861),
.A2(n_360),
.A3(n_362),
.B1(n_358),
.B2(n_359),
.B3(n_361),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_3038),
.Y(n_3098)
);

NAND2xp5_ASAP7_75t_L g3099 ( 
.A(n_3065),
.B(n_2870),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_3024),
.B(n_2777),
.Y(n_3100)
);

AND2x2_ASAP7_75t_L g3101 ( 
.A(n_3014),
.B(n_2923),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_2957),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2959),
.Y(n_3103)
);

AOI21xp33_ASAP7_75t_L g3104 ( 
.A1(n_3052),
.A2(n_2930),
.B(n_2913),
.Y(n_3104)
);

AND2x2_ASAP7_75t_L g3105 ( 
.A(n_2991),
.B(n_2926),
.Y(n_3105)
);

NAND2x1p5_ASAP7_75t_L g3106 ( 
.A(n_3031),
.B(n_3001),
.Y(n_3106)
);

AND2x2_ASAP7_75t_L g3107 ( 
.A(n_3061),
.B(n_2931),
.Y(n_3107)
);

AOI22xp33_ASAP7_75t_L g3108 ( 
.A1(n_2986),
.A2(n_2798),
.B1(n_2799),
.B2(n_2863),
.Y(n_3108)
);

HB1xp67_ASAP7_75t_L g3109 ( 
.A(n_3094),
.Y(n_3109)
);

INVx1_ASAP7_75t_SL g3110 ( 
.A(n_2958),
.Y(n_3110)
);

AND2x2_ASAP7_75t_L g3111 ( 
.A(n_2968),
.B(n_2932),
.Y(n_3111)
);

INVx2_ASAP7_75t_L g3112 ( 
.A(n_3029),
.Y(n_3112)
);

NAND4xp25_ASAP7_75t_SL g3113 ( 
.A(n_3081),
.B(n_2879),
.C(n_2937),
.D(n_2936),
.Y(n_3113)
);

OAI22xp33_ASAP7_75t_L g3114 ( 
.A1(n_2989),
.A2(n_2939),
.B1(n_2767),
.B2(n_2816),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2970),
.Y(n_3115)
);

NOR2xp33_ASAP7_75t_L g3116 ( 
.A(n_3060),
.B(n_2811),
.Y(n_3116)
);

AND2x2_ASAP7_75t_L g3117 ( 
.A(n_2973),
.B(n_2933),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_2972),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_L g3119 ( 
.A(n_3079),
.B(n_2940),
.Y(n_3119)
);

NAND2x1p5_ASAP7_75t_L g3120 ( 
.A(n_2980),
.B(n_2948),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_L g3121 ( 
.A(n_3063),
.B(n_2949),
.Y(n_3121)
);

INVxp67_ASAP7_75t_L g3122 ( 
.A(n_3046),
.Y(n_3122)
);

NAND2x1_ASAP7_75t_L g3123 ( 
.A(n_3020),
.B(n_2955),
.Y(n_3123)
);

HB1xp67_ASAP7_75t_L g3124 ( 
.A(n_2969),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_2976),
.Y(n_3125)
);

AND2x2_ASAP7_75t_L g3126 ( 
.A(n_3092),
.B(n_2956),
.Y(n_3126)
);

INVxp67_ASAP7_75t_L g3127 ( 
.A(n_3030),
.Y(n_3127)
);

INVx1_ASAP7_75t_SL g3128 ( 
.A(n_2965),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_2977),
.Y(n_3129)
);

OR2x2_ASAP7_75t_L g3130 ( 
.A(n_3078),
.B(n_2827),
.Y(n_3130)
);

OR2x2_ASAP7_75t_L g3131 ( 
.A(n_3084),
.B(n_2833),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2978),
.Y(n_3132)
);

NOR2xp33_ASAP7_75t_L g3133 ( 
.A(n_3007),
.B(n_2856),
.Y(n_3133)
);

INVx2_ASAP7_75t_L g3134 ( 
.A(n_3090),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_L g3135 ( 
.A(n_3056),
.B(n_2780),
.Y(n_3135)
);

AND2x2_ASAP7_75t_L g3136 ( 
.A(n_3074),
.B(n_3087),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2983),
.Y(n_3137)
);

OAI21xp33_ASAP7_75t_L g3138 ( 
.A1(n_3008),
.A2(n_2853),
.B(n_2801),
.Y(n_3138)
);

INVx1_ASAP7_75t_SL g3139 ( 
.A(n_2960),
.Y(n_3139)
);

INVx2_ASAP7_75t_L g3140 ( 
.A(n_3013),
.Y(n_3140)
);

AOI22xp5_ASAP7_75t_L g3141 ( 
.A1(n_2975),
.A2(n_2929),
.B1(n_2953),
.B2(n_2920),
.Y(n_3141)
);

INVx2_ASAP7_75t_L g3142 ( 
.A(n_3013),
.Y(n_3142)
);

BUFx2_ASAP7_75t_L g3143 ( 
.A(n_2979),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_L g3144 ( 
.A(n_3091),
.B(n_2814),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2992),
.Y(n_3145)
);

AND2x2_ASAP7_75t_SL g3146 ( 
.A(n_3043),
.B(n_2787),
.Y(n_3146)
);

AND2x2_ASAP7_75t_L g3147 ( 
.A(n_3093),
.B(n_2792),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_L g3148 ( 
.A(n_3095),
.B(n_3082),
.Y(n_3148)
);

INVx2_ASAP7_75t_L g3149 ( 
.A(n_3023),
.Y(n_3149)
);

OR2x2_ASAP7_75t_L g3150 ( 
.A(n_2987),
.B(n_2810),
.Y(n_3150)
);

INVx2_ASAP7_75t_SL g3151 ( 
.A(n_2994),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_2997),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2998),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_2999),
.Y(n_3154)
);

HB1xp67_ASAP7_75t_L g3155 ( 
.A(n_3040),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_3004),
.Y(n_3156)
);

NAND2x1p5_ASAP7_75t_L g3157 ( 
.A(n_2995),
.B(n_2806),
.Y(n_3157)
);

INVx1_ASAP7_75t_SL g3158 ( 
.A(n_2984),
.Y(n_3158)
);

AND2x2_ASAP7_75t_L g3159 ( 
.A(n_2996),
.B(n_2858),
.Y(n_3159)
);

AOI21xp33_ASAP7_75t_L g3160 ( 
.A1(n_2990),
.A2(n_2888),
.B(n_2849),
.Y(n_3160)
);

NOR2xp33_ASAP7_75t_L g3161 ( 
.A(n_3034),
.B(n_2848),
.Y(n_3161)
);

INVx2_ASAP7_75t_L g3162 ( 
.A(n_3023),
.Y(n_3162)
);

AND2x2_ASAP7_75t_L g3163 ( 
.A(n_3039),
.B(n_3058),
.Y(n_3163)
);

INVx2_ASAP7_75t_L g3164 ( 
.A(n_2981),
.Y(n_3164)
);

AND2x2_ASAP7_75t_L g3165 ( 
.A(n_2985),
.B(n_2830),
.Y(n_3165)
);

AND2x2_ASAP7_75t_L g3166 ( 
.A(n_3054),
.B(n_2835),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_L g3167 ( 
.A(n_2966),
.B(n_362),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_3005),
.Y(n_3168)
);

NAND2x1_ASAP7_75t_L g3169 ( 
.A(n_3010),
.B(n_363),
.Y(n_3169)
);

OR2x2_ASAP7_75t_L g3170 ( 
.A(n_2967),
.B(n_363),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_3006),
.Y(n_3171)
);

OR2x2_ASAP7_75t_L g3172 ( 
.A(n_2961),
.B(n_364),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_L g3173 ( 
.A(n_3036),
.B(n_3044),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_3011),
.Y(n_3174)
);

NAND2xp33_ASAP7_75t_L g3175 ( 
.A(n_2964),
.B(n_364),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_3012),
.Y(n_3176)
);

AND2x4_ASAP7_75t_L g3177 ( 
.A(n_3021),
.B(n_365),
.Y(n_3177)
);

AND2x2_ASAP7_75t_L g3178 ( 
.A(n_2982),
.B(n_366),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_3155),
.Y(n_3179)
);

NOR2xp33_ASAP7_75t_L g3180 ( 
.A(n_3139),
.B(n_3158),
.Y(n_3180)
);

OAI21xp5_ASAP7_75t_L g3181 ( 
.A1(n_3175),
.A2(n_3022),
.B(n_3055),
.Y(n_3181)
);

OR2x2_ASAP7_75t_L g3182 ( 
.A(n_3128),
.B(n_3026),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_3109),
.Y(n_3183)
);

OR2x2_ASAP7_75t_L g3184 ( 
.A(n_3148),
.B(n_3098),
.Y(n_3184)
);

AOI221xp5_ASAP7_75t_L g3185 ( 
.A1(n_3110),
.A2(n_3042),
.B1(n_3104),
.B2(n_3124),
.C(n_3049),
.Y(n_3185)
);

OA21x2_ASAP7_75t_L g3186 ( 
.A1(n_3127),
.A2(n_2962),
.B(n_3000),
.Y(n_3186)
);

AOI221xp5_ASAP7_75t_L g3187 ( 
.A1(n_3114),
.A2(n_3016),
.B1(n_3003),
.B2(n_3019),
.C(n_2963),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_3146),
.B(n_3050),
.Y(n_3188)
);

AND2x2_ASAP7_75t_L g3189 ( 
.A(n_3101),
.B(n_3071),
.Y(n_3189)
);

OAI211xp5_ASAP7_75t_L g3190 ( 
.A1(n_3122),
.A2(n_3088),
.B(n_3025),
.C(n_2971),
.Y(n_3190)
);

AND2x2_ASAP7_75t_L g3191 ( 
.A(n_3105),
.B(n_3071),
.Y(n_3191)
);

INVx2_ASAP7_75t_L g3192 ( 
.A(n_3143),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_3136),
.Y(n_3193)
);

XNOR2xp5_ASAP7_75t_L g3194 ( 
.A(n_3141),
.B(n_2988),
.Y(n_3194)
);

INVx2_ASAP7_75t_L g3195 ( 
.A(n_3106),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_3130),
.Y(n_3196)
);

OAI21xp33_ASAP7_75t_L g3197 ( 
.A1(n_3134),
.A2(n_3099),
.B(n_3112),
.Y(n_3197)
);

NOR2xp33_ASAP7_75t_L g3198 ( 
.A(n_3119),
.B(n_3041),
.Y(n_3198)
);

OR2x2_ASAP7_75t_L g3199 ( 
.A(n_3140),
.B(n_3072),
.Y(n_3199)
);

INVx2_ASAP7_75t_L g3200 ( 
.A(n_3151),
.Y(n_3200)
);

OAI221xp5_ASAP7_75t_L g3201 ( 
.A1(n_3123),
.A2(n_3085),
.B1(n_3066),
.B2(n_3089),
.C(n_3077),
.Y(n_3201)
);

AOI21xp33_ASAP7_75t_L g3202 ( 
.A1(n_3131),
.A2(n_3064),
.B(n_3059),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_3107),
.B(n_3009),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_3165),
.B(n_3017),
.Y(n_3204)
);

A2O1A1Ixp33_ASAP7_75t_L g3205 ( 
.A1(n_3169),
.A2(n_3097),
.B(n_3028),
.C(n_3051),
.Y(n_3205)
);

OAI222xp33_ASAP7_75t_L g3206 ( 
.A1(n_3120),
.A2(n_2974),
.B1(n_3035),
.B2(n_3067),
.C1(n_3070),
.C2(n_3068),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_SL g3207 ( 
.A(n_3142),
.B(n_3048),
.Y(n_3207)
);

AND2x2_ASAP7_75t_L g3208 ( 
.A(n_3111),
.B(n_2993),
.Y(n_3208)
);

AOI21xp33_ASAP7_75t_L g3209 ( 
.A1(n_3164),
.A2(n_3073),
.B(n_3032),
.Y(n_3209)
);

AND2x2_ASAP7_75t_L g3210 ( 
.A(n_3117),
.B(n_3002),
.Y(n_3210)
);

AND2x2_ASAP7_75t_L g3211 ( 
.A(n_3126),
.B(n_3037),
.Y(n_3211)
);

OAI22xp5_ASAP7_75t_L g3212 ( 
.A1(n_3108),
.A2(n_3018),
.B1(n_3033),
.B2(n_3053),
.Y(n_3212)
);

AOI221xp5_ASAP7_75t_L g3213 ( 
.A1(n_3138),
.A2(n_3083),
.B1(n_3027),
.B2(n_3045),
.C(n_3047),
.Y(n_3213)
);

INVxp67_ASAP7_75t_L g3214 ( 
.A(n_3161),
.Y(n_3214)
);

XOR2x2_ASAP7_75t_L g3215 ( 
.A(n_3157),
.B(n_3080),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_L g3216 ( 
.A(n_3166),
.B(n_3015),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_3147),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_3149),
.B(n_3162),
.Y(n_3218)
);

OAI21xp5_ASAP7_75t_SL g3219 ( 
.A1(n_3116),
.A2(n_3069),
.B(n_3096),
.Y(n_3219)
);

AOI22xp5_ASAP7_75t_L g3220 ( 
.A1(n_3133),
.A2(n_3113),
.B1(n_3159),
.B2(n_3121),
.Y(n_3220)
);

NAND2xp33_ASAP7_75t_L g3221 ( 
.A(n_3173),
.B(n_3062),
.Y(n_3221)
);

OAI221xp5_ASAP7_75t_L g3222 ( 
.A1(n_3100),
.A2(n_3057),
.B1(n_3076),
.B2(n_3086),
.C(n_3075),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_3163),
.B(n_366),
.Y(n_3223)
);

AOI21xp5_ASAP7_75t_L g3224 ( 
.A1(n_3135),
.A2(n_367),
.B(n_368),
.Y(n_3224)
);

OAI322xp33_ASAP7_75t_L g3225 ( 
.A1(n_3102),
.A2(n_374),
.A3(n_373),
.B1(n_371),
.B2(n_369),
.C1(n_370),
.C2(n_372),
.Y(n_3225)
);

AOI21xp33_ASAP7_75t_SL g3226 ( 
.A1(n_3150),
.A2(n_3160),
.B(n_3144),
.Y(n_3226)
);

OR2x2_ASAP7_75t_L g3227 ( 
.A(n_3172),
.B(n_369),
.Y(n_3227)
);

NAND2xp5_ASAP7_75t_L g3228 ( 
.A(n_3177),
.B(n_370),
.Y(n_3228)
);

AOI221xp5_ASAP7_75t_SL g3229 ( 
.A1(n_3103),
.A2(n_373),
.B1(n_371),
.B2(n_372),
.C(n_375),
.Y(n_3229)
);

INVx1_ASAP7_75t_SL g3230 ( 
.A(n_3178),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_3115),
.Y(n_3231)
);

NOR2x1p5_ASAP7_75t_L g3232 ( 
.A(n_3167),
.B(n_375),
.Y(n_3232)
);

INVx2_ASAP7_75t_L g3233 ( 
.A(n_3177),
.Y(n_3233)
);

AOI21xp5_ASAP7_75t_L g3234 ( 
.A1(n_3170),
.A2(n_3125),
.B(n_3118),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_3129),
.Y(n_3235)
);

AOI21xp33_ASAP7_75t_SL g3236 ( 
.A1(n_3132),
.A2(n_376),
.B(n_378),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_3137),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_3145),
.B(n_378),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_3183),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_3218),
.Y(n_3240)
);

OAI322xp33_ASAP7_75t_L g3241 ( 
.A1(n_3188),
.A2(n_3180),
.A3(n_3179),
.B1(n_3184),
.B2(n_3220),
.C1(n_3201),
.C2(n_3198),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_3227),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_3193),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_3217),
.Y(n_3244)
);

OAI21xp33_ASAP7_75t_SL g3245 ( 
.A1(n_3185),
.A2(n_3153),
.B(n_3152),
.Y(n_3245)
);

OR2x2_ASAP7_75t_L g3246 ( 
.A(n_3203),
.B(n_3154),
.Y(n_3246)
);

OAI22xp33_ASAP7_75t_L g3247 ( 
.A1(n_3181),
.A2(n_3168),
.B1(n_3171),
.B2(n_3156),
.Y(n_3247)
);

OAI21xp5_ASAP7_75t_L g3248 ( 
.A1(n_3221),
.A2(n_3205),
.B(n_3224),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_SL g3249 ( 
.A(n_3187),
.B(n_3174),
.Y(n_3249)
);

AOI21xp33_ASAP7_75t_SL g3250 ( 
.A1(n_3194),
.A2(n_3176),
.B(n_379),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_3230),
.B(n_380),
.Y(n_3251)
);

OAI21xp33_ASAP7_75t_L g3252 ( 
.A1(n_3197),
.A2(n_380),
.B(n_381),
.Y(n_3252)
);

XOR2x2_ASAP7_75t_L g3253 ( 
.A(n_3215),
.B(n_381),
.Y(n_3253)
);

AOI21xp33_ASAP7_75t_L g3254 ( 
.A1(n_3195),
.A2(n_382),
.B(n_383),
.Y(n_3254)
);

INVxp67_ASAP7_75t_L g3255 ( 
.A(n_3189),
.Y(n_3255)
);

OAI21xp5_ASAP7_75t_L g3256 ( 
.A1(n_3190),
.A2(n_382),
.B(n_384),
.Y(n_3256)
);

INVx1_ASAP7_75t_SL g3257 ( 
.A(n_3191),
.Y(n_3257)
);

OAI211xp5_ASAP7_75t_SL g3258 ( 
.A1(n_3214),
.A2(n_387),
.B(n_385),
.C(n_386),
.Y(n_3258)
);

OAI221xp5_ASAP7_75t_L g3259 ( 
.A1(n_3213),
.A2(n_389),
.B1(n_387),
.B2(n_388),
.C(n_390),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_3196),
.Y(n_3260)
);

OAI32xp33_ASAP7_75t_L g3261 ( 
.A1(n_3182),
.A2(n_390),
.A3(n_388),
.B1(n_389),
.B2(n_391),
.Y(n_3261)
);

AND2x2_ASAP7_75t_L g3262 ( 
.A(n_3208),
.B(n_391),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_3210),
.B(n_393),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_L g3264 ( 
.A(n_3200),
.B(n_393),
.Y(n_3264)
);

AND2x2_ASAP7_75t_L g3265 ( 
.A(n_3211),
.B(n_394),
.Y(n_3265)
);

NOR2xp33_ASAP7_75t_R g3266 ( 
.A(n_3192),
.B(n_394),
.Y(n_3266)
);

OAI21xp33_ASAP7_75t_SL g3267 ( 
.A1(n_3202),
.A2(n_3207),
.B(n_3209),
.Y(n_3267)
);

NAND4xp25_ASAP7_75t_L g3268 ( 
.A(n_3226),
.B(n_397),
.C(n_395),
.D(n_396),
.Y(n_3268)
);

INVx2_ASAP7_75t_SL g3269 ( 
.A(n_3233),
.Y(n_3269)
);

NOR2xp33_ASAP7_75t_L g3270 ( 
.A(n_3219),
.B(n_3222),
.Y(n_3270)
);

AOI31xp33_ASAP7_75t_L g3271 ( 
.A1(n_3229),
.A2(n_3236),
.A3(n_3199),
.B(n_3234),
.Y(n_3271)
);

XOR2x2_ASAP7_75t_L g3272 ( 
.A(n_3204),
.B(n_397),
.Y(n_3272)
);

AOI221xp5_ASAP7_75t_L g3273 ( 
.A1(n_3206),
.A2(n_400),
.B1(n_398),
.B2(n_399),
.C(n_401),
.Y(n_3273)
);

NAND2xp5_ASAP7_75t_L g3274 ( 
.A(n_3232),
.B(n_398),
.Y(n_3274)
);

OAI322xp33_ASAP7_75t_L g3275 ( 
.A1(n_3231),
.A2(n_406),
.A3(n_405),
.B1(n_403),
.B2(n_399),
.C1(n_402),
.C2(n_404),
.Y(n_3275)
);

OAI22xp5_ASAP7_75t_L g3276 ( 
.A1(n_3212),
.A2(n_405),
.B1(n_403),
.B2(n_404),
.Y(n_3276)
);

NAND5xp2_ASAP7_75t_L g3277 ( 
.A(n_3270),
.B(n_3216),
.C(n_3237),
.D(n_3235),
.E(n_3223),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_3269),
.Y(n_3278)
);

AOI21xp5_ASAP7_75t_L g3279 ( 
.A1(n_3248),
.A2(n_3186),
.B(n_3238),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_3262),
.Y(n_3280)
);

AND2x2_ASAP7_75t_L g3281 ( 
.A(n_3257),
.B(n_3186),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_3265),
.Y(n_3282)
);

NAND3xp33_ASAP7_75t_L g3283 ( 
.A(n_3273),
.B(n_3228),
.C(n_3225),
.Y(n_3283)
);

AOI21xp5_ASAP7_75t_L g3284 ( 
.A1(n_3241),
.A2(n_3249),
.B(n_3256),
.Y(n_3284)
);

AOI22xp5_ASAP7_75t_L g3285 ( 
.A1(n_3259),
.A2(n_409),
.B1(n_407),
.B2(n_408),
.Y(n_3285)
);

AOI22xp5_ASAP7_75t_L g3286 ( 
.A1(n_3267),
.A2(n_411),
.B1(n_408),
.B2(n_410),
.Y(n_3286)
);

AOI211xp5_ASAP7_75t_L g3287 ( 
.A1(n_3245),
.A2(n_413),
.B(n_410),
.C(n_412),
.Y(n_3287)
);

AOI211xp5_ASAP7_75t_L g3288 ( 
.A1(n_3247),
.A2(n_415),
.B(n_413),
.C(n_414),
.Y(n_3288)
);

INVxp67_ASAP7_75t_L g3289 ( 
.A(n_3274),
.Y(n_3289)
);

OAI32xp33_ASAP7_75t_L g3290 ( 
.A1(n_3268),
.A2(n_416),
.A3(n_414),
.B1(n_415),
.B2(n_417),
.Y(n_3290)
);

AOI22xp33_ASAP7_75t_L g3291 ( 
.A1(n_3253),
.A2(n_420),
.B1(n_418),
.B2(n_419),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_3264),
.Y(n_3292)
);

O2A1O1Ixp33_ASAP7_75t_L g3293 ( 
.A1(n_3271),
.A2(n_421),
.B(n_418),
.C(n_420),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_3242),
.Y(n_3294)
);

OAI21xp33_ASAP7_75t_L g3295 ( 
.A1(n_3255),
.A2(n_421),
.B(n_422),
.Y(n_3295)
);

AOI221xp5_ASAP7_75t_L g3296 ( 
.A1(n_3250),
.A2(n_3239),
.B1(n_3260),
.B2(n_3275),
.C(n_3261),
.Y(n_3296)
);

AOI221xp5_ASAP7_75t_L g3297 ( 
.A1(n_3276),
.A2(n_424),
.B1(n_422),
.B2(n_423),
.C(n_425),
.Y(n_3297)
);

AOI22xp5_ASAP7_75t_L g3298 ( 
.A1(n_3272),
.A2(n_426),
.B1(n_424),
.B2(n_425),
.Y(n_3298)
);

AOI221xp5_ASAP7_75t_L g3299 ( 
.A1(n_3244),
.A2(n_428),
.B1(n_426),
.B2(n_427),
.C(n_429),
.Y(n_3299)
);

AOI322xp5_ASAP7_75t_L g3300 ( 
.A1(n_3252),
.A2(n_433),
.A3(n_432),
.B1(n_430),
.B2(n_427),
.C1(n_428),
.C2(n_431),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_3263),
.Y(n_3301)
);

O2A1O1Ixp33_ASAP7_75t_SL g3302 ( 
.A1(n_3254),
.A2(n_435),
.B(n_432),
.C(n_433),
.Y(n_3302)
);

OAI221xp5_ASAP7_75t_SL g3303 ( 
.A1(n_3246),
.A2(n_437),
.B1(n_435),
.B2(n_436),
.C(n_438),
.Y(n_3303)
);

AOI222xp33_ASAP7_75t_L g3304 ( 
.A1(n_3240),
.A2(n_439),
.B1(n_441),
.B2(n_436),
.C1(n_438),
.C2(n_440),
.Y(n_3304)
);

AND2x2_ASAP7_75t_L g3305 ( 
.A(n_3266),
.B(n_440),
.Y(n_3305)
);

HB1xp67_ASAP7_75t_L g3306 ( 
.A(n_3251),
.Y(n_3306)
);

A2O1A1Ixp33_ASAP7_75t_L g3307 ( 
.A1(n_3258),
.A2(n_443),
.B(n_441),
.C(n_442),
.Y(n_3307)
);

AOI322xp5_ASAP7_75t_L g3308 ( 
.A1(n_3243),
.A2(n_449),
.A3(n_448),
.B1(n_446),
.B2(n_443),
.C1(n_444),
.C2(n_447),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_3269),
.B(n_444),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_3269),
.Y(n_3310)
);

AND2x2_ASAP7_75t_L g3311 ( 
.A(n_3257),
.B(n_446),
.Y(n_3311)
);

AOI22xp5_ASAP7_75t_L g3312 ( 
.A1(n_3249),
.A2(n_450),
.B1(n_448),
.B2(n_449),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_3269),
.Y(n_3313)
);

INVx1_ASAP7_75t_SL g3314 ( 
.A(n_3281),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_SL g3315 ( 
.A(n_3284),
.B(n_450),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_3311),
.B(n_451),
.Y(n_3316)
);

AOI211xp5_ASAP7_75t_L g3317 ( 
.A1(n_3293),
.A2(n_453),
.B(n_451),
.C(n_452),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_L g3318 ( 
.A(n_3278),
.B(n_452),
.Y(n_3318)
);

AOI22xp5_ASAP7_75t_L g3319 ( 
.A1(n_3312),
.A2(n_455),
.B1(n_549),
.B2(n_547),
.Y(n_3319)
);

OA22x2_ASAP7_75t_L g3320 ( 
.A1(n_3286),
.A2(n_455),
.B1(n_551),
.B2(n_550),
.Y(n_3320)
);

AOI21xp5_ASAP7_75t_L g3321 ( 
.A1(n_3279),
.A2(n_552),
.B(n_553),
.Y(n_3321)
);

OAI22xp5_ASAP7_75t_L g3322 ( 
.A1(n_3291),
.A2(n_557),
.B1(n_555),
.B2(n_556),
.Y(n_3322)
);

OA22x2_ASAP7_75t_L g3323 ( 
.A1(n_3310),
.A2(n_562),
.B1(n_558),
.B2(n_560),
.Y(n_3323)
);

AOI211x1_ASAP7_75t_SL g3324 ( 
.A1(n_3283),
.A2(n_567),
.B(n_564),
.C(n_566),
.Y(n_3324)
);

AOI21xp5_ASAP7_75t_L g3325 ( 
.A1(n_3287),
.A2(n_568),
.B(n_569),
.Y(n_3325)
);

NOR2x1_ASAP7_75t_L g3326 ( 
.A(n_3313),
.B(n_570),
.Y(n_3326)
);

NOR2xp33_ASAP7_75t_L g3327 ( 
.A(n_3280),
.B(n_865),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_3282),
.B(n_571),
.Y(n_3328)
);

NAND2x1_ASAP7_75t_SL g3329 ( 
.A(n_3305),
.B(n_573),
.Y(n_3329)
);

AOI211x1_ASAP7_75t_L g3330 ( 
.A1(n_3290),
.A2(n_577),
.B(n_574),
.C(n_576),
.Y(n_3330)
);

AND3x2_ASAP7_75t_L g3331 ( 
.A(n_3288),
.B(n_578),
.C(n_579),
.Y(n_3331)
);

AOI211x1_ASAP7_75t_L g3332 ( 
.A1(n_3294),
.A2(n_3309),
.B(n_3295),
.C(n_3301),
.Y(n_3332)
);

INVx1_ASAP7_75t_L g3333 ( 
.A(n_3306),
.Y(n_3333)
);

NOR3xp33_ASAP7_75t_L g3334 ( 
.A(n_3277),
.B(n_3289),
.C(n_3296),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_3292),
.Y(n_3335)
);

AND2x2_ASAP7_75t_L g3336 ( 
.A(n_3298),
.B(n_584),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_L g3337 ( 
.A(n_3304),
.B(n_585),
.Y(n_3337)
);

AOI22xp5_ASAP7_75t_L g3338 ( 
.A1(n_3334),
.A2(n_3285),
.B1(n_3297),
.B2(n_3299),
.Y(n_3338)
);

NOR4xp25_ASAP7_75t_L g3339 ( 
.A(n_3315),
.B(n_3303),
.C(n_3302),
.D(n_3307),
.Y(n_3339)
);

AOI221xp5_ASAP7_75t_L g3340 ( 
.A1(n_3314),
.A2(n_3308),
.B1(n_3300),
.B2(n_592),
.C(n_588),
.Y(n_3340)
);

NOR2xp33_ASAP7_75t_L g3341 ( 
.A(n_3329),
.B(n_591),
.Y(n_3341)
);

NOR2x1_ASAP7_75t_L g3342 ( 
.A(n_3326),
.B(n_594),
.Y(n_3342)
);

OAI21xp33_ASAP7_75t_L g3343 ( 
.A1(n_3333),
.A2(n_595),
.B(n_596),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_L g3344 ( 
.A(n_3317),
.B(n_599),
.Y(n_3344)
);

AND4x1_ASAP7_75t_L g3345 ( 
.A(n_3324),
.B(n_604),
.C(n_601),
.D(n_603),
.Y(n_3345)
);

O2A1O1Ixp33_ASAP7_75t_SL g3346 ( 
.A1(n_3316),
.A2(n_864),
.B(n_607),
.C(n_605),
.Y(n_3346)
);

NOR2xp67_ASAP7_75t_L g3347 ( 
.A(n_3318),
.B(n_606),
.Y(n_3347)
);

A2O1A1Ixp33_ASAP7_75t_L g3348 ( 
.A1(n_3321),
.A2(n_612),
.B(n_609),
.C(n_611),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_3330),
.B(n_614),
.Y(n_3349)
);

OR2x2_ASAP7_75t_L g3350 ( 
.A(n_3339),
.B(n_3337),
.Y(n_3350)
);

NOR3xp33_ASAP7_75t_L g3351 ( 
.A(n_3340),
.B(n_3335),
.C(n_3328),
.Y(n_3351)
);

INVxp33_ASAP7_75t_L g3352 ( 
.A(n_3342),
.Y(n_3352)
);

INVx2_ASAP7_75t_L g3353 ( 
.A(n_3344),
.Y(n_3353)
);

NOR3xp33_ASAP7_75t_L g3354 ( 
.A(n_3338),
.B(n_3327),
.C(n_3322),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_3350),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_3353),
.Y(n_3356)
);

AND4x1_ASAP7_75t_L g3357 ( 
.A(n_3355),
.B(n_3351),
.C(n_3354),
.D(n_3341),
.Y(n_3357)
);

AOI21xp33_ASAP7_75t_L g3358 ( 
.A1(n_3356),
.A2(n_3352),
.B(n_3320),
.Y(n_3358)
);

INVxp67_ASAP7_75t_SL g3359 ( 
.A(n_3357),
.Y(n_3359)
);

INVx1_ASAP7_75t_SL g3360 ( 
.A(n_3358),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_3357),
.B(n_3332),
.Y(n_3361)
);

CKINVDCx5p33_ASAP7_75t_R g3362 ( 
.A(n_3360),
.Y(n_3362)
);

OAI222xp33_ASAP7_75t_L g3363 ( 
.A1(n_3361),
.A2(n_3325),
.B1(n_3349),
.B2(n_3323),
.C1(n_3319),
.C2(n_3336),
.Y(n_3363)
);

INVx2_ASAP7_75t_L g3364 ( 
.A(n_3359),
.Y(n_3364)
);

OAI221xp5_ASAP7_75t_L g3365 ( 
.A1(n_3362),
.A2(n_3347),
.B1(n_3343),
.B2(n_3348),
.C(n_3345),
.Y(n_3365)
);

NOR3xp33_ASAP7_75t_SL g3366 ( 
.A(n_3363),
.B(n_3346),
.C(n_3331),
.Y(n_3366)
);

INVxp67_ASAP7_75t_SL g3367 ( 
.A(n_3365),
.Y(n_3367)
);

NOR3xp33_ASAP7_75t_L g3368 ( 
.A(n_3367),
.B(n_3364),
.C(n_3366),
.Y(n_3368)
);

OAI22xp5_ASAP7_75t_SL g3369 ( 
.A1(n_3368),
.A2(n_619),
.B1(n_616),
.B2(n_617),
.Y(n_3369)
);

INVx3_ASAP7_75t_L g3370 ( 
.A(n_3369),
.Y(n_3370)
);

AOI21xp5_ASAP7_75t_L g3371 ( 
.A1(n_3370),
.A2(n_620),
.B(n_621),
.Y(n_3371)
);

AOI322xp5_ASAP7_75t_L g3372 ( 
.A1(n_3371),
.A2(n_637),
.A3(n_633),
.B1(n_629),
.B2(n_622),
.C1(n_625),
.C2(n_631),
.Y(n_3372)
);

AOI22xp5_ASAP7_75t_L g3373 ( 
.A1(n_3372),
.A2(n_640),
.B1(n_638),
.B2(n_639),
.Y(n_3373)
);

AOI31xp33_ASAP7_75t_L g3374 ( 
.A1(n_3373),
.A2(n_644),
.A3(n_642),
.B(n_643),
.Y(n_3374)
);


endmodule