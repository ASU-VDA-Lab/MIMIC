module fake_jpeg_14238_n_138 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_138);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_138;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx3_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_38),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_40),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_15),
.B(n_29),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_0),
.B(n_10),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_5),
.B(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_9),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_12),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_60),
.A2(n_52),
.B1(n_44),
.B2(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_1),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_61),
.B(n_65),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_63),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_3),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_67),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx5_ASAP7_75t_SL g68 ( 
.A(n_48),
.Y(n_68)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_69),
.A2(n_23),
.B(n_37),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_53),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_56),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_62),
.A2(n_42),
.B1(n_44),
.B2(n_54),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_74),
.A2(n_50),
.B1(n_55),
.B2(n_46),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_43),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_82),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_58),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_72),
.B(n_25),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_95),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_86),
.B(n_89),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_78),
.A2(n_72),
.B1(n_74),
.B2(n_76),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_88),
.B(n_39),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_78),
.A2(n_45),
.B1(n_4),
.B2(n_5),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_75),
.C(n_79),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_26),
.C(n_36),
.Y(n_102)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

FAx1_ASAP7_75t_SL g93 ( 
.A(n_79),
.B(n_3),
.CI(n_6),
.CON(n_93),
.SN(n_93)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_94),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_98),
.Y(n_104)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_100),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_114),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_8),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_106),
.B(n_107),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_10),
.Y(n_107)
);

MAJx2_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_11),
.C(n_13),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_108),
.A2(n_84),
.B(n_33),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_14),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_110),
.B(n_111),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_18),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_86),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_27),
.C(n_30),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_34),
.Y(n_125)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_121),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_104),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_108),
.C(n_102),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_103),
.B(n_32),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_125),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_122),
.A2(n_109),
.B(n_112),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_127),
.A2(n_120),
.B1(n_105),
.B2(n_113),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_128),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_132),
.B(n_129),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_117),
.C(n_112),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_131),
.C(n_118),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_135),
.B(n_131),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

AOI221xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_120),
.B1(n_115),
.B2(n_35),
.C(n_114),
.Y(n_138)
);


endmodule