module fake_jpeg_8546_n_59 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_59);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_59;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_38;
wire n_36;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx2_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_6),
.B(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_11),
.B(n_15),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_25),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_23),
.B(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_30),
.B(n_35),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_41),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_0),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_29),
.A2(n_12),
.B1(n_2),
.B2(n_3),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_44),
.Y(n_49)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_29),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_1),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_31),
.B(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_50),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_49),
.A2(n_42),
.B1(n_34),
.B2(n_8),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_52),
.B(n_47),
.Y(n_54)
);

FAx1_ASAP7_75t_SL g55 ( 
.A(n_54),
.B(n_53),
.CI(n_51),
.CON(n_55),
.SN(n_55)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_4),
.B(n_7),
.Y(n_56)
);

AOI21x1_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_55),
.B(n_13),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_10),
.B(n_14),
.C(n_17),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_SL g59 ( 
.A1(n_58),
.A2(n_26),
.B(n_21),
.C(n_22),
.Y(n_59)
);


endmodule