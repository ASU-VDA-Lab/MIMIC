module fake_jpeg_32109_n_328 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_44),
.B(n_60),
.Y(n_88)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_45),
.Y(n_114)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_17),
.B(n_13),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_50),
.B(n_62),
.Y(n_115)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_68),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_17),
.B(n_29),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_55),
.B(n_58),
.Y(n_110)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_57),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_18),
.B(n_26),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_18),
.B(n_0),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_37),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_61),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_26),
.B(n_9),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_32),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_64),
.Y(n_101)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_30),
.B(n_0),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_67),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_29),
.B(n_1),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_35),
.B(n_36),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_21),
.B(n_1),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_70),
.B(n_71),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_37),
.B(n_1),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_35),
.B(n_9),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_77),
.Y(n_92)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_36),
.B(n_2),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_71),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_27),
.B(n_8),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_61),
.A2(n_25),
.B1(n_21),
.B2(n_15),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_79),
.A2(n_82),
.B1(n_90),
.B2(n_109),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_52),
.A2(n_25),
.B1(n_32),
.B2(n_15),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_24),
.B1(n_25),
.B2(n_33),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_86),
.A2(n_57),
.B1(n_51),
.B2(n_56),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_55),
.B(n_33),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_95),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_61),
.A2(n_15),
.B1(n_28),
.B2(n_39),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_70),
.A2(n_32),
.B1(n_28),
.B2(n_39),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_91),
.A2(n_93),
.B1(n_125),
.B2(n_31),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_60),
.A2(n_32),
.B1(n_24),
.B2(n_20),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_24),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_38),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_106),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_77),
.B(n_22),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_38),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_121),
.Y(n_143)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_44),
.A2(n_22),
.B1(n_41),
.B2(n_40),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_111),
.B(n_28),
.Y(n_152)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_64),
.A2(n_28),
.B1(n_39),
.B2(n_20),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_119),
.A2(n_81),
.B1(n_72),
.B2(n_63),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_38),
.Y(n_121)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_67),
.B(n_43),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_38),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_66),
.A2(n_41),
.B1(n_40),
.B2(n_20),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_129),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_74),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_150),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_100),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_133),
.B(n_152),
.Y(n_182)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_137),
.A2(n_153),
.B1(n_103),
.B2(n_89),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_48),
.B(n_8),
.C(n_75),
.Y(n_138)
);

OAI32xp33_ASAP7_75t_L g175 ( 
.A1(n_138),
.A2(n_110),
.A3(n_39),
.B1(n_114),
.B2(n_83),
.Y(n_175)
);

NOR2x1_ASAP7_75t_R g141 ( 
.A(n_122),
.B(n_42),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_141),
.B(n_147),
.Y(n_193)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_145),
.B(n_146),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_80),
.B(n_38),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_149),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_45),
.Y(n_150)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_86),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_156),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_157),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_92),
.B(n_53),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_90),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_115),
.B(n_39),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_158),
.B(n_31),
.Y(n_186)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_79),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_161),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_91),
.B(n_53),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_165),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_85),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_163),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_120),
.A2(n_46),
.B1(n_69),
.B2(n_63),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_164),
.A2(n_99),
.B1(n_116),
.B2(n_96),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_115),
.B(n_72),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_130),
.C(n_154),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_168),
.B(n_181),
.C(n_183),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_173),
.A2(n_177),
.B1(n_189),
.B2(n_196),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_161),
.A2(n_100),
.B1(n_117),
.B2(n_89),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_174),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_153),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_162),
.A2(n_116),
.B1(n_96),
.B2(n_123),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_143),
.C(n_165),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_112),
.C(n_108),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_184),
.A2(n_197),
.B1(n_136),
.B2(n_140),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_186),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_157),
.A2(n_117),
.B1(n_126),
.B2(n_118),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_135),
.Y(n_191)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_191),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_155),
.B(n_126),
.C(n_118),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_153),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_147),
.A2(n_105),
.B1(n_85),
.B2(n_104),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_139),
.A2(n_104),
.B1(n_105),
.B2(n_94),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_142),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_198),
.Y(n_201)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_148),
.Y(n_199)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_199),
.Y(n_206)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_160),
.Y(n_200)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_203),
.Y(n_236)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_207),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_182),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_218),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_192),
.A2(n_138),
.B(n_132),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_210),
.A2(n_185),
.B(n_199),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_167),
.B(n_153),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_216),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_214),
.A2(n_219),
.B1(n_196),
.B2(n_189),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_169),
.B(n_127),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_215),
.B(n_223),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_167),
.B(n_134),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_170),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_195),
.A2(n_134),
.B1(n_164),
.B2(n_94),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_131),
.B1(n_140),
.B2(n_128),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_221),
.A2(n_227),
.B1(n_184),
.B2(n_169),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_171),
.B(n_159),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_224),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_168),
.B(n_128),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_178),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_131),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_225),
.B(n_228),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_144),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_193),
.C(n_194),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_193),
.A2(n_151),
.B1(n_144),
.B2(n_31),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_183),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_187),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_181),
.B(n_3),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_230),
.B(n_185),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_211),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_233),
.A2(n_235),
.B1(n_246),
.B2(n_219),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_208),
.B(n_175),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_239),
.B(n_240),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_215),
.Y(n_240)
);

AOI221xp5_ASAP7_75t_L g255 ( 
.A1(n_241),
.A2(n_242),
.B1(n_244),
.B2(n_210),
.C(n_216),
.Y(n_255)
);

OA21x2_ASAP7_75t_SL g244 ( 
.A1(n_225),
.A2(n_178),
.B(n_177),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_212),
.A2(n_200),
.B1(n_188),
.B2(n_191),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

INVxp67_ASAP7_75t_SL g254 ( 
.A(n_247),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_213),
.A2(n_187),
.B(n_179),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_250),
.A2(n_204),
.B(n_206),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_180),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_252),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_206),
.B(n_224),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_245),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_259),
.Y(n_274)
);

XNOR2x1_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_249),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_211),
.C(n_228),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_263),
.C(n_266),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_232),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_257),
.B(n_260),
.Y(n_271)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_251),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_232),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_235),
.A2(n_213),
.B1(n_204),
.B2(n_202),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_262),
.A2(n_270),
.B1(n_246),
.B2(n_243),
.Y(n_282)
);

NAND2x1_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_226),
.Y(n_265)
);

A2O1A1Ixp33_ASAP7_75t_SL g273 ( 
.A1(n_265),
.A2(n_269),
.B(n_242),
.C(n_244),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_227),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_268),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_240),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_273),
.A2(n_265),
.B(n_250),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_231),
.C(n_234),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_283),
.C(n_284),
.Y(n_290)
);

OAI321xp33_ASAP7_75t_L g276 ( 
.A1(n_264),
.A2(n_249),
.A3(n_236),
.B1(n_239),
.B2(n_234),
.C(n_261),
.Y(n_276)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_269),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_270),
.B(n_238),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_205),
.Y(n_293)
);

NOR3xp33_ASAP7_75t_SL g279 ( 
.A(n_261),
.B(n_238),
.C(n_241),
.Y(n_279)
);

NOR3xp33_ASAP7_75t_SL g294 ( 
.A(n_279),
.B(n_233),
.C(n_217),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_282),
.A2(n_248),
.B1(n_201),
.B2(n_207),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_256),
.B(n_242),
.C(n_237),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_237),
.C(n_246),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_281),
.A2(n_262),
.B1(n_258),
.B2(n_259),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_285),
.B(n_287),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_267),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_290),
.C(n_289),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_287),
.B(n_289),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_288),
.A2(n_296),
.B(n_166),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_265),
.Y(n_289)
);

XNOR2x1_ASAP7_75t_SL g292 ( 
.A(n_273),
.B(n_254),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_292),
.A2(n_297),
.B1(n_273),
.B2(n_279),
.Y(n_298)
);

OAI21x1_ASAP7_75t_L g302 ( 
.A1(n_293),
.A2(n_294),
.B(n_295),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_217),
.Y(n_295)
);

AOI321xp33_ASAP7_75t_L g296 ( 
.A1(n_277),
.A2(n_233),
.A3(n_253),
.B1(n_201),
.B2(n_248),
.C(n_180),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_298),
.A2(n_299),
.B1(n_292),
.B2(n_296),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_300),
.B(n_301),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_272),
.C(n_274),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_273),
.C(n_248),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_304),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_291),
.A2(n_188),
.B1(n_198),
.B2(n_176),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_220),
.C(n_176),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_307),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_166),
.C(n_172),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_308),
.A2(n_294),
.B(n_299),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_312),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_311),
.A2(n_306),
.B(n_163),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_302),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_306),
.A2(n_163),
.B1(n_4),
.B2(n_5),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_3),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_317),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_313),
.B(n_163),
.Y(n_317)
);

OAI321xp33_ASAP7_75t_L g318 ( 
.A1(n_311),
.A2(n_314),
.A3(n_315),
.B1(n_309),
.B2(n_310),
.C(n_7),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_318),
.A2(n_320),
.B1(n_3),
.B2(n_4),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_319),
.B(n_3),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_322),
.B(n_5),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_4),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_324),
.A2(n_325),
.B(n_6),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_321),
.C(n_6),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_6),
.C(n_42),
.Y(n_328)
);


endmodule