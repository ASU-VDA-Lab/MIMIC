module fake_jpeg_11451_n_133 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_133);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_14),
.B(n_31),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_4),
.B(n_12),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_33),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_9),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_54),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_0),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_59),
.B(n_41),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_50),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_64),
.Y(n_70)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_49),
.B1(n_42),
.B2(n_47),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_68),
.B(n_49),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_20),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_67),
.Y(n_69)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_42),
.A2(n_17),
.B1(n_37),
.B2(n_35),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_16),
.B(n_34),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_68),
.B(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_75),
.B(n_77),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_53),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_2),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_81),
.A2(n_2),
.B(n_3),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_44),
.Y(n_90)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_62),
.B1(n_61),
.B2(n_48),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_87),
.B1(n_89),
.B2(n_73),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_69),
.A2(n_44),
.B1(n_52),
.B2(n_55),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_80),
.B1(n_70),
.B2(n_82),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_91),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_58),
.Y(n_91)
);

AO22x1_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_50),
.B1(n_38),
.B2(n_30),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_92),
.B(n_94),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_50),
.B(n_3),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_95),
.C(n_98),
.Y(n_99)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_5),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_97),
.B(n_6),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_73),
.A2(n_28),
.B(n_27),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_107),
.B1(n_10),
.B2(n_11),
.Y(n_117)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_105),
.Y(n_121)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_5),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_110),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_87),
.A2(n_86),
.B1(n_96),
.B2(n_92),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_108),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_114)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_7),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_112),
.C(n_113),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_7),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_8),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_115),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_93),
.C(n_22),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_117),
.A2(n_118),
.B1(n_120),
.B2(n_99),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_12),
.B1(n_13),
.B2(n_21),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_23),
.C(n_24),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_102),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_104),
.A2(n_13),
.B1(n_26),
.B2(n_99),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_124),
.C(n_116),
.Y(n_127)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_126),
.A2(n_122),
.B1(n_105),
.B2(n_103),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_128),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_121),
.B(n_122),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_115),
.B(n_125),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_124),
.C(n_102),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_109),
.Y(n_133)
);


endmodule