module fake_jpeg_20192_n_42 (n_3, n_2, n_1, n_0, n_4, n_5, n_42);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_42;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

INVx3_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_0),
.B(n_2),
.Y(n_8)
);

INVx5_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx2_ASAP7_75t_SL g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_10),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_14)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_14),
.A2(n_16),
.B1(n_9),
.B2(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_10),
.A2(n_1),
.B1(n_5),
.B2(n_9),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_11),
.B(n_1),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_18),
.B(n_10),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_15),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_5),
.B(n_14),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_26),
.B1(n_27),
.B2(n_21),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_19),
.A2(n_18),
.B(n_11),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_21),
.C(n_6),
.Y(n_33)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_17),
.B1(n_23),
.B2(n_6),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_28),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_34),
.A2(n_23),
.B1(n_32),
.B2(n_29),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_36),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_30),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_28),
.Y(n_39)
);

BUFx24_ASAP7_75t_SL g40 ( 
.A(n_39),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_38),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_41),
.A2(n_37),
.B(n_7),
.Y(n_42)
);


endmodule