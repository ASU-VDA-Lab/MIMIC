module fake_jpeg_20929_n_213 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_213);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_213;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_165;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_33;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_37),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_30),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_19),
.B(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_41),
.Y(n_58)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_42),
.Y(n_54)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

OR2x4_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_40),
.Y(n_53)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_52),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_36),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_31),
.B1(n_28),
.B2(n_17),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_55),
.A2(n_24),
.B1(n_23),
.B2(n_16),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_37),
.B(n_41),
.Y(n_72)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_28),
.B1(n_30),
.B2(n_27),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_63),
.A2(n_45),
.B1(n_42),
.B2(n_24),
.Y(n_95)
);

BUFx8_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_64),
.Y(n_78)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_17),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_27),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_72),
.A2(n_82),
.B(n_2),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_94),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_70),
.B1(n_67),
.B2(n_58),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_74),
.A2(n_89),
.B1(n_98),
.B2(n_100),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_56),
.A2(n_29),
.B1(n_16),
.B2(n_40),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_75),
.A2(n_6),
.B(n_10),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_36),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_96),
.Y(n_114)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_47),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_91),
.B(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_64),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_65),
.B1(n_59),
.B2(n_64),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_57),
.B(n_42),
.Y(n_96)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_54),
.A2(n_23),
.B1(n_29),
.B2(n_27),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_60),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_4),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_54),
.A2(n_21),
.B1(n_27),
.B2(n_33),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_59),
.Y(n_101)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx3_ASAP7_75t_SL g133 ( 
.A(n_103),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_33),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_119),
.C(n_86),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_105),
.A2(n_110),
.B1(n_122),
.B2(n_123),
.Y(n_132)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_79),
.A2(n_33),
.B1(n_22),
.B2(n_18),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_1),
.B(n_2),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_113),
.A2(n_115),
.B(n_124),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_11),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_118),
.B(n_12),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_22),
.Y(n_119)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_89),
.A2(n_18),
.B1(n_5),
.B2(n_4),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_85),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_123)
);

NAND2xp67_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_5),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_75),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_126),
.B(n_128),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_124),
.A2(n_81),
.B1(n_99),
.B2(n_86),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_105),
.B1(n_117),
.B2(n_116),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_93),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_130),
.B(n_131),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_111),
.B(n_12),
.Y(n_131)
);

BUFx12_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_134),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_81),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_140),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_136),
.A2(n_142),
.B(n_123),
.Y(n_160)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_83),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_92),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_83),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_144),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_108),
.B(n_90),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_76),
.Y(n_163)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_146),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_149),
.B(n_156),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_125),
.C(n_122),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_159),
.C(n_129),
.Y(n_166)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_141),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_138),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_157),
.A2(n_160),
.B(n_136),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_110),
.C(n_106),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_106),
.B1(n_117),
.B2(n_92),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_142),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_155),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_164),
.B(n_171),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_167),
.C(n_169),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_135),
.C(n_142),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_143),
.B(n_129),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_151),
.Y(n_177)
);

NOR2x1p5_ASAP7_75t_SL g171 ( 
.A(n_154),
.B(n_132),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_173),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_137),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_174),
.B(n_175),
.Y(n_187)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_177),
.A2(n_146),
.B(n_134),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_160),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_139),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_176),
.A2(n_132),
.B1(n_161),
.B2(n_147),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_182),
.A2(n_185),
.B1(n_167),
.B2(n_147),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_150),
.C(n_159),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_173),
.C(n_148),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_186),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_176),
.A2(n_170),
.B1(n_168),
.B2(n_153),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_158),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_192),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_191),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_152),
.Y(n_191)
);

NOR2xp67_ASAP7_75t_SL g196 ( 
.A(n_193),
.B(n_194),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_139),
.C(n_87),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_133),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_195),
.A2(n_78),
.B1(n_77),
.B2(n_14),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_190),
.A2(n_180),
.B1(n_184),
.B2(n_178),
.Y(n_197)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_192),
.A2(n_187),
.B1(n_133),
.B2(n_87),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_195),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_201),
.B(n_200),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_204),
.Y(n_206)
);

FAx1_ASAP7_75t_SL g203 ( 
.A(n_197),
.B(n_191),
.CI(n_13),
.CON(n_203),
.SN(n_203)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_203),
.B(n_199),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_207),
.A2(n_208),
.B(n_206),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_199),
.Y(n_208)
);

AO21x1_ASAP7_75t_L g211 ( 
.A1(n_209),
.A2(n_210),
.B(n_203),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_208),
.A2(n_205),
.B(n_203),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_211),
.B(n_196),
.Y(n_212)
);

BUFx24_ASAP7_75t_SL g213 ( 
.A(n_212),
.Y(n_213)
);


endmodule