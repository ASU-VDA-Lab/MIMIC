module fake_ariane_2168_n_72 (n_8, n_3, n_2, n_11, n_7, n_16, n_5, n_14, n_1, n_0, n_12, n_15, n_6, n_13, n_9, n_17, n_4, n_10, n_72);

input n_8;
input n_3;
input n_2;
input n_11;
input n_7;
input n_16;
input n_5;
input n_14;
input n_1;
input n_0;
input n_12;
input n_15;
input n_6;
input n_13;
input n_9;
input n_17;
input n_4;
input n_10;

output n_72;

wire n_66;
wire n_56;
wire n_60;
wire n_24;
wire n_22;
wire n_71;
wire n_43;
wire n_49;
wire n_20;
wire n_27;
wire n_48;
wire n_29;
wire n_64;
wire n_41;
wire n_50;
wire n_38;
wire n_55;
wire n_62;
wire n_47;
wire n_32;
wire n_18;
wire n_28;
wire n_37;
wire n_58;
wire n_65;
wire n_51;
wire n_67;
wire n_45;
wire n_34;
wire n_69;
wire n_26;
wire n_46;
wire n_52;
wire n_36;
wire n_68;
wire n_33;
wire n_44;
wire n_19;
wire n_30;
wire n_40;
wire n_39;
wire n_59;
wire n_31;
wire n_42;
wire n_57;
wire n_63;
wire n_53;
wire n_21;
wire n_70;
wire n_23;
wire n_61;
wire n_35;
wire n_54;
wire n_25;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_5),
.B(n_17),
.Y(n_19)
);

OAI22xp33_ASAP7_75t_L g20 ( 
.A1(n_9),
.A2(n_12),
.B1(n_0),
.B2(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_15),
.A2(n_3),
.B1(n_2),
.B2(n_5),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_16),
.A2(n_3),
.B1(n_10),
.B2(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_13),
.A2(n_6),
.B1(n_1),
.B2(n_4),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_1),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_7),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_7),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2x1_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_19),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_19),
.B(n_30),
.C(n_23),
.Y(n_38)
);

AND2x4_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_32),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

OR2x6_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_26),
.Y(n_41)
);

O2A1O1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_23),
.B(n_30),
.C(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

OAI21x1_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_29),
.B(n_21),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_40),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_38),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_28),
.B1(n_18),
.B2(n_27),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

AO21x2_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_42),
.B(n_41),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_24),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_48),
.B1(n_46),
.B2(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_53),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_48),
.B1(n_44),
.B2(n_54),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_58),
.B(n_55),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_51),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_57),
.B(n_59),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_44),
.B(n_47),
.C(n_50),
.Y(n_64)
);

AOI221xp5_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_47),
.B1(n_51),
.B2(n_50),
.C(n_52),
.Y(n_65)
);

NAND4xp75_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_53),
.C(n_57),
.D(n_51),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_51),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_24),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_53),
.B1(n_44),
.B2(n_24),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_18),
.B1(n_68),
.B2(n_67),
.Y(n_71)
);

OR2x6_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_18),
.Y(n_72)
);


endmodule