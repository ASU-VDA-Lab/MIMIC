module fake_jpeg_970_n_536 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_536);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_536;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_361;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_341;
wire n_151;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_4),
.B(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_14),
.B(n_13),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_46),
.B(n_47),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_13),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_12),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_48),
.B(n_56),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_50),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_53),
.Y(n_122)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_54),
.Y(n_124)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_33),
.B(n_11),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_57),
.B(n_60),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

NOR2xp67_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_10),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_61),
.Y(n_141)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_19),
.B(n_9),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_63),
.B(n_65),
.Y(n_138)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_44),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_66),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx5_ASAP7_75t_SL g123 ( 
.A(n_68),
.Y(n_123)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_69),
.Y(n_160)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_70),
.Y(n_139)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_19),
.B(n_9),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_87),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_29),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_78),
.B(n_80),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_22),
.B(n_0),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_81),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

BUFx24_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_17),
.B(n_0),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_83),
.Y(n_129)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_21),
.B(n_9),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_24),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

BUFx16f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_89),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_21),
.B(n_9),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_95),
.Y(n_107)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_26),
.B(n_1),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_85),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_100),
.B(n_135),
.Y(n_183)
);

O2A1O1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_50),
.A2(n_43),
.B(n_42),
.C(n_35),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_103),
.B(n_121),
.Y(n_199)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_109),
.Y(n_172)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_118),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_57),
.B(n_34),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_65),
.B(n_34),
.Y(n_135)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_142),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_94),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_144),
.B(n_145),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_54),
.Y(n_145)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_58),
.Y(n_149)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_67),
.Y(n_153)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_153),
.Y(n_198)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_64),
.Y(n_154)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_78),
.B(n_30),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_156),
.B(n_36),
.Y(n_209)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_71),
.Y(n_157)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_84),
.Y(n_158)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_73),
.Y(n_159)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_113),
.B(n_83),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_162),
.Y(n_229)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_105),
.Y(n_164)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_164),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_83),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_166),
.B(n_202),
.Y(n_224)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

INVx13_ASAP7_75t_L g243 ( 
.A(n_167),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_72),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_171),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_88),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_185),
.Y(n_215)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_176),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_131),
.A2(n_25),
.B1(n_15),
.B2(n_39),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_177),
.A2(n_189),
.B1(n_28),
.B2(n_42),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_106),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_178),
.Y(n_216)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_125),
.Y(n_180)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_180),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_127),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_181),
.Y(n_219)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_110),
.Y(n_182)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_113),
.B(n_80),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_184),
.B(n_204),
.Y(n_227)
);

INVx5_ASAP7_75t_SL g185 ( 
.A(n_130),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_129),
.A2(n_96),
.B1(n_81),
.B2(n_75),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_186),
.A2(n_161),
.B1(n_122),
.B2(n_117),
.Y(n_211)
);

INVx4_ASAP7_75t_SL g187 ( 
.A(n_130),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_190),
.Y(n_223)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_143),
.Y(n_188)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_188),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_138),
.A2(n_25),
.B1(n_39),
.B2(n_15),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_116),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_127),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_192),
.B(n_193),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_148),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_132),
.Y(n_194)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_194),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_115),
.B(n_70),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_195),
.B(n_62),
.C(n_160),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_107),
.B(n_91),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_196),
.B(n_197),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_99),
.Y(n_197)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_200),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_115),
.B(n_31),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_104),
.Y(n_203)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_203),
.Y(n_247)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_119),
.Y(n_204)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_152),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_205),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_148),
.Y(n_206)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_206),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_137),
.B(n_50),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_207),
.B(n_208),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_99),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_36),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_114),
.A2(n_89),
.B1(n_97),
.B2(n_69),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_210),
.A2(n_111),
.B1(n_90),
.B2(n_61),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_211),
.A2(n_213),
.B1(n_214),
.B2(n_218),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_195),
.A2(n_133),
.B1(n_124),
.B2(n_161),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_186),
.A2(n_133),
.B1(n_124),
.B2(n_79),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_202),
.A2(n_128),
.B1(n_117),
.B2(n_122),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_199),
.A2(n_134),
.B1(n_136),
.B2(n_128),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_233),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_207),
.A2(n_101),
.B(n_102),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_230),
.A2(n_232),
.B(n_164),
.Y(n_261)
);

A2O1A1Ixp33_ASAP7_75t_L g232 ( 
.A1(n_166),
.A2(n_147),
.B(n_30),
.C(n_26),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_184),
.A2(n_146),
.B1(n_136),
.B2(n_134),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_245),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_191),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

INVxp33_ASAP7_75t_L g267 ( 
.A(n_240),
.Y(n_267)
);

AOI32xp33_ASAP7_75t_L g245 ( 
.A1(n_162),
.A2(n_108),
.A3(n_141),
.B1(n_86),
.B2(n_123),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_184),
.B(n_139),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_162),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_249),
.B(n_252),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_250),
.B(n_227),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_165),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_251),
.B(n_232),
.C(n_231),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_183),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_171),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_255),
.B(n_256),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_168),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_169),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_259),
.Y(n_290)
);

INVx8_ASAP7_75t_L g258 ( 
.A(n_243),
.Y(n_258)
);

INVx5_ASAP7_75t_L g301 ( 
.A(n_258),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_174),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_174),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_271),
.Y(n_292)
);

AO21x1_ASAP7_75t_L g309 ( 
.A1(n_261),
.A2(n_273),
.B(n_278),
.Y(n_309)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_212),
.Y(n_262)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_262),
.Y(n_282)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_263),
.Y(n_285)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_264),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_223),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_268),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_223),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_247),
.Y(n_269)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

INVx13_ASAP7_75t_L g270 ( 
.A(n_243),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_270),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_227),
.B(n_203),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_217),
.Y(n_272)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_272),
.Y(n_295)
);

AND2x6_ASAP7_75t_L g273 ( 
.A(n_229),
.B(n_185),
.Y(n_273)
);

INVx13_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_274),
.A2(n_187),
.B1(n_217),
.B2(n_200),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_226),
.A2(n_164),
.B(n_206),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_275),
.A2(n_215),
.B(n_231),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_216),
.Y(n_276)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_216),
.Y(n_277)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_277),
.Y(n_300)
);

AND2x6_ASAP7_75t_L g278 ( 
.A(n_229),
.B(n_167),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_266),
.A2(n_214),
.B1(n_218),
.B2(n_235),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_279),
.A2(n_280),
.B1(n_303),
.B2(n_308),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_266),
.A2(n_232),
.B1(n_226),
.B2(n_227),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_256),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_283),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_284),
.B(n_298),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_288),
.A2(n_296),
.B(n_307),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_252),
.A2(n_220),
.B1(n_230),
.B2(n_246),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_291),
.A2(n_248),
.B1(n_262),
.B2(n_225),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_265),
.B(n_234),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_293),
.B(n_304),
.Y(n_320)
);

BUFx12f_ASAP7_75t_L g317 ( 
.A(n_294),
.Y(n_317)
);

OR2x4_ASAP7_75t_L g296 ( 
.A(n_261),
.B(n_245),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_251),
.B(n_215),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_302),
.B(n_305),
.C(n_249),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_253),
.A2(n_211),
.B1(n_233),
.B2(n_198),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_255),
.B(n_219),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_250),
.B(n_219),
.C(n_247),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_275),
.A2(n_237),
.B(n_212),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_253),
.A2(n_221),
.B1(n_237),
.B2(n_222),
.Y(n_308)
);

OAI32xp33_ASAP7_75t_L g310 ( 
.A1(n_257),
.A2(n_221),
.A3(n_222),
.B1(n_169),
.B2(n_204),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_271),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_259),
.Y(n_311)
);

OAI221xp5_ASAP7_75t_L g354 ( 
.A1(n_311),
.A2(n_313),
.B1(n_316),
.B2(n_333),
.C(n_314),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_301),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_312),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_260),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_286),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_314),
.B(n_315),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_283),
.B(n_242),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_285),
.Y(n_318)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_318),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_306),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_319),
.B(n_323),
.Y(n_355)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_301),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_321),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_290),
.B(n_272),
.Y(n_322)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_322),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_306),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_285),
.Y(n_324)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_324),
.Y(n_357)
);

AND2x6_ASAP7_75t_L g325 ( 
.A(n_296),
.B(n_273),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_325),
.B(n_330),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_326),
.B(n_339),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_309),
.A2(n_273),
.B(n_254),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_327),
.A2(n_309),
.B(n_307),
.Y(n_346)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_287),
.Y(n_328)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_328),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_292),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_290),
.B(n_263),
.Y(n_332)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_332),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_302),
.B(n_242),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_287),
.Y(n_335)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_335),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_281),
.B(n_264),
.Y(n_336)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_336),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_298),
.B(n_278),
.C(n_269),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_337),
.B(n_342),
.C(n_182),
.Y(n_373)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_289),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_338),
.B(n_236),
.Y(n_374)
);

XOR2x1_ASAP7_75t_L g339 ( 
.A(n_288),
.B(n_278),
.Y(n_339)
);

FAx1_ASAP7_75t_SL g340 ( 
.A(n_284),
.B(n_267),
.CI(n_248),
.CON(n_340),
.SN(n_340)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_340),
.B(n_281),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_341),
.A2(n_282),
.B1(n_300),
.B2(n_297),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_305),
.B(n_225),
.C(n_262),
.Y(n_342)
);

AO22x1_ASAP7_75t_L g344 ( 
.A1(n_334),
.A2(n_309),
.B1(n_303),
.B2(n_279),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_344),
.B(n_340),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_346),
.A2(n_352),
.B(n_360),
.Y(n_377)
);

OAI21x1_ASAP7_75t_L g389 ( 
.A1(n_350),
.A2(n_366),
.B(n_370),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_334),
.A2(n_308),
.B1(n_280),
.B2(n_292),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_351),
.A2(n_358),
.B1(n_328),
.B2(n_324),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_329),
.A2(n_327),
.B(n_315),
.Y(n_352)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_354),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_331),
.B(n_289),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_356),
.B(n_373),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_330),
.A2(n_295),
.B1(n_300),
.B2(n_297),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_329),
.A2(n_282),
.B(n_295),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_320),
.B(n_228),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_362),
.B(n_365),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_363),
.A2(n_367),
.B1(n_318),
.B2(n_277),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_343),
.B(n_236),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_331),
.B(n_310),
.Y(n_366)
);

MAJx2_ASAP7_75t_L g382 ( 
.A(n_366),
.B(n_337),
.C(n_340),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_341),
.A2(n_277),
.B1(n_276),
.B2(n_258),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_322),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_368),
.B(n_372),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_332),
.A2(n_258),
.B(n_270),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_369),
.A2(n_371),
.B(n_274),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_339),
.A2(n_205),
.B(n_170),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_336),
.Y(n_372)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_374),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_378),
.A2(n_393),
.B1(n_398),
.B2(n_375),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_356),
.B(n_342),
.C(n_326),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_379),
.B(n_384),
.C(n_390),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_376),
.B(n_319),
.Y(n_380)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_380),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_349),
.B(n_321),
.Y(n_381)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_381),
.Y(n_423)
);

XNOR2x1_ASAP7_75t_L g427 ( 
.A(n_382),
.B(n_176),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_355),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_383),
.B(n_389),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_373),
.B(n_323),
.C(n_335),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_376),
.B(n_338),
.Y(n_385)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_385),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_386),
.A2(n_394),
.B1(n_405),
.B2(n_367),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_349),
.B(n_348),
.Y(n_387)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_387),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_388),
.A2(n_360),
.B(n_371),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_SL g390 ( 
.A(n_364),
.B(n_325),
.C(n_317),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_364),
.Y(n_392)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_392),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_351),
.A2(n_317),
.B1(n_276),
.B2(n_172),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_355),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_395),
.B(n_399),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_345),
.B(n_180),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_396),
.B(n_345),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_344),
.A2(n_317),
.B1(n_172),
.B2(n_201),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_370),
.B(n_358),
.Y(n_399)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_347),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_402),
.B(n_403),
.Y(n_421)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_347),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_353),
.A2(n_317),
.B1(n_201),
.B2(n_198),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_369),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_406),
.B(n_274),
.Y(n_432)
);

INVx13_ASAP7_75t_L g407 ( 
.A(n_383),
.Y(n_407)
);

INVx13_ASAP7_75t_L g446 ( 
.A(n_407),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_408),
.B(n_427),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_401),
.B(n_352),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_409),
.B(n_425),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_410),
.A2(n_416),
.B1(n_420),
.B2(n_429),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_414),
.A2(n_377),
.B(n_388),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_379),
.B(n_346),
.C(n_348),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_415),
.B(n_430),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_386),
.A2(n_344),
.B1(n_353),
.B2(n_363),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_417),
.A2(n_419),
.B1(n_406),
.B2(n_380),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_397),
.Y(n_418)
);

NOR3xp33_ASAP7_75t_L g448 ( 
.A(n_418),
.B(n_400),
.C(n_405),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_391),
.A2(n_375),
.B1(n_361),
.B2(n_357),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_395),
.A2(n_361),
.B1(n_357),
.B2(n_359),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_401),
.B(n_359),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_399),
.A2(n_179),
.B1(n_216),
.B2(n_146),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_384),
.B(n_175),
.C(n_194),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_404),
.B(n_228),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_431),
.B(n_433),
.Y(n_457)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_432),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_396),
.B(n_175),
.C(n_178),
.Y(n_433)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_434),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_423),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_435),
.B(n_445),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_441),
.A2(n_444),
.B(n_434),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_425),
.B(n_390),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_442),
.B(n_427),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_417),
.A2(n_378),
.B1(n_394),
.B2(n_398),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_443),
.A2(n_448),
.B1(n_450),
.B2(n_451),
.Y(n_473)
);

OAI21xp33_ASAP7_75t_L g444 ( 
.A1(n_411),
.A2(n_377),
.B(n_385),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_415),
.B(n_382),
.C(n_393),
.Y(n_445)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_421),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_447),
.B(n_449),
.Y(n_470)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_419),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_410),
.A2(n_179),
.B1(n_270),
.B2(n_140),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_416),
.A2(n_140),
.B1(n_126),
.B2(n_151),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_411),
.A2(n_170),
.B(n_120),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_452),
.A2(n_432),
.B(n_424),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_420),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_453),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_412),
.B(n_188),
.C(n_160),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_454),
.B(n_455),
.Y(n_466)
);

AOI322xp5_ASAP7_75t_L g455 ( 
.A1(n_428),
.A2(n_126),
.A3(n_77),
.B1(n_98),
.B2(n_27),
.C1(n_31),
.C2(n_228),
.Y(n_455)
);

AOI321xp33_ASAP7_75t_L g456 ( 
.A1(n_414),
.A2(n_163),
.A3(n_112),
.B1(n_152),
.B2(n_123),
.C(n_86),
.Y(n_456)
);

INVxp33_ASAP7_75t_SL g461 ( 
.A(n_456),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_440),
.B(n_412),
.C(n_409),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_458),
.B(n_464),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_459),
.B(n_462),
.Y(n_493)
);

AOI21xp33_ASAP7_75t_SL g482 ( 
.A1(n_462),
.A2(n_444),
.B(n_441),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_463),
.B(n_439),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_445),
.B(n_408),
.C(n_430),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_438),
.B(n_424),
.C(n_422),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_465),
.B(n_467),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_438),
.B(n_422),
.C(n_413),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_R g469 ( 
.A(n_436),
.B(n_426),
.C(n_407),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_469),
.B(n_471),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_453),
.B(n_433),
.C(n_429),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_457),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_472),
.B(n_476),
.Y(n_484)
);

INVx11_ASAP7_75t_L g474 ( 
.A(n_446),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_474),
.A2(n_477),
.B1(n_473),
.B2(n_471),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_442),
.B(n_49),
.C(n_31),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_437),
.A2(n_93),
.B1(n_31),
.B2(n_27),
.Y(n_477)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_479),
.Y(n_503)
);

AOI21xp33_ASAP7_75t_L g504 ( 
.A1(n_482),
.A2(n_483),
.B(n_493),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_468),
.B(n_454),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_458),
.B(n_443),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_485),
.B(n_486),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_465),
.B(n_451),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_487),
.B(n_59),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_464),
.B(n_439),
.C(n_446),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_488),
.B(n_489),
.C(n_463),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_467),
.B(n_456),
.C(n_82),
.Y(n_489)
);

OAI221xp5_ASAP7_75t_L g490 ( 
.A1(n_470),
.A2(n_28),
.B1(n_16),
.B2(n_35),
.C(n_42),
.Y(n_490)
);

AOI31xp67_ASAP7_75t_L g499 ( 
.A1(n_490),
.A2(n_35),
.A3(n_16),
.B(n_3),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_466),
.B(n_475),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_491),
.B(n_492),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_460),
.B(n_469),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_461),
.B(n_476),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_494),
.B(n_1),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_495),
.B(n_496),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_481),
.A2(n_474),
.B1(n_477),
.B2(n_28),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_497),
.B(n_502),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_499),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_478),
.A2(n_51),
.B(n_55),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_501),
.A2(n_482),
.B(n_489),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_480),
.A2(n_68),
.B1(n_43),
.B2(n_40),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_488),
.A2(n_43),
.B1(n_40),
.B2(n_23),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_505),
.B(n_479),
.C(n_20),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_483),
.B(n_23),
.C(n_40),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_506),
.B(n_507),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_484),
.B(n_20),
.C(n_2),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_508),
.B(n_1),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_510),
.B(n_513),
.Y(n_521)
);

NAND3xp33_ASAP7_75t_L g512 ( 
.A(n_503),
.B(n_498),
.C(n_504),
.Y(n_512)
);

NAND3xp33_ASAP7_75t_SL g522 ( 
.A(n_512),
.B(n_519),
.C(n_2),
.Y(n_522)
);

INVxp33_ASAP7_75t_L g525 ( 
.A(n_516),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_500),
.B(n_2),
.Y(n_517)
);

O2A1O1Ixp33_ASAP7_75t_SL g520 ( 
.A1(n_517),
.A2(n_518),
.B(n_508),
.C(n_506),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_495),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_496),
.A2(n_20),
.B(n_3),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_SL g529 ( 
.A1(n_520),
.A2(n_522),
.B(n_524),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_515),
.B(n_20),
.C(n_3),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_523),
.B(n_526),
.Y(n_527)
);

O2A1O1Ixp33_ASAP7_75t_SL g524 ( 
.A1(n_512),
.A2(n_20),
.B(n_4),
.C(n_5),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_518),
.B(n_2),
.C(n_4),
.Y(n_526)
);

AOI322xp5_ASAP7_75t_L g528 ( 
.A1(n_522),
.A2(n_514),
.A3(n_511),
.B1(n_509),
.B2(n_7),
.C1(n_6),
.C2(n_5),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_528),
.A2(n_521),
.B1(n_5),
.B2(n_6),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_525),
.B(n_4),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_530),
.B(n_4),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_531),
.Y(n_533)
);

OAI33xp33_ASAP7_75t_L g534 ( 
.A1(n_533),
.A2(n_529),
.A3(n_527),
.B1(n_532),
.B2(n_6),
.B3(n_5),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_534),
.B(n_6),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_535),
.B(n_7),
.Y(n_536)
);


endmodule