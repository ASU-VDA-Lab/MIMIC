module fake_ibex_2060_n_539 (n_64, n_3, n_73, n_65, n_55, n_63, n_29, n_2, n_76, n_8, n_67, n_9, n_38, n_37, n_47, n_10, n_21, n_27, n_16, n_78, n_60, n_70, n_7, n_20, n_69, n_75, n_48, n_57, n_59, n_28, n_39, n_5, n_62, n_71, n_13, n_61, n_14, n_0, n_12, n_42, n_77, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_58, n_43, n_22, n_4, n_33, n_30, n_6, n_72, n_26, n_34, n_15, n_24, n_52, n_1, n_25, n_36, n_41, n_45, n_18, n_32, n_53, n_50, n_11, n_68, n_79, n_35, n_31, n_56, n_23, n_54, n_19, n_539);

input n_64;
input n_3;
input n_73;
input n_65;
input n_55;
input n_63;
input n_29;
input n_2;
input n_76;
input n_8;
input n_67;
input n_9;
input n_38;
input n_37;
input n_47;
input n_10;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_70;
input n_7;
input n_20;
input n_69;
input n_75;
input n_48;
input n_57;
input n_59;
input n_28;
input n_39;
input n_5;
input n_62;
input n_71;
input n_13;
input n_61;
input n_14;
input n_0;
input n_12;
input n_42;
input n_77;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_58;
input n_43;
input n_22;
input n_4;
input n_33;
input n_30;
input n_6;
input n_72;
input n_26;
input n_34;
input n_15;
input n_24;
input n_52;
input n_1;
input n_25;
input n_36;
input n_41;
input n_45;
input n_18;
input n_32;
input n_53;
input n_50;
input n_11;
input n_68;
input n_79;
input n_35;
input n_31;
input n_56;
input n_23;
input n_54;
input n_19;

output n_539;

wire n_151;
wire n_85;
wire n_507;
wire n_395;
wire n_84;
wire n_171;
wire n_103;
wire n_529;
wire n_389;
wire n_204;
wire n_274;
wire n_387;
wire n_130;
wire n_177;
wire n_273;
wire n_330;
wire n_309;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_124;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_446;
wire n_108;
wire n_350;
wire n_165;
wire n_452;
wire n_86;
wire n_255;
wire n_175;
wire n_398;
wire n_125;
wire n_304;
wire n_191;
wire n_153;
wire n_194;
wire n_249;
wire n_334;
wire n_312;
wire n_478;
wire n_239;
wire n_134;
wire n_94;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_357;
wire n_88;
wire n_412;
wire n_457;
wire n_494;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_90;
wire n_449;
wire n_176;
wire n_216;
wire n_421;
wire n_475;
wire n_166;
wire n_163;
wire n_500;
wire n_114;
wire n_236;
wire n_376;
wire n_377;
wire n_531;
wire n_189;
wire n_498;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_105;
wire n_187;
wire n_154;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_89;
wire n_170;
wire n_144;
wire n_270;
wire n_346;
wire n_383;
wire n_113;
wire n_117;
wire n_417;
wire n_471;
wire n_265;
wire n_504;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_210;
wire n_348;
wire n_220;
wire n_91;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_228;
wire n_147;
wire n_251;
wire n_384;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_426;
wire n_323;
wire n_469;
wire n_143;
wire n_106;
wire n_386;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_333;
wire n_110;
wire n_306;
wire n_400;
wire n_169;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_109;
wire n_127;
wire n_121;
wire n_527;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_434;
wire n_296;
wire n_120;
wire n_168;
wire n_526;
wire n_155;
wire n_315;
wire n_441;
wire n_122;
wire n_523;
wire n_116;
wire n_370;
wire n_431;
wire n_289;
wire n_515;
wire n_150;
wire n_286;
wire n_321;
wire n_133;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_136;
wire n_261;
wire n_521;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_437;
wire n_355;
wire n_474;
wire n_490;
wire n_102;
wire n_407;
wire n_448;
wire n_99;
wire n_466;
wire n_269;
wire n_156;
wire n_126;
wire n_530;
wire n_356;
wire n_104;
wire n_420;
wire n_483;
wire n_141;
wire n_487;
wire n_222;
wire n_186;
wire n_524;
wire n_349;
wire n_454;
wire n_295;
wire n_331;
wire n_230;
wire n_96;
wire n_185;
wire n_388;
wire n_536;
wire n_352;
wire n_290;
wire n_174;
wire n_467;
wire n_427;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_438;
wire n_167;
wire n_128;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_205;
wire n_488;
wire n_139;
wire n_514;
wire n_429;
wire n_275;
wire n_98;
wire n_129;
wire n_267;
wire n_245;
wire n_229;
wire n_209;
wire n_472;
wire n_347;
wire n_473;
wire n_445;
wire n_335;
wire n_413;
wire n_82;
wire n_263;
wire n_353;
wire n_359;
wire n_299;
wire n_87;
wire n_262;
wire n_439;
wire n_433;
wire n_137;
wire n_338;
wire n_173;
wire n_477;
wire n_363;
wire n_402;
wire n_180;
wire n_369;
wire n_201;
wire n_351;
wire n_368;
wire n_456;
wire n_257;
wire n_401;
wire n_305;
wire n_307;
wire n_192;
wire n_140;
wire n_484;
wire n_480;
wire n_416;
wire n_365;
wire n_100;
wire n_179;
wire n_392;
wire n_206;
wire n_354;
wire n_516;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_199;
wire n_495;
wire n_410;
wire n_308;
wire n_463;
wire n_411;
wire n_135;
wire n_520;
wire n_512;
wire n_283;
wire n_366;
wire n_397;
wire n_111;
wire n_322;
wire n_227;
wire n_499;
wire n_115;
wire n_248;
wire n_92;
wire n_451;
wire n_101;
wire n_190;
wire n_138;
wire n_409;
wire n_238;
wire n_214;
wire n_332;
wire n_517;
wire n_211;
wire n_218;
wire n_314;
wire n_132;
wire n_277;
wire n_337;
wire n_522;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_535;
wire n_382;
wire n_502;
wire n_532;
wire n_95;
wire n_405;
wire n_415;
wire n_285;
wire n_288;
wire n_247;
wire n_320;
wire n_379;
wire n_291;
wire n_318;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_148;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_118;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_217;
wire n_324;
wire n_391;
wire n_537;
wire n_390;
wire n_178;
wire n_509;
wire n_303;
wire n_362;
wire n_93;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_501;
wire n_266;
wire n_294;
wire n_112;
wire n_485;
wire n_284;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_476;
wire n_461;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_119;
wire n_361;
wire n_455;
wire n_419;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_311;
wire n_406;
wire n_97;
wire n_197;
wire n_528;
wire n_181;
wire n_131;
wire n_123;
wire n_260;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_252;
wire n_396;
wire n_83;
wire n_107;
wire n_149;
wire n_489;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_81;
wire n_364;
wire n_159;
wire n_231;
wire n_202;
wire n_298;
wire n_160;
wire n_184;
wire n_492;
wire n_232;
wire n_380;
wire n_281;
wire n_425;

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_37),
.Y(n_81)
);

CKINVDCx5p33_ASAP7_75t_R g82 ( 
.A(n_70),
.Y(n_82)
);

CKINVDCx5p33_ASAP7_75t_R g83 ( 
.A(n_56),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_43),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_44),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_54),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g90 ( 
.A(n_75),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

CKINVDCx5p33_ASAP7_75t_R g92 ( 
.A(n_58),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

CKINVDCx5p33_ASAP7_75t_R g94 ( 
.A(n_45),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_23),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_18),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

CKINVDCx5p33_ASAP7_75t_R g100 ( 
.A(n_4),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_59),
.Y(n_101)
);

CKINVDCx5p33_ASAP7_75t_R g102 ( 
.A(n_72),
.Y(n_102)
);

NOR2xp67_ASAP7_75t_L g103 ( 
.A(n_17),
.B(n_6),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_11),
.Y(n_104)
);

BUFx10_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_33),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_42),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

CKINVDCx5p33_ASAP7_75t_R g110 ( 
.A(n_68),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_4),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_46),
.Y(n_113)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_57),
.Y(n_114)
);

NOR2xp67_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_52),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_32),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_74),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g118 ( 
.A(n_25),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_5),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_14),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_38),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_80),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_7),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_30),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_35),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_11),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_26),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_13),
.Y(n_129)
);

BUFx2_ASAP7_75t_SL g130 ( 
.A(n_79),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_50),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_36),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_62),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_13),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_1),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_10),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_27),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_51),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

AND2x4_ASAP7_75t_L g141 ( 
.A(n_97),
.B(n_0),
.Y(n_141)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

AND2x4_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_0),
.Y(n_145)
);

AND2x6_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_73),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_123),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_123),
.Y(n_148)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_134),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_91),
.B(n_2),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_112),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_88),
.Y(n_154)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_91),
.B(n_7),
.Y(n_156)
);

OAI21x1_ASAP7_75t_L g157 ( 
.A1(n_99),
.A2(n_34),
.B(n_66),
.Y(n_157)
);

OA21x2_ASAP7_75t_L g158 ( 
.A1(n_99),
.A2(n_29),
.B(n_64),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_8),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_88),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_9),
.Y(n_162)
);

AND2x4_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_9),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_12),
.Y(n_164)
);

AND2x4_ASAP7_75t_L g165 ( 
.A(n_124),
.B(n_12),
.Y(n_165)
);

AND2x4_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_14),
.Y(n_166)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_104),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_86),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_87),
.B(n_15),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_109),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_109),
.Y(n_171)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_82),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_109),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_109),
.Y(n_174)
);

AND2x4_ASAP7_75t_L g175 ( 
.A(n_93),
.B(n_15),
.Y(n_175)
);

BUFx8_ASAP7_75t_SL g176 ( 
.A(n_112),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_81),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g178 ( 
.A(n_126),
.Y(n_178)
);

BUFx8_ASAP7_75t_L g179 ( 
.A(n_96),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_85),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_98),
.Y(n_181)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_111),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_129),
.Y(n_184)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_111),
.Y(n_185)
);

AND2x6_ASAP7_75t_L g186 ( 
.A(n_121),
.B(n_67),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_136),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_89),
.Y(n_188)
);

AND2x4_ASAP7_75t_L g189 ( 
.A(n_133),
.B(n_16),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_137),
.Y(n_190)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_111),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_108),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_192)
);

OAI22x1_ASAP7_75t_R g193 ( 
.A1(n_122),
.A2(n_22),
.B1(n_40),
.B2(n_48),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_130),
.Y(n_194)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_127),
.Y(n_195)
);

AND2x4_ASAP7_75t_L g196 ( 
.A(n_103),
.B(n_49),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_83),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_142),
.B(n_114),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_142),
.B(n_110),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_152),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_163),
.Y(n_203)
);

AO21x2_ASAP7_75t_L g204 ( 
.A1(n_151),
.A2(n_115),
.B(n_132),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_106),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_163),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_102),
.Y(n_208)
);

AO21x2_ASAP7_75t_L g209 ( 
.A1(n_151),
.A2(n_127),
.B(n_138),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_140),
.B(n_101),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_140),
.B(n_116),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_156),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_156),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_160),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_170),
.Y(n_215)
);

AOI21x1_ASAP7_75t_L g216 ( 
.A1(n_159),
.A2(n_127),
.B(n_131),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_162),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_167),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_165),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_162),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_164),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_95),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_164),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_196),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_145),
.A2(n_141),
.B1(n_192),
.B2(n_150),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_175),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_147),
.Y(n_228)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_146),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_161),
.B(n_94),
.Y(n_230)
);

AND2x6_ASAP7_75t_L g231 ( 
.A(n_175),
.B(n_127),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_172),
.B(n_92),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_148),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_177),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_189),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_194),
.B(n_167),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_141),
.B(n_117),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_178),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_171),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_146),
.Y(n_240)
);

CKINVDCx6p67_ASAP7_75t_R g241 ( 
.A(n_184),
.Y(n_241)
);

NOR2x1p5_ASAP7_75t_L g242 ( 
.A(n_176),
.B(n_90),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_169),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_169),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_182),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_180),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_173),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_182),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_139),
.B(n_118),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_174),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_182),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_191),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_191),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_143),
.B(n_144),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_149),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_190),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_149),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_149),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_149),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_190),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_181),
.B(n_53),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_158),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_212),
.B(n_186),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_244),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_213),
.Y(n_265)
);

BUFx6f_ASAP7_75t_SL g266 ( 
.A(n_231),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_229),
.B(n_179),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_213),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_226),
.A2(n_179),
.B1(n_153),
.B2(n_183),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_245),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_217),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_217),
.B(n_168),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_248),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_240),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_220),
.B(n_146),
.Y(n_275)
);

INVxp33_ASAP7_75t_L g276 ( 
.A(n_222),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_220),
.B(n_186),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_221),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_241),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_221),
.B(n_223),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_248),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_223),
.B(n_186),
.Y(n_282)
);

AOI222xp33_ASAP7_75t_L g283 ( 
.A1(n_254),
.A2(n_176),
.B1(n_193),
.B2(n_155),
.C1(n_185),
.C2(n_195),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_251),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_251),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_155),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_256),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_252),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_240),
.Y(n_289)
);

BUFx5_ASAP7_75t_L g290 ( 
.A(n_240),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_224),
.B(n_55),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_241),
.B(n_60),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_252),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_260),
.Y(n_294)
);

O2A1O1Ixp5_ASAP7_75t_L g295 ( 
.A1(n_216),
.A2(n_198),
.B(n_262),
.C(n_236),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_253),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_230),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_225),
.B(n_227),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_225),
.B(n_227),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_218),
.B(n_237),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_253),
.Y(n_301)
);

NOR3xp33_ASAP7_75t_L g302 ( 
.A(n_246),
.B(n_234),
.C(n_208),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_210),
.B(n_211),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_206),
.B(n_232),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_235),
.B(n_203),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_203),
.B(n_207),
.Y(n_306)
);

INVx8_ASAP7_75t_L g307 ( 
.A(n_231),
.Y(n_307)
);

OAI22x1_ASAP7_75t_L g308 ( 
.A1(n_269),
.A2(n_242),
.B1(n_238),
.B2(n_201),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_263),
.A2(n_262),
.B(n_198),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_280),
.B(n_219),
.Y(n_310)
);

OAI21xp33_ASAP7_75t_L g311 ( 
.A1(n_268),
.A2(n_249),
.B(n_201),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_280),
.B(n_200),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_307),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_295),
.A2(n_216),
.B(n_261),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_263),
.A2(n_231),
.B(n_199),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_282),
.A2(n_209),
.B(n_204),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_279),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_265),
.B(n_233),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_271),
.B(n_204),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_282),
.A2(n_209),
.B(n_204),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_278),
.B(n_231),
.Y(n_321)
);

AOI21xp33_ASAP7_75t_L g322 ( 
.A1(n_275),
.A2(n_209),
.B(n_259),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_297),
.A2(n_242),
.B1(n_228),
.B2(n_202),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_277),
.A2(n_255),
.B(n_258),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_276),
.B(n_257),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_300),
.B(n_257),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_307),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_272),
.B(n_304),
.Y(n_328)
);

AND2x4_ASAP7_75t_L g329 ( 
.A(n_292),
.B(n_247),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_283),
.B(n_205),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_307),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_303),
.B(n_250),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_306),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_298),
.A2(n_299),
.B(n_291),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_270),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_302),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_287),
.B(n_214),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_R g338 ( 
.A(n_266),
.B(n_215),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_266),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_305),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_286),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_294),
.Y(n_342)
);

AND2x4_ASAP7_75t_L g343 ( 
.A(n_267),
.B(n_239),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_274),
.Y(n_344)
);

NOR2xp67_ASAP7_75t_L g345 ( 
.A(n_273),
.B(n_281),
.Y(n_345)
);

BUFx12f_ASAP7_75t_L g346 ( 
.A(n_274),
.Y(n_346)
);

BUFx12f_ASAP7_75t_L g347 ( 
.A(n_289),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_284),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_285),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_328),
.B(n_288),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_310),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_334),
.A2(n_293),
.B(n_296),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_310),
.B(n_301),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_336),
.A2(n_290),
.B1(n_330),
.B2(n_311),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_346),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_342),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_316),
.A2(n_320),
.B(n_314),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_325),
.B(n_341),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_322),
.A2(n_324),
.B(n_312),
.Y(n_359)
);

AND2x4_ASAP7_75t_L g360 ( 
.A(n_333),
.B(n_340),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_313),
.B(n_331),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_332),
.A2(n_315),
.B(n_321),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_347),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_308),
.B(n_323),
.Y(n_364)
);

AND2x4_ASAP7_75t_L g365 ( 
.A(n_327),
.B(n_313),
.Y(n_365)
);

BUFx12f_ASAP7_75t_L g366 ( 
.A(n_329),
.Y(n_366)
);

AO22x1_ASAP7_75t_L g367 ( 
.A1(n_339),
.A2(n_329),
.B1(n_335),
.B2(n_326),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_345),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_348),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_338),
.B(n_344),
.Y(n_370)
);

OAI21x1_ASAP7_75t_SL g371 ( 
.A1(n_349),
.A2(n_344),
.B(n_318),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_337),
.B(n_343),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_328),
.B(n_264),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_316),
.A2(n_320),
.B(n_295),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_328),
.B(n_264),
.Y(n_375)
);

AO31x2_ASAP7_75t_L g376 ( 
.A1(n_316),
.A2(n_320),
.A3(n_319),
.B(n_198),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_342),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_328),
.B(n_264),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_328),
.B(n_264),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_346),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_309),
.A2(n_320),
.B(n_316),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_328),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_342),
.Y(n_383)
);

OAI21x1_ASAP7_75t_SL g384 ( 
.A1(n_328),
.A2(n_280),
.B(n_310),
.Y(n_384)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_328),
.B(n_188),
.Y(n_385)
);

AO31x2_ASAP7_75t_L g386 ( 
.A1(n_316),
.A2(n_320),
.A3(n_319),
.B(n_198),
.Y(n_386)
);

AOI21xp33_ASAP7_75t_L g387 ( 
.A1(n_328),
.A2(n_276),
.B(n_297),
.Y(n_387)
);

INVxp33_ASAP7_75t_L g388 ( 
.A(n_328),
.Y(n_388)
);

AO31x2_ASAP7_75t_L g389 ( 
.A1(n_316),
.A2(n_320),
.A3(n_319),
.B(n_198),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_342),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_328),
.B(n_264),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_328),
.Y(n_392)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_346),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_342),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_346),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_328),
.B(n_264),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_328),
.B(n_264),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_328),
.B(n_264),
.Y(n_398)
);

INVx2_ASAP7_75t_SL g399 ( 
.A(n_317),
.Y(n_399)
);

AO21x2_ASAP7_75t_L g400 ( 
.A1(n_314),
.A2(n_322),
.B(n_320),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_355),
.Y(n_401)
);

INVx6_ASAP7_75t_L g402 ( 
.A(n_393),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_382),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_388),
.B(n_392),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_392),
.Y(n_405)
);

NAND2x1p5_ASAP7_75t_L g406 ( 
.A(n_375),
.B(n_379),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_379),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_366),
.Y(n_408)
);

OA21x2_ASAP7_75t_L g409 ( 
.A1(n_357),
.A2(n_374),
.B(n_381),
.Y(n_409)
);

AO21x2_ASAP7_75t_L g410 ( 
.A1(n_359),
.A2(n_400),
.B(n_384),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_373),
.B(n_378),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_391),
.B(n_396),
.Y(n_412)
);

INVx6_ASAP7_75t_L g413 ( 
.A(n_393),
.Y(n_413)
);

OR2x6_ASAP7_75t_L g414 ( 
.A(n_397),
.B(n_398),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_351),
.Y(n_415)
);

NAND2x1p5_ASAP7_75t_L g416 ( 
.A(n_360),
.B(n_351),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_358),
.B(n_387),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_356),
.Y(n_418)
);

OAI21x1_ASAP7_75t_L g419 ( 
.A1(n_352),
.A2(n_371),
.B(n_362),
.Y(n_419)
);

INVx8_ASAP7_75t_L g420 ( 
.A(n_363),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_377),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_350),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_363),
.Y(n_423)
);

OA21x2_ASAP7_75t_L g424 ( 
.A1(n_354),
.A2(n_364),
.B(n_386),
.Y(n_424)
);

AO31x2_ASAP7_75t_L g425 ( 
.A1(n_376),
.A2(n_386),
.A3(n_389),
.B(n_394),
.Y(n_425)
);

BUFx2_ASAP7_75t_SL g426 ( 
.A(n_380),
.Y(n_426)
);

NAND2x1p5_ASAP7_75t_L g427 ( 
.A(n_365),
.B(n_370),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_395),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_383),
.Y(n_429)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_399),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_390),
.B(n_372),
.Y(n_431)
);

NAND3xp33_ASAP7_75t_L g432 ( 
.A(n_367),
.B(n_368),
.C(n_385),
.Y(n_432)
);

OAI21x1_ASAP7_75t_L g433 ( 
.A1(n_361),
.A2(n_369),
.B(n_353),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_392),
.B(n_375),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_388),
.B(n_382),
.Y(n_435)
);

NOR2xp67_ASAP7_75t_L g436 ( 
.A(n_393),
.B(n_382),
.Y(n_436)
);

INVx5_ASAP7_75t_L g437 ( 
.A(n_375),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_355),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_392),
.B(n_375),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_355),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_414),
.A2(n_422),
.B1(n_412),
.B2(n_411),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_425),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_422),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_411),
.B(n_412),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_417),
.A2(n_434),
.B1(n_439),
.B2(n_404),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_432),
.A2(n_435),
.B(n_433),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_418),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_421),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_406),
.A2(n_416),
.B(n_404),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_409),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_415),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_437),
.B(n_410),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_438),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_437),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_440),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_429),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_450),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_452),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_442),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g460 ( 
.A(n_443),
.B(n_424),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_454),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_451),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_454),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_452),
.B(n_419),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_441),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_453),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_459),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_461),
.B(n_455),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_462),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_462),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_458),
.B(n_452),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_457),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_465),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_461),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_458),
.B(n_464),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_472),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_473),
.B(n_465),
.Y(n_477)
);

INVxp67_ASAP7_75t_SL g478 ( 
.A(n_472),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_469),
.B(n_445),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_470),
.B(n_460),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_475),
.B(n_458),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_467),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_474),
.B(n_461),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_477),
.B(n_479),
.Y(n_484)
);

INVx3_ASAP7_75t_SL g485 ( 
.A(n_483),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_481),
.B(n_475),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_478),
.B(n_474),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_481),
.B(n_475),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_480),
.B(n_471),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_476),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_476),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_490),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_484),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_485),
.A2(n_449),
.B1(n_468),
.B2(n_463),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_491),
.Y(n_495)
);

AOI222xp33_ASAP7_75t_L g496 ( 
.A1(n_485),
.A2(n_444),
.B1(n_403),
.B2(n_447),
.C1(n_456),
.C2(n_448),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_491),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_489),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_493),
.B(n_487),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_495),
.Y(n_500)
);

OAI21xp33_ASAP7_75t_L g501 ( 
.A1(n_494),
.A2(n_487),
.B(n_486),
.Y(n_501)
);

AOI221xp5_ASAP7_75t_L g502 ( 
.A1(n_498),
.A2(n_482),
.B1(n_488),
.B2(n_446),
.C(n_444),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_499),
.B(n_497),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_501),
.B(n_496),
.Y(n_504)
);

OAI221xp5_ASAP7_75t_L g505 ( 
.A1(n_502),
.A2(n_496),
.B1(n_492),
.B2(n_449),
.C(n_466),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_504),
.B(n_500),
.Y(n_506)
);

OAI211xp5_ASAP7_75t_SL g507 ( 
.A1(n_505),
.A2(n_445),
.B(n_435),
.C(n_423),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_506),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_507),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_508),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_509),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_510),
.B(n_503),
.Y(n_512)
);

NAND4xp75_ASAP7_75t_L g513 ( 
.A(n_511),
.B(n_436),
.C(n_438),
.D(n_426),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_513),
.A2(n_510),
.B1(n_428),
.B2(n_402),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_512),
.Y(n_515)
);

AND3x4_ASAP7_75t_L g516 ( 
.A(n_513),
.B(n_401),
.C(n_440),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_515),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_514),
.Y(n_518)
);

NOR2x1_ASAP7_75t_L g519 ( 
.A(n_516),
.B(n_408),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_515),
.A2(n_402),
.B1(n_413),
.B2(n_428),
.Y(n_520)
);

AO21x1_ASAP7_75t_L g521 ( 
.A1(n_515),
.A2(n_430),
.B(n_413),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_516),
.A2(n_402),
.B1(n_413),
.B2(n_401),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_517),
.Y(n_523)
);

AO22x2_ASAP7_75t_L g524 ( 
.A1(n_519),
.A2(n_430),
.B1(n_423),
.B2(n_420),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_518),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_521),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_522),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_520),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_518),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_518),
.Y(n_530)
);

AO21x2_ASAP7_75t_L g531 ( 
.A1(n_529),
.A2(n_420),
.B(n_431),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_530),
.A2(n_525),
.B1(n_528),
.B2(n_527),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_523),
.Y(n_533)
);

OAI21x1_ASAP7_75t_SL g534 ( 
.A1(n_532),
.A2(n_526),
.B(n_523),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_533),
.A2(n_524),
.B1(n_531),
.B2(n_420),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_535),
.A2(n_431),
.B(n_405),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_536),
.A2(n_534),
.B(n_427),
.Y(n_537)
);

OR2x6_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_454),
.Y(n_538)
);

AOI21xp33_ASAP7_75t_SL g539 ( 
.A1(n_538),
.A2(n_407),
.B(n_427),
.Y(n_539)
);


endmodule