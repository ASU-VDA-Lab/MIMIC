module fake_jpeg_23749_n_282 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_282);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_282;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_7),
.B(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_30),
.B(n_36),
.Y(n_52)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_33),
.Y(n_40)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_35),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_20),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_22),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_37),
.A2(n_18),
.B1(n_28),
.B2(n_21),
.Y(n_43)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NAND2xp33_ASAP7_75t_SL g39 ( 
.A(n_33),
.B(n_17),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_39),
.A2(n_43),
.B(n_16),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_18),
.B1(n_21),
.B2(n_28),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_41),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_21),
.B1(n_28),
.B2(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_31),
.A2(n_18),
.B1(n_19),
.B2(n_23),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_31),
.A2(n_19),
.B1(n_23),
.B2(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_55),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_29),
.A2(n_19),
.B1(n_23),
.B2(n_27),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_53),
.A2(n_29),
.B1(n_24),
.B2(n_14),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_36),
.B(n_27),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_57),
.B(n_17),
.Y(n_80)
);

BUFx2_ASAP7_75t_R g58 ( 
.A(n_33),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_58),
.Y(n_73)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_60),
.Y(n_103)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_54),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_53),
.B(n_14),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_63),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_64),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_69),
.A2(n_75),
.B1(n_78),
.B2(n_79),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_52),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_70),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_47),
.A2(n_27),
.B1(n_16),
.B2(n_14),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_71),
.A2(n_77),
.B(n_25),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_72),
.A2(n_62),
.B1(n_75),
.B2(n_61),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_52),
.B(n_24),
.Y(n_74)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_45),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_85),
.B(n_17),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_SL g87 ( 
.A1(n_68),
.A2(n_39),
.B(n_41),
.C(n_35),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_87),
.A2(n_91),
.B(n_97),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_48),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_38),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_69),
.A2(n_68),
.B1(n_63),
.B2(n_70),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_92),
.A2(n_93),
.B1(n_99),
.B2(n_100),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_60),
.A2(n_42),
.B1(n_49),
.B2(n_55),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_95),
.A2(n_96),
.B1(n_101),
.B2(n_35),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_67),
.A2(n_73),
.B1(n_59),
.B2(n_49),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_67),
.A2(n_48),
.B(n_50),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_61),
.A2(n_37),
.B1(n_34),
.B2(n_56),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_51),
.B1(n_35),
.B2(n_37),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_80),
.A2(n_34),
.B1(n_37),
.B2(n_30),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_50),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_65),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_73),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_113),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_65),
.B(n_30),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_106),
.A2(n_112),
.B(n_117),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_84),
.A2(n_75),
.B1(n_79),
.B2(n_66),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

INVxp33_ASAP7_75t_SL g109 ( 
.A(n_94),
.Y(n_109)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_123),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_34),
.B1(n_64),
.B2(n_66),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_85),
.A2(n_57),
.B(n_24),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_76),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_25),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_119),
.Y(n_133)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_116),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_38),
.B1(n_40),
.B2(n_64),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_97),
.C(n_101),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_87),
.A2(n_38),
.B1(n_40),
.B2(n_78),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_66),
.B1(n_40),
.B2(n_76),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_89),
.B(n_13),
.Y(n_122)
);

BUFx24_ASAP7_75t_SL g137 ( 
.A(n_122),
.Y(n_137)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_32),
.Y(n_124)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_83),
.A2(n_82),
.B(n_81),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_125),
.A2(n_88),
.B(n_94),
.Y(n_150)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_142),
.C(n_32),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_124),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_129),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_113),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_130),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_125),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_132),
.B(n_105),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_149),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_107),
.B(n_82),
.Y(n_135)
);

AOI32xp33_ASAP7_75t_L g151 ( 
.A1(n_135),
.A2(n_104),
.A3(n_112),
.B1(n_110),
.B2(n_117),
.Y(n_151)
);

AO21x2_ASAP7_75t_SL g140 ( 
.A1(n_111),
.A2(n_96),
.B(n_87),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_140),
.A2(n_141),
.B(n_148),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_107),
.A2(n_86),
.B(n_81),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_88),
.C(n_102),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_118),
.A2(n_87),
.B1(n_93),
.B2(n_99),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_144),
.A2(n_147),
.B1(n_26),
.B2(n_15),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_120),
.A2(n_95),
.B1(n_89),
.B2(n_96),
.Y(n_147)
);

AOI21x1_ASAP7_75t_SL g148 ( 
.A1(n_123),
.A2(n_96),
.B(n_32),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_96),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_150),
.A2(n_17),
.B(n_15),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_151),
.B(n_149),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_140),
.A2(n_126),
.B1(n_116),
.B2(n_115),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_154),
.A2(n_148),
.B1(n_131),
.B2(n_143),
.Y(n_183)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_163),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_121),
.Y(n_156)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_140),
.A2(n_105),
.B1(n_122),
.B2(n_84),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_157),
.A2(n_159),
.B1(n_168),
.B2(n_170),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_134),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_141),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_161),
.Y(n_189)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_174),
.C(n_142),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_128),
.B(n_17),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_145),
.B(n_17),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_171),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_32),
.Y(n_165)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_169),
.Y(n_181)
);

AOI322xp5_ASAP7_75t_L g169 ( 
.A1(n_135),
.A2(n_26),
.A3(n_15),
.B1(n_13),
.B2(n_12),
.C1(n_10),
.C2(n_9),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_170),
.A2(n_173),
.B1(n_143),
.B2(n_146),
.Y(n_179)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_13),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_140),
.A2(n_134),
.B1(n_144),
.B2(n_147),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_127),
.B(n_15),
.C(n_1),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_161),
.C(n_10),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_133),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_184),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_179),
.A2(n_196),
.B1(n_171),
.B2(n_156),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_SL g209 ( 
.A(n_180),
.B(n_194),
.C(n_156),
.Y(n_209)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_183),
.A2(n_185),
.B1(n_182),
.B2(n_187),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_138),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_154),
.A2(n_138),
.B1(n_137),
.B2(n_2),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_153),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_186),
.Y(n_206)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_167),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_193),
.Y(n_213)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

NOR2xp67_ASAP7_75t_SL g194 ( 
.A(n_160),
.B(n_12),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_12),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_157),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_174),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_201),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_215),
.C(n_185),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_189),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_203),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_159),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_184),
.B(n_173),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_202),
.B(n_209),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_175),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_205),
.B(n_207),
.Y(n_223)
);

MAJx2_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_152),
.C(n_155),
.Y(n_210)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_210),
.Y(n_216)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_214),
.Y(n_217)
);

INVxp33_ASAP7_75t_L g214 ( 
.A(n_190),
.Y(n_214)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_214),
.Y(n_221)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_206),
.B(n_211),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_218),
.B(n_225),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_210),
.Y(n_219)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_181),
.C(n_9),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_200),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_1),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_183),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_228),
.Y(n_235)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_215),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_0),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_208),
.A2(n_179),
.B1(n_196),
.B2(n_201),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_232),
.A2(n_199),
.B1(n_195),
.B2(n_198),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_232),
.B(n_198),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_3),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_237),
.B1(n_220),
.B2(n_227),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_220),
.A2(n_216),
.B1(n_223),
.B2(n_221),
.Y(n_237)
);

BUFx24_ASAP7_75t_SL g238 ( 
.A(n_230),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_246),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_222),
.B(n_181),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_240),
.B(n_227),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_245),
.C(n_3),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_242),
.A2(n_244),
.B(n_2),
.Y(n_249)
);

NOR2x1_ASAP7_75t_R g244 ( 
.A(n_231),
.B(n_0),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_0),
.C(n_1),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_254),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_249),
.B(n_253),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_230),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_250),
.B(n_251),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_2),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_257),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_235),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_255),
.B(n_4),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_243),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_4),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_4),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_241),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_263),
.Y(n_267)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_261),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_248),
.A2(n_244),
.B1(n_5),
.B2(n_6),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_265),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_5),
.Y(n_265)
);

OAI21x1_ASAP7_75t_L g268 ( 
.A1(n_258),
.A2(n_247),
.B(n_255),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_270),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_256),
.C(n_6),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_5),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_271),
.B(n_262),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_273),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_272),
.B(n_262),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_274),
.A2(n_275),
.B(n_269),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_267),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_R g279 ( 
.A(n_278),
.B(n_276),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_277),
.C(n_7),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_8),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_8),
.Y(n_282)
);


endmodule