module fake_aes_8261_n_11 (n_1, n_2, n_0, n_11);
input n_1;
input n_2;
input n_0;
output n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
OR2x6_ASAP7_75t_L g3 ( .A(n_1), .B(n_0), .Y(n_3) );
NAND2xp5_ASAP7_75t_SL g4 ( .A(n_2), .B(n_0), .Y(n_4) );
OR2x2_ASAP7_75t_L g5 ( .A(n_3), .B(n_0), .Y(n_5) );
INVx1_ASAP7_75t_L g6 ( .A(n_3), .Y(n_6) );
BUFx2_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
A2O1A1Ixp33_ASAP7_75t_L g8 ( .A1(n_7), .A2(n_6), .B(n_4), .C(n_1), .Y(n_8) );
OAI211xp5_ASAP7_75t_L g9 ( .A1(n_8), .A2(n_2), .B(n_0), .C(n_1), .Y(n_9) );
HB1xp67_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
AO21x2_ASAP7_75t_L g11 ( .A1(n_10), .A2(n_2), .B(n_1), .Y(n_11) );
endmodule