module fake_jpeg_136_n_437 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_437);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_437;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_0),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_SL g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_44),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_46),
.B(n_50),
.Y(n_91)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_47),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_48),
.Y(n_132)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_51),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_18),
.B(n_1),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_57),
.Y(n_86)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_18),
.B(n_1),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_73),
.Y(n_95)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_62),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_27),
.B(n_1),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_67),
.Y(n_98)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_69),
.Y(n_108)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_70),
.Y(n_128)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

HAxp5_ASAP7_75t_SL g107 ( 
.A(n_71),
.B(n_2),
.CON(n_107),
.SN(n_107)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_72),
.B(n_75),
.Y(n_120)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_76),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_79),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_80),
.Y(n_87)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_41),
.B(n_1),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_83),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_37),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_82),
.A2(n_16),
.B(n_3),
.Y(n_126)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_33),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_84),
.B(n_85),
.Y(n_130)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_43),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_92),
.B(n_100),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_62),
.A2(n_37),
.B1(n_20),
.B2(n_39),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_93),
.A2(n_103),
.B1(n_114),
.B2(n_131),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_34),
.B1(n_42),
.B2(n_38),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_99),
.A2(n_54),
.B1(n_9),
.B2(n_10),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_52),
.B(n_43),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_51),
.B(n_43),
.C(n_24),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_102),
.B(n_67),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_45),
.A2(n_24),
.B1(n_38),
.B2(n_34),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_39),
.B(n_32),
.C(n_23),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_104),
.B(n_127),
.Y(n_147)
);

INVx6_ASAP7_75t_SL g146 ( 
.A(n_107),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_48),
.B(n_24),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_111),
.B(n_115),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_71),
.A2(n_32),
.B(n_23),
.C(n_20),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_65),
.A2(n_16),
.B1(n_38),
.B2(n_42),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_69),
.B(n_19),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_75),
.B(n_19),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_122),
.B(n_125),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_78),
.B(n_80),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_126),
.A2(n_133),
.B1(n_70),
.B2(n_8),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_58),
.B(n_42),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_2),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_129),
.B(n_6),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_53),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_55),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_133)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_134),
.Y(n_184)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_135),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_67),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_136),
.B(n_145),
.Y(n_190)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_137),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g213 ( 
.A1(n_138),
.A2(n_148),
.B1(n_153),
.B2(n_172),
.Y(n_213)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_139),
.Y(n_183)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_140),
.Y(n_218)
);

AND2x2_ASAP7_75t_SL g201 ( 
.A(n_141),
.B(n_118),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_113),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_142),
.B(n_156),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_144),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_98),
.Y(n_145)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_149),
.Y(n_208)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_105),
.Y(n_150)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_150),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_100),
.A2(n_54),
.B1(n_10),
.B2(n_11),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_151),
.A2(n_160),
.B1(n_170),
.B2(n_171),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_131),
.A2(n_6),
.B1(n_10),
.B2(n_11),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_152),
.A2(n_159),
.B1(n_164),
.B2(n_165),
.Y(n_193)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_153),
.Y(n_194)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_88),
.Y(n_154)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_154),
.Y(n_199)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_110),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_157),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_95),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_169),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_101),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_92),
.A2(n_12),
.B1(n_13),
.B2(n_97),
.Y(n_160)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_106),
.Y(n_162)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_162),
.Y(n_220)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_106),
.Y(n_163)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_103),
.B1(n_111),
.B2(n_115),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_122),
.A2(n_126),
.B1(n_102),
.B2(n_125),
.Y(n_165)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_109),
.Y(n_166)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_166),
.Y(n_212)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_89),
.Y(n_167)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_167),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_130),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_98),
.A2(n_86),
.B1(n_108),
.B2(n_128),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_116),
.Y(n_171)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_171),
.Y(n_219)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_89),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_175),
.Y(n_179)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_109),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_174),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_86),
.B(n_120),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_120),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_108),
.A2(n_87),
.B1(n_117),
.B2(n_127),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_177),
.A2(n_112),
.B1(n_132),
.B2(n_88),
.Y(n_182)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_117),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_119),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_147),
.A2(n_87),
.B1(n_128),
.B2(n_104),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_180),
.A2(n_182),
.B1(n_188),
.B2(n_214),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_185),
.B(n_212),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_168),
.B(n_119),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_186),
.B(n_197),
.C(n_206),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_142),
.A2(n_112),
.B1(n_96),
.B2(n_88),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_155),
.A2(n_133),
.B1(n_132),
.B2(n_123),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_191),
.A2(n_198),
.B1(n_200),
.B2(n_197),
.Y(n_249)
);

AO21x2_ASAP7_75t_SL g192 ( 
.A1(n_146),
.A2(n_123),
.B(n_96),
.Y(n_192)
);

AOI22x1_ASAP7_75t_L g231 ( 
.A1(n_192),
.A2(n_162),
.B1(n_163),
.B2(n_157),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_132),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_175),
.A2(n_138),
.B1(n_176),
.B2(n_161),
.Y(n_198)
);

AO21x2_ASAP7_75t_L g200 ( 
.A1(n_146),
.A2(n_94),
.B(n_118),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_201),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_94),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_205),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_110),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_141),
.B(n_174),
.C(n_167),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_178),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_215),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_218),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_141),
.A2(n_148),
.B1(n_140),
.B2(n_139),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_149),
.B(n_150),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_221),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_144),
.B(n_134),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_214),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_222),
.B(n_250),
.Y(n_268)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_183),
.Y(n_225)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_225),
.Y(n_264)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_226),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_198),
.A2(n_154),
.B1(n_173),
.B2(n_137),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_228),
.A2(n_249),
.B1(n_252),
.B2(n_255),
.Y(n_293)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_183),
.Y(n_229)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_229),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_190),
.B(n_135),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_230),
.B(n_244),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_231),
.Y(n_273)
);

INVxp33_ASAP7_75t_L g233 ( 
.A(n_192),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_233),
.Y(n_269)
);

XNOR2x2_ASAP7_75t_SL g263 ( 
.A(n_234),
.B(n_257),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_209),
.A2(n_166),
.B(n_196),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_235),
.A2(n_236),
.B(n_256),
.Y(n_271)
);

A2O1A1O1Ixp25_ASAP7_75t_L g236 ( 
.A1(n_206),
.A2(n_186),
.B(n_203),
.C(n_205),
.D(n_179),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_208),
.Y(n_237)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_237),
.Y(n_272)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_238),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_195),
.Y(n_239)
);

INVx13_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_185),
.Y(n_240)
);

INVx4_ASAP7_75t_SL g277 ( 
.A(n_240),
.Y(n_277)
);

INVxp33_ASAP7_75t_L g242 ( 
.A(n_192),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_242),
.B(n_247),
.Y(n_282)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_208),
.Y(n_243)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_243),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_179),
.B(n_194),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_194),
.B(n_217),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_253),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_200),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_246),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_192),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_219),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_220),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_251),
.B(n_258),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_191),
.A2(n_180),
.B1(n_213),
.B2(n_201),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_201),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_202),
.Y(n_254)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_254),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_193),
.A2(n_200),
.B1(n_213),
.B2(n_187),
.Y(n_255)
);

NAND5xp2_ASAP7_75t_L g256 ( 
.A(n_200),
.B(n_207),
.C(n_187),
.D(n_204),
.E(n_184),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_204),
.B(n_199),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_181),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_259),
.B(n_181),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_211),
.C(n_189),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_260),
.B(n_227),
.C(n_245),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_257),
.Y(n_261)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_261),
.Y(n_302)
);

INVxp33_ASAP7_75t_SL g262 ( 
.A(n_223),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_262),
.B(n_281),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_230),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_280),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_258),
.Y(n_267)
);

INVxp67_ASAP7_75t_SL g317 ( 
.A(n_267),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_248),
.B(n_200),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_276),
.B(n_278),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_232),
.B(n_211),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_239),
.B(n_235),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_234),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_253),
.A2(n_184),
.B(n_199),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_286),
.Y(n_322)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_225),
.Y(n_288)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_288),
.Y(n_304)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_289),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_240),
.B(n_189),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_291),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_232),
.A2(n_222),
.B1(n_247),
.B2(n_241),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_292),
.A2(n_249),
.B1(n_252),
.B2(n_244),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_246),
.A2(n_255),
.B1(n_227),
.B2(n_224),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_294),
.A2(n_229),
.B1(n_226),
.B2(n_238),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_297),
.B(n_312),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_231),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_300),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_282),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_301),
.B(n_303),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_266),
.Y(n_303)
);

OAI21x1_ASAP7_75t_R g305 ( 
.A1(n_269),
.A2(n_256),
.B(n_231),
.Y(n_305)
);

A2O1A1Ixp33_ASAP7_75t_SL g345 ( 
.A1(n_305),
.A2(n_319),
.B(n_263),
.C(n_277),
.Y(n_345)
);

XNOR2x1_ASAP7_75t_SL g306 ( 
.A(n_274),
.B(n_236),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_306),
.B(n_271),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_307),
.B(n_315),
.C(n_271),
.Y(n_332)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_264),
.Y(n_308)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_308),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_292),
.A2(n_256),
.B1(n_224),
.B2(n_241),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_309),
.A2(n_293),
.B1(n_281),
.B2(n_286),
.Y(n_349)
);

HB1xp67_ASAP7_75t_SL g311 ( 
.A(n_276),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_311),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g312 ( 
.A(n_287),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_264),
.Y(n_313)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_313),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_273),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_260),
.B(n_228),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_287),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_316),
.B(n_277),
.Y(n_348)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_270),
.Y(n_318)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_318),
.Y(n_337)
);

OA21x2_ASAP7_75t_L g319 ( 
.A1(n_274),
.A2(n_237),
.B(n_243),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_270),
.Y(n_320)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_320),
.Y(n_340)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_288),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_321),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_266),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_323),
.B(n_277),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_319),
.Y(n_324)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_324),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_327),
.A2(n_322),
.B1(n_305),
.B2(n_342),
.Y(n_356)
);

CKINVDCx14_ASAP7_75t_R g369 ( 
.A(n_330),
.Y(n_369)
);

INVx13_ASAP7_75t_L g331 ( 
.A(n_305),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_331),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_332),
.B(n_307),
.C(n_310),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_296),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_334),
.B(n_341),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_295),
.B(n_279),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_335),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_336),
.B(n_309),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_312),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_338),
.B(n_344),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_298),
.B(n_285),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_296),
.B(n_285),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_343),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_299),
.B(n_267),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_345),
.B(n_348),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_299),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_346),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_315),
.B(n_268),
.Y(n_347)
);

NOR2xp67_ASAP7_75t_SL g352 ( 
.A(n_347),
.B(n_297),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_349),
.A2(n_293),
.B1(n_300),
.B2(n_273),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_350),
.B(n_363),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_332),
.B(n_310),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_351),
.B(n_345),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_369),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_336),
.B(n_306),
.C(n_317),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_355),
.B(n_361),
.C(n_329),
.Y(n_378)
);

XNOR2x1_ASAP7_75t_L g385 ( 
.A(n_356),
.B(n_358),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_342),
.A2(n_322),
.B(n_302),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_359),
.A2(n_365),
.B(n_324),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_326),
.B(n_278),
.C(n_319),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_349),
.B(n_263),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_339),
.A2(n_300),
.B(n_269),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_367),
.A2(n_327),
.B1(n_339),
.B2(n_338),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_345),
.A2(n_261),
.B(n_316),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_370),
.A2(n_348),
.B(n_327),
.Y(n_373)
);

OR2x2_ASAP7_75t_L g398 ( 
.A(n_371),
.B(n_373),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_360),
.B(n_335),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_372),
.B(n_381),
.Y(n_392)
);

OAI211xp5_ASAP7_75t_L g388 ( 
.A1(n_375),
.A2(n_357),
.B(n_370),
.C(n_368),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_376),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_360),
.A2(n_328),
.B1(n_334),
.B2(n_344),
.Y(n_377)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_377),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_378),
.B(n_380),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_379),
.B(n_382),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_361),
.B(n_329),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_366),
.B(n_304),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_355),
.B(n_345),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_358),
.B(n_345),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_383),
.B(n_384),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_364),
.B(n_362),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_350),
.B(n_272),
.C(n_283),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_386),
.B(n_387),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_357),
.Y(n_387)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_388),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_386),
.B(n_351),
.C(n_362),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_389),
.B(n_395),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_371),
.A2(n_368),
.B(n_359),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_390),
.A2(n_331),
.B(n_312),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_374),
.B(n_363),
.C(n_356),
.Y(n_395)
);

AOI321xp33_ASAP7_75t_L g399 ( 
.A1(n_374),
.A2(n_353),
.A3(n_325),
.B1(n_337),
.B2(n_340),
.C(n_333),
.Y(n_399)
);

BUFx24_ASAP7_75t_SL g404 ( 
.A(n_399),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_400),
.B(n_380),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_401),
.B(n_405),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_397),
.A2(n_354),
.B1(n_385),
.B2(n_382),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_402),
.B(n_316),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_391),
.A2(n_367),
.B1(n_340),
.B2(n_337),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_398),
.A2(n_383),
.B(n_379),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_406),
.A2(n_411),
.B(n_402),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_389),
.B(n_378),
.C(n_385),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_407),
.B(n_408),
.C(n_393),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_397),
.A2(n_365),
.B1(n_333),
.B2(n_325),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_392),
.B(n_254),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_410),
.B(n_412),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_396),
.B(n_308),
.Y(n_412)
);

AOI322xp5_ASAP7_75t_L g413 ( 
.A1(n_409),
.A2(n_394),
.A3(n_398),
.B1(n_393),
.B2(n_395),
.C1(n_318),
.C2(n_313),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_413),
.B(n_420),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_401),
.B(n_321),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_415),
.B(n_417),
.Y(n_425)
);

OAI21x1_ASAP7_75t_L g428 ( 
.A1(n_418),
.A2(n_419),
.B(n_284),
.Y(n_428)
);

MAJx2_ASAP7_75t_L g420 ( 
.A(n_403),
.B(n_407),
.C(n_404),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_406),
.B(n_272),
.C(n_283),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_421),
.B(n_275),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_416),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_422),
.B(n_424),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_414),
.B(n_419),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_426),
.B(n_428),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_413),
.A2(n_320),
.B(n_284),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_427),
.B(n_275),
.C(n_259),
.Y(n_429)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_429),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_425),
.B(n_275),
.Y(n_432)
);

AO21x1_ASAP7_75t_L g433 ( 
.A1(n_432),
.A2(n_423),
.B(n_431),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_433),
.B(n_430),
.C(n_423),
.Y(n_435)
);

BUFx24_ASAP7_75t_SL g436 ( 
.A(n_435),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_436),
.B(n_434),
.Y(n_437)
);


endmodule