module real_jpeg_14044_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_285, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_285;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_243;
wire n_105;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_200;
wire n_164;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_211;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_244;
wire n_202;
wire n_128;
wire n_179;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_273;
wire n_253;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_0),
.A2(n_23),
.B1(n_26),
.B2(n_36),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_0),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_0),
.A2(n_36),
.B1(n_45),
.B2(n_46),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_0),
.A2(n_8),
.B(n_32),
.C(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_0),
.A2(n_36),
.B1(n_56),
.B2(n_57),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_0),
.B(n_37),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_0),
.B(n_54),
.C(n_57),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_0),
.B(n_44),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_0),
.B(n_29),
.C(n_33),
.Y(n_167)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_3),
.Y(n_100)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_40),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_6),
.A2(n_23),
.B1(n_26),
.B2(n_40),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_6),
.A2(n_40),
.B1(n_56),
.B2(n_57),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_6),
.A2(n_40),
.B1(n_45),
.B2(n_46),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

AO22x1_ASAP7_75t_L g44 ( 
.A1(n_8),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

INVxp33_ASAP7_75t_L g282 ( 
.A(n_9),
.Y(n_282)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_11),
.A2(n_23),
.B1(n_26),
.B2(n_48),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_11),
.A2(n_48),
.B1(n_56),
.B2(n_57),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_12),
.A2(n_15),
.B(n_281),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_12),
.B(n_282),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_13),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_13),
.A2(n_25),
.B1(n_32),
.B2(n_33),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_13),
.A2(n_25),
.B1(n_45),
.B2(n_46),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_13),
.A2(n_25),
.B1(n_56),
.B2(n_57),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_74),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_72),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_69),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_18),
.B(n_69),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_62),
.C(n_66),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_19),
.B(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_38),
.C(n_49),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_20),
.A2(n_107),
.B1(n_117),
.B2(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_20),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_20),
.B(n_117),
.C(n_180),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_20),
.A2(n_83),
.B1(n_84),
.B2(n_182),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_20),
.A2(n_182),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_27),
.B1(n_35),
.B2(n_37),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OA21x2_ASAP7_75t_L g170 ( 
.A1(n_22),
.A2(n_31),
.B(n_68),
.Y(n_170)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_26),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_27),
.B(n_35),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_27),
.B(n_37),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_29),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_31),
.A2(n_67),
.B(n_68),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_31),
.A2(n_67),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_42),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

INVxp33_ASAP7_75t_L g238 ( 
.A(n_35),
.Y(n_238)
);

OAI21xp33_ASAP7_75t_SL g96 ( 
.A1(n_36),
.A2(n_42),
.B(n_45),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_36),
.B(n_103),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_36),
.B(n_60),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_38),
.A2(n_49),
.B1(n_256),
.B2(n_270),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_38),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_41),
.B1(n_44),
.B2(n_47),
.Y(n_38)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_39),
.Y(n_258)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_41),
.B(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_46),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_46),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_49),
.A2(n_256),
.B1(n_257),
.B2(n_259),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_49),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_49),
.B(n_170),
.C(n_257),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_60),
.B(n_61),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_50),
.A2(n_60),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_92),
.Y(n_91)
);

AO22x1_ASAP7_75t_SL g122 ( 
.A1(n_51),
.A2(n_55),
.B1(n_90),
.B2(n_92),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_51),
.A2(n_55),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

NOR2x1_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

AO22x1_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_56),
.B(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_57),
.B(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OA21x2_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_89),
.B(n_91),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_60),
.A2(n_91),
.B(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_61),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_62),
.B(n_66),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_64),
.A2(n_65),
.B1(n_85),
.B2(n_108),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_64),
.A2(n_65),
.B(n_108),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_85),
.B(n_86),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_65),
.A2(n_86),
.B(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_276),
.B(n_280),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_248),
.B(n_273),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_226),
.B(n_247),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_209),
.B(n_225),
.Y(n_77)
);

OAI321xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_177),
.A3(n_204),
.B1(n_207),
.B2(n_208),
.C(n_285),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_159),
.B(n_176),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_125),
.B(n_158),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_104),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_82),
.B(n_104),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_88),
.C(n_93),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_83),
.A2(n_84),
.B1(n_88),
.B2(n_142),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_83),
.A2(n_84),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_84),
.B(n_169),
.C(n_174),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_84),
.B(n_182),
.C(n_214),
.Y(n_246)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_88),
.B(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_88),
.A2(n_129),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_88),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_88),
.A2(n_142),
.B1(n_184),
.B2(n_186),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_92),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_93),
.A2(n_94),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_97),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_98),
.A2(n_102),
.B1(n_103),
.B2(n_114),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_99),
.B(n_202),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_102),
.A2(n_103),
.B1(n_185),
.B2(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_114),
.B(n_115),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_103),
.A2(n_115),
.B(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_119),
.B2(n_120),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_105),
.B(n_122),
.C(n_123),
.Y(n_160)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_109),
.B1(n_117),
.B2(n_118),
.Y(n_106)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_107),
.B(n_110),
.C(n_113),
.Y(n_163)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_112),
.B(n_140),
.Y(n_150)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_113),
.B(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_117),
.A2(n_242),
.B(n_245),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_117),
.B(n_242),
.Y(n_245)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_121),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_122),
.A2(n_124),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_134),
.C(n_136),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_122),
.A2(n_124),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_122),
.B(n_201),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_152),
.B(n_157),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_138),
.B(n_151),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_131),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_128),
.B(n_131),
.Y(n_151)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_131)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_133),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_136),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_136),
.B(n_148),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_136),
.B(n_165),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_143),
.B(n_150),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_142),
.B(n_184),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_147),
.B(n_149),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_153),
.B(n_154),
.Y(n_157)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_160),
.B(n_161),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_168),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_163),
.B(n_164),
.C(n_168),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_169),
.A2(n_170),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_169),
.B(n_192),
.C(n_197),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_169),
.A2(n_170),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_169),
.A2(n_170),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_170),
.B(n_267),
.C(n_271),
.Y(n_279)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_188),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_188),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.C(n_187),
.Y(n_178)
);

FAx1_ASAP7_75t_SL g206 ( 
.A(n_179),
.B(n_183),
.CI(n_187),
.CON(n_206),
.SN(n_206)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_184),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_203),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_198),
.B2(n_199),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_199),
.C(n_203),
.Y(n_224)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_205),
.B(n_206),
.Y(n_207)
);

BUFx24_ASAP7_75t_SL g284 ( 
.A(n_206),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_224),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_224),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_213),
.C(n_218),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_218),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_223),
.Y(n_218)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_219),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_221),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_219),
.A2(n_223),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_223),
.A2(n_232),
.B(n_237),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_228),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_246),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_240),
.B2(n_241),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_240),
.C(n_246),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_245),
.A2(n_252),
.B1(n_253),
.B2(n_260),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_245),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_263),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_262),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_262),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_261),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_260),
.C(n_261),
.Y(n_272)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_257),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_263),
.A2(n_274),
.B(n_275),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_272),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_272),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_271),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_279),
.Y(n_280)
);


endmodule