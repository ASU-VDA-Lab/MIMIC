module fake_jpeg_27371_n_309 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_309);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_309;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_44),
.B(n_46),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_26),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_18),
.B1(n_19),
.B2(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_29),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_26),
.Y(n_56)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_31),
.Y(n_59)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_26),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_64),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_33),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_49),
.A2(n_25),
.B1(n_31),
.B2(n_24),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_74),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_36),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_84),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_49),
.A2(n_25),
.B1(n_24),
.B2(n_33),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_90),
.B1(n_55),
.B2(n_37),
.Y(n_93)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_82),
.Y(n_95)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_36),
.Y(n_84)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

AO22x2_ASAP7_75t_SL g90 ( 
.A1(n_58),
.A2(n_41),
.B1(n_37),
.B2(n_34),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_90),
.A2(n_53),
.B1(n_47),
.B2(n_55),
.Y(n_113)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_93),
.A2(n_88),
.B1(n_91),
.B2(n_67),
.Y(n_137)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_98),
.B(n_100),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_78),
.B(n_27),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_111),
.C(n_118),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_103),
.A2(n_113),
.B1(n_71),
.B2(n_80),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_109),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_24),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_108),
.B(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_41),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_76),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_43),
.C(n_39),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_116),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_72),
.B(n_19),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_27),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_43),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_53),
.B1(n_32),
.B2(n_17),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_118),
.A2(n_88),
.B1(n_82),
.B2(n_77),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_106),
.B(n_103),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_132),
.B(n_140),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g121 ( 
.A(n_108),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_121),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_122),
.B(n_62),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_113),
.A2(n_18),
.B1(n_19),
.B2(n_22),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_124),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_126),
.A2(n_104),
.B1(n_86),
.B2(n_17),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_99),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_127),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_128),
.A2(n_137),
.B1(n_32),
.B2(n_22),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_131),
.B(n_134),
.Y(n_157)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_98),
.B(n_71),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_135),
.Y(n_147)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

O2A1O1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_109),
.A2(n_47),
.B(n_77),
.C(n_75),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_139),
.Y(n_161)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

OA21x2_ASAP7_75t_L g140 ( 
.A1(n_97),
.A2(n_40),
.B(n_51),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_94),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_141),
.Y(n_160)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_144),
.Y(n_164)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_102),
.C(n_100),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_146),
.B(n_148),
.C(n_149),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_96),
.C(n_105),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_96),
.C(n_105),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_103),
.B(n_94),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_151),
.A2(n_170),
.B(n_22),
.Y(n_179)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_166),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_117),
.C(n_115),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_154),
.B(n_163),
.C(n_120),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_27),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_163),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_156),
.A2(n_158),
.B1(n_129),
.B2(n_141),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_128),
.A2(n_104),
.B1(n_86),
.B2(n_17),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_136),
.A2(n_17),
.B1(n_32),
.B2(n_22),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_159),
.A2(n_129),
.B1(n_135),
.B2(n_142),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_165),
.A2(n_152),
.B1(n_166),
.B2(n_150),
.Y(n_196)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_125),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_167),
.B(n_168),
.Y(n_182)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_127),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_169),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_140),
.A2(n_0),
.B(n_1),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_175),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

AO22x2_ASAP7_75t_L g174 ( 
.A1(n_145),
.A2(n_140),
.B1(n_124),
.B2(n_126),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_174),
.A2(n_183),
.B1(n_172),
.B2(n_193),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_164),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_176),
.A2(n_183),
.B1(n_193),
.B2(n_196),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_131),
.Y(n_177)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_177),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_178),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_179),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_L g180 ( 
.A1(n_151),
.A2(n_138),
.B(n_121),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_192),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_187),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_145),
.A2(n_161),
.B(n_170),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_132),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_62),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_171),
.B(n_138),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_189),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_161),
.A2(n_132),
.B(n_144),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_191),
.A2(n_169),
.B1(n_162),
.B2(n_150),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_171),
.B(n_132),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_168),
.A2(n_120),
.B1(n_32),
.B2(n_28),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_155),
.Y(n_200)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_147),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_20),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_146),
.C(n_154),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_200),
.C(n_202),
.Y(n_225)
);

NAND2xp33_ASAP7_75t_SL g201 ( 
.A(n_174),
.B(n_152),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_201),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_153),
.C(n_157),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_204),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_158),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_188),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_162),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_207),
.A2(n_0),
.B(n_33),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_174),
.A2(n_156),
.B1(n_159),
.B2(n_18),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_174),
.A2(n_28),
.B1(n_30),
.B2(n_29),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_216),
.B(n_185),
.Y(n_224)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_218),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_185),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_191),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_43),
.C(n_62),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_195),
.C(n_181),
.Y(n_228)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_221),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_229),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_208),
.A2(n_187),
.B(n_179),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_223),
.Y(n_245)
);

MAJx2_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_202),
.C(n_220),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_197),
.B(n_184),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_226),
.B(n_235),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_234),
.C(n_224),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_178),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_219),
.Y(n_230)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_230),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_231),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_28),
.B1(n_30),
.B2(n_29),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_232),
.A2(n_238),
.B1(n_212),
.B2(n_16),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_199),
.B(n_43),
.C(n_23),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_20),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_217),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_237),
.B(n_239),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_206),
.A2(n_30),
.B1(n_23),
.B2(n_20),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_215),
.B(n_2),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_209),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_240),
.B(n_205),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_242),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_243),
.A2(n_254),
.B1(n_20),
.B2(n_27),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_251),
.C(n_255),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_238),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_216),
.C(n_203),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_227),
.A2(n_211),
.B1(n_213),
.B2(n_210),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_234),
.C(n_229),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_203),
.C(n_23),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_23),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_252),
.A2(n_236),
.B1(n_233),
.B2(n_223),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_257),
.A2(n_265),
.B1(n_21),
.B2(n_4),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_255),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_232),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_260),
.B(n_264),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_247),
.B(n_2),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_270),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_233),
.Y(n_263)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_244),
.A2(n_20),
.B1(n_23),
.B2(n_5),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_267),
.A2(n_21),
.B1(n_6),
.B2(n_7),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_3),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_269),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_241),
.B(n_251),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_253),
.B(n_3),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_245),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_273),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_266),
.A2(n_250),
.B(n_246),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_281),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_21),
.C(n_4),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_279),
.C(n_257),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_282),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_21),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_3),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_262),
.Y(n_283)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_283),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_286),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_272),
.A2(n_4),
.B(n_6),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_288),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_7),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_276),
.B(n_275),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_291),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_8),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_279),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_295),
.A2(n_10),
.B(n_12),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_284),
.B(n_276),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_298),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_8),
.Y(n_298)
);

A2O1A1O1Ixp25_ASAP7_75t_L g299 ( 
.A1(n_292),
.A2(n_285),
.B(n_11),
.C(n_12),
.D(n_13),
.Y(n_299)
);

AOI221xp5_ASAP7_75t_SL g303 ( 
.A1(n_299),
.A2(n_301),
.B1(n_302),
.B2(n_300),
.C(n_13),
.Y(n_303)
);

AO21x1_ASAP7_75t_L g302 ( 
.A1(n_295),
.A2(n_10),
.B(n_13),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_303),
.B(n_304),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_293),
.C(n_297),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_294),
.C(n_14),
.Y(n_306)
);

NAND3xp33_ASAP7_75t_SL g307 ( 
.A(n_306),
.B(n_10),
.C(n_14),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_15),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_15),
.Y(n_309)
);


endmodule