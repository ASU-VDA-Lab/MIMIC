module real_aes_16030_n_297 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_286, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_287, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_293, n_124, n_22, n_173, n_191, n_209, n_296, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_288, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_295, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_294, n_227, n_67, n_92, n_33, n_206, n_258, n_291, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_292, n_116, n_94, n_229, n_289, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_290, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_297);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_286;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_287;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_293;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_296;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_288;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_295;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_294;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_291;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_292;
input n_116;
input n_94;
input n_229;
input n_289;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_290;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_297;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_1487;
wire n_939;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_334;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_1524;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1175;
wire n_778;
wire n_1170;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_1268;
wire n_852;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1496;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_1049;
wire n_559;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1252;
wire n_430;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1280;
wire n_394;
wire n_729;
wire n_1352;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp5_ASAP7_75t_L g1314 ( .A1(n_0), .A2(n_224), .B1(n_1287), .B2(n_1291), .Y(n_1314) );
OAI22xp33_ASAP7_75t_SL g698 ( .A1(n_1), .A2(n_133), .B1(n_445), .B2(n_448), .Y(n_698) );
OAI22xp33_ASAP7_75t_L g709 ( .A1(n_1), .A2(n_22), .B1(n_458), .B2(n_459), .Y(n_709) );
INVx1_ASAP7_75t_L g906 ( .A(n_2), .Y(n_906) );
INVx1_ASAP7_75t_L g1268 ( .A(n_3), .Y(n_1268) );
OAI22xp5_ASAP7_75t_L g1111 ( .A1(n_4), .A2(n_204), .B1(n_841), .B2(n_1112), .Y(n_1111) );
INVxp67_ASAP7_75t_SL g1129 ( .A(n_4), .Y(n_1129) );
AOI22xp33_ASAP7_75t_L g1323 ( .A1(n_5), .A2(n_54), .B1(n_1287), .B2(n_1291), .Y(n_1323) );
OAI22xp33_ASAP7_75t_L g1217 ( .A1(n_6), .A2(n_193), .B1(n_439), .B2(n_448), .Y(n_1217) );
OAI22xp33_ASAP7_75t_SL g1227 ( .A1(n_6), .A2(n_193), .B1(n_458), .B2(n_548), .Y(n_1227) );
OAI211xp5_ASAP7_75t_L g1494 ( .A1(n_7), .A2(n_422), .B(n_963), .C(n_1495), .Y(n_1494) );
INVx1_ASAP7_75t_L g1504 ( .A(n_7), .Y(n_1504) );
INVx1_ASAP7_75t_L g576 ( .A(n_8), .Y(n_576) );
INVx1_ASAP7_75t_L g1252 ( .A(n_9), .Y(n_1252) );
INVx1_ASAP7_75t_L g1044 ( .A(n_10), .Y(n_1044) );
INVx1_ASAP7_75t_L g312 ( .A(n_11), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_11), .B(n_322), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g681 ( .A(n_12), .Y(n_681) );
OAI22xp33_ASAP7_75t_L g832 ( .A1(n_13), .A2(n_236), .B1(n_314), .B2(n_544), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g850 ( .A1(n_13), .A2(n_236), .B1(n_851), .B2(n_853), .Y(n_850) );
CKINVDCx5p33_ASAP7_75t_R g671 ( .A(n_14), .Y(n_671) );
CKINVDCx5p33_ASAP7_75t_R g675 ( .A(n_15), .Y(n_675) );
INVx1_ASAP7_75t_L g955 ( .A(n_16), .Y(n_955) );
INVx1_ASAP7_75t_L g1509 ( .A(n_17), .Y(n_1509) );
INVx1_ASAP7_75t_L g739 ( .A(n_18), .Y(n_739) );
INVx2_ASAP7_75t_L g1290 ( .A(n_19), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_19), .B(n_112), .Y(n_1292) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_19), .B(n_1296), .Y(n_1298) );
AOI22xp33_ASAP7_75t_SL g611 ( .A1(n_20), .A2(n_284), .B1(n_593), .B2(n_596), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_20), .A2(n_23), .B1(n_621), .B2(n_626), .Y(n_636) );
INVx1_ASAP7_75t_L g647 ( .A(n_21), .Y(n_647) );
OAI22xp33_ASAP7_75t_SL g695 ( .A1(n_22), .A2(n_268), .B1(n_439), .B2(n_696), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_23), .A2(n_198), .B1(n_599), .B2(n_604), .Y(n_598) );
AO22x2_ASAP7_75t_L g1189 ( .A1(n_24), .A2(n_1190), .B1(n_1233), .B2(n_1234), .Y(n_1189) );
INVx1_ASAP7_75t_L g1233 ( .A(n_24), .Y(n_1233) );
AOI22xp5_ASAP7_75t_L g1308 ( .A1(n_24), .A2(n_33), .B1(n_1294), .B2(n_1297), .Y(n_1308) );
OAI22xp33_ASAP7_75t_L g1269 ( .A1(n_25), .A2(n_248), .B1(n_458), .B2(n_1151), .Y(n_1269) );
OAI22xp33_ASAP7_75t_L g1278 ( .A1(n_25), .A2(n_290), .B1(n_439), .B2(n_544), .Y(n_1278) );
INVx1_ASAP7_75t_L g573 ( .A(n_26), .Y(n_573) );
OAI22xp33_ASAP7_75t_L g521 ( .A1(n_27), .A2(n_170), .B1(n_448), .B2(n_522), .Y(n_521) );
OAI22xp33_ASAP7_75t_L g524 ( .A1(n_27), .A2(n_286), .B1(n_458), .B2(n_459), .Y(n_524) );
XOR2xp5_ASAP7_75t_L g666 ( .A(n_28), .B(n_667), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g1313 ( .A1(n_28), .A2(n_132), .B1(n_1294), .B2(n_1297), .Y(n_1313) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_29), .A2(n_188), .B1(n_314), .B2(n_448), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_29), .A2(n_188), .B1(n_459), .B2(n_651), .Y(n_650) );
CKINVDCx5p33_ASAP7_75t_R g497 ( .A(n_30), .Y(n_497) );
OAI22xp33_ASAP7_75t_L g543 ( .A1(n_31), .A2(n_156), .B1(n_439), .B2(n_544), .Y(n_543) );
OAI22xp33_ASAP7_75t_SL g547 ( .A1(n_31), .A2(n_156), .B1(n_458), .B2(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g1195 ( .A(n_32), .Y(n_1195) );
OAI22xp33_ASAP7_75t_L g438 ( .A1(n_34), .A2(n_222), .B1(n_439), .B2(n_441), .Y(n_438) );
OAI22xp33_ASAP7_75t_L g457 ( .A1(n_34), .A2(n_106), .B1(n_458), .B2(n_459), .Y(n_457) );
CKINVDCx5p33_ASAP7_75t_R g679 ( .A(n_35), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g1372 ( .A1(n_36), .A2(n_111), .B1(n_1287), .B2(n_1373), .Y(n_1372) );
INVx1_ASAP7_75t_L g897 ( .A(n_37), .Y(n_897) );
AOI22xp5_ASAP7_75t_L g1300 ( .A1(n_38), .A2(n_104), .B1(n_1287), .B2(n_1301), .Y(n_1300) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_39), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g1020 ( .A(n_40), .Y(n_1020) );
CKINVDCx5p33_ASAP7_75t_R g494 ( .A(n_41), .Y(n_494) );
XOR2x2_ASAP7_75t_L g927 ( .A(n_42), .B(n_928), .Y(n_927) );
XOR2x2_ASAP7_75t_L g588 ( .A(n_43), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g1091 ( .A(n_44), .Y(n_1091) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_45), .A2(n_197), .B1(n_459), .B2(n_480), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_45), .A2(n_47), .B1(n_522), .B2(n_542), .Y(n_748) );
INVx1_ASAP7_75t_L g642 ( .A(n_46), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_47), .A2(n_293), .B1(n_458), .B2(n_479), .Y(n_732) );
INVx1_ASAP7_75t_L g1093 ( .A(n_48), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_48), .A2(n_88), .B1(n_610), .B2(n_1121), .Y(n_1126) );
OAI22xp33_ASAP7_75t_L g1493 ( .A1(n_49), .A2(n_137), .B1(n_522), .B2(n_542), .Y(n_1493) );
OAI22xp33_ASAP7_75t_L g1505 ( .A1(n_49), .A2(n_59), .B1(n_459), .B2(n_480), .Y(n_1505) );
INVx1_ASAP7_75t_L g540 ( .A(n_50), .Y(n_540) );
INVx1_ASAP7_75t_L g347 ( .A(n_51), .Y(n_347) );
INVx1_ASAP7_75t_L g354 ( .A(n_51), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g871 ( .A1(n_52), .A2(n_151), .B1(n_851), .B2(n_872), .Y(n_871) );
OAI22xp33_ASAP7_75t_L g890 ( .A1(n_52), .A2(n_151), .B1(n_314), .B2(n_448), .Y(n_890) );
AOI22xp5_ASAP7_75t_L g1319 ( .A1(n_53), .A2(n_142), .B1(n_1287), .B2(n_1301), .Y(n_1319) );
XOR2xp5_ASAP7_75t_L g1238 ( .A(n_55), .B(n_1239), .Y(n_1238) );
INVx1_ASAP7_75t_L g813 ( .A(n_56), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g1374 ( .A1(n_57), .A2(n_250), .B1(n_1294), .B2(n_1297), .Y(n_1374) );
OAI22xp33_ASAP7_75t_L g1224 ( .A1(n_58), .A2(n_116), .B1(n_522), .B2(n_1225), .Y(n_1224) );
OAI22xp33_ASAP7_75t_L g1232 ( .A1(n_58), .A2(n_116), .B1(n_479), .B2(n_480), .Y(n_1232) );
OAI22xp33_ASAP7_75t_L g1498 ( .A1(n_59), .A2(n_230), .B1(n_439), .B2(n_544), .Y(n_1498) );
INVx1_ASAP7_75t_L g797 ( .A(n_60), .Y(n_797) );
INVx1_ASAP7_75t_L g1060 ( .A(n_61), .Y(n_1060) );
OAI211xp5_ASAP7_75t_L g420 ( .A1(n_62), .A2(n_421), .B(n_422), .C(n_428), .Y(n_420) );
INVx1_ASAP7_75t_L g477 ( .A(n_62), .Y(n_477) );
INVx1_ASAP7_75t_L g305 ( .A(n_63), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g994 ( .A1(n_64), .A2(n_179), .B1(n_887), .B2(n_936), .Y(n_994) );
OAI22xp5_ASAP7_75t_L g997 ( .A1(n_64), .A2(n_179), .B1(n_862), .B2(n_863), .Y(n_997) );
INVx2_ASAP7_75t_L g340 ( .A(n_65), .Y(n_340) );
XNOR2x2_ASAP7_75t_L g785 ( .A(n_66), .B(n_786), .Y(n_785) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_67), .A2(n_271), .B1(n_655), .B2(n_715), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_67), .A2(n_202), .B1(n_766), .B2(n_768), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g845 ( .A1(n_68), .A2(n_252), .B1(n_846), .B2(n_847), .Y(n_845) );
OAI22xp33_ASAP7_75t_L g861 ( .A1(n_68), .A2(n_252), .B1(n_862), .B2(n_863), .Y(n_861) );
INVx1_ASAP7_75t_L g1101 ( .A(n_69), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g1163 ( .A1(n_70), .A2(n_220), .B1(n_1157), .B2(n_1164), .Y(n_1163) );
AOI22xp33_ASAP7_75t_L g1181 ( .A1(n_70), .A2(n_234), .B1(n_1175), .B2(n_1179), .Y(n_1181) );
INVx1_ASAP7_75t_L g1245 ( .A(n_71), .Y(n_1245) );
INVx1_ASAP7_75t_L g738 ( .A(n_72), .Y(n_738) );
INVx1_ASAP7_75t_L g1497 ( .A(n_73), .Y(n_1497) );
INVx1_ASAP7_75t_L g735 ( .A(n_74), .Y(n_735) );
XNOR2xp5_ASAP7_75t_L g1081 ( .A(n_75), .B(n_1082), .Y(n_1081) );
INVx1_ASAP7_75t_L g799 ( .A(n_76), .Y(n_799) );
OAI222xp33_ASAP7_75t_L g1152 ( .A1(n_77), .A2(n_118), .B1(n_266), .B2(n_702), .C1(n_1131), .C2(n_1153), .Y(n_1152) );
OAI222xp33_ASAP7_75t_L g1188 ( .A1(n_77), .A2(n_118), .B1(n_266), .B2(n_841), .C1(n_963), .C2(n_1112), .Y(n_1188) );
INVx1_ASAP7_75t_L g1512 ( .A(n_78), .Y(n_1512) );
OAI22xp33_ASAP7_75t_L g444 ( .A1(n_79), .A2(n_106), .B1(n_445), .B2(n_448), .Y(n_444) );
OAI22xp33_ASAP7_75t_L g478 ( .A1(n_79), .A2(n_222), .B1(n_479), .B2(n_480), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g1071 ( .A1(n_80), .A2(n_259), .B1(n_887), .B2(n_936), .Y(n_1071) );
OAI22xp33_ASAP7_75t_L g1080 ( .A1(n_80), .A2(n_259), .B1(n_862), .B2(n_939), .Y(n_1080) );
INVx1_ASAP7_75t_L g564 ( .A(n_81), .Y(n_564) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_82), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g1159 ( .A1(n_83), .A2(n_294), .B1(n_1160), .B2(n_1162), .Y(n_1159) );
AOI22xp33_ASAP7_75t_SL g1182 ( .A1(n_83), .A2(n_150), .B1(n_772), .B2(n_1183), .Y(n_1182) );
OAI22xp33_ASAP7_75t_L g930 ( .A1(n_84), .A2(n_122), .B1(n_314), .B2(n_448), .Y(n_930) );
OAI22xp33_ASAP7_75t_L g946 ( .A1(n_84), .A2(n_122), .B1(n_947), .B2(n_949), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g1166 ( .A1(n_85), .A2(n_150), .B1(n_719), .B2(n_1167), .Y(n_1166) );
AOI22xp33_ASAP7_75t_SL g1174 ( .A1(n_85), .A2(n_294), .B1(n_1175), .B2(n_1179), .Y(n_1174) );
AOI221xp5_ASAP7_75t_L g717 ( .A1(n_86), .A2(n_292), .B1(n_718), .B2(n_719), .C(n_721), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_86), .A2(n_148), .B1(n_771), .B2(n_772), .Y(n_770) );
INVx1_ASAP7_75t_L g538 ( .A(n_87), .Y(n_538) );
INVx1_ASAP7_75t_L g1097 ( .A(n_88), .Y(n_1097) );
AOI22xp33_ASAP7_75t_SL g609 ( .A1(n_89), .A2(n_241), .B1(n_604), .B2(n_610), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_89), .A2(n_91), .B1(n_511), .B2(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g692 ( .A(n_90), .Y(n_692) );
OAI211xp5_ASAP7_75t_SL g701 ( .A1(n_90), .A2(n_662), .B(n_702), .C(n_703), .Y(n_701) );
AOI22xp33_ASAP7_75t_SL g592 ( .A1(n_91), .A2(n_186), .B1(n_593), .B2(n_596), .Y(n_592) );
INVx1_ASAP7_75t_L g933 ( .A(n_92), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g1286 ( .A1(n_93), .A2(n_115), .B1(n_1287), .B2(n_1291), .Y(n_1286) );
XOR2x2_ASAP7_75t_L g532 ( .A(n_94), .B(n_533), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g1339 ( .A1(n_95), .A2(n_134), .B1(n_1294), .B2(n_1297), .Y(n_1339) );
OAI22xp33_ASAP7_75t_L g995 ( .A1(n_96), .A2(n_103), .B1(n_314), .B2(n_448), .Y(n_995) );
OAI22xp33_ASAP7_75t_L g1003 ( .A1(n_96), .A2(n_103), .B1(n_872), .B2(n_947), .Y(n_1003) );
INVx1_ASAP7_75t_L g791 ( .A(n_97), .Y(n_791) );
OAI211xp5_ASAP7_75t_L g833 ( .A1(n_98), .A2(n_834), .B(n_837), .C(n_843), .Y(n_833) );
INVx1_ASAP7_75t_L g860 ( .A(n_98), .Y(n_860) );
INVx1_ASAP7_75t_L g329 ( .A(n_99), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_100), .A2(n_187), .B1(n_522), .B2(n_542), .Y(n_541) );
OAI22xp33_ASAP7_75t_L g557 ( .A1(n_100), .A2(n_187), .B1(n_479), .B2(n_480), .Y(n_557) );
OAI221xp5_ASAP7_75t_L g1263 ( .A1(n_101), .A2(n_290), .B1(n_459), .B2(n_479), .C(n_1264), .Y(n_1263) );
INVx1_ASAP7_75t_L g1276 ( .A(n_101), .Y(n_1276) );
INVx1_ASAP7_75t_L g902 ( .A(n_102), .Y(n_902) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_105), .Y(n_307) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_105), .B(n_305), .Y(n_1288) );
CKINVDCx5p33_ASAP7_75t_R g991 ( .A(n_107), .Y(n_991) );
INVx1_ASAP7_75t_L g1049 ( .A(n_108), .Y(n_1049) );
INVx1_ASAP7_75t_L g1247 ( .A(n_109), .Y(n_1247) );
INVx1_ASAP7_75t_L g1050 ( .A(n_110), .Y(n_1050) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_112), .B(n_1290), .Y(n_1289) );
INVx1_ASAP7_75t_L g1296 ( .A(n_112), .Y(n_1296) );
AOI22xp5_ASAP7_75t_L g1318 ( .A1(n_113), .A2(n_184), .B1(n_1294), .B2(n_1297), .Y(n_1318) );
INVx1_ASAP7_75t_L g1089 ( .A(n_114), .Y(n_1089) );
OAI22xp33_ASAP7_75t_SL g935 ( .A1(n_117), .A2(n_272), .B1(n_887), .B2(n_936), .Y(n_935) );
OAI22xp5_ASAP7_75t_L g938 ( .A1(n_117), .A2(n_272), .B1(n_862), .B2(n_939), .Y(n_938) );
INVx1_ASAP7_75t_L g1249 ( .A(n_119), .Y(n_1249) );
INVx1_ASAP7_75t_L g1086 ( .A(n_120), .Y(n_1086) );
AOI22xp33_ASAP7_75t_L g1119 ( .A1(n_120), .A2(n_237), .B1(n_1120), .B2(n_1121), .Y(n_1119) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_121), .Y(n_499) );
INVx1_ASAP7_75t_L g960 ( .A(n_123), .Y(n_960) );
INVx1_ASAP7_75t_L g1208 ( .A(n_124), .Y(n_1208) );
OAI22xp33_ASAP7_75t_L g1072 ( .A1(n_125), .A2(n_240), .B1(n_314), .B2(n_448), .Y(n_1072) );
OAI22xp33_ASAP7_75t_L g1074 ( .A1(n_125), .A2(n_240), .B1(n_872), .B2(n_1075), .Y(n_1074) );
OAI22xp5_ASAP7_75t_L g1149 ( .A1(n_126), .A2(n_256), .B1(n_1150), .B2(n_1151), .Y(n_1149) );
OAI22xp5_ASAP7_75t_L g1187 ( .A1(n_126), .A2(n_256), .B1(n_696), .B2(n_846), .Y(n_1187) );
INVx2_ASAP7_75t_L g339 ( .A(n_127), .Y(n_339) );
INVx1_ASAP7_75t_L g387 ( .A(n_127), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_128), .Y(n_348) );
INVx1_ASAP7_75t_L g1515 ( .A(n_129), .Y(n_1515) );
INVx1_ASAP7_75t_L g562 ( .A(n_130), .Y(n_562) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_131), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_133), .A2(n_268), .B1(n_479), .B2(n_480), .Y(n_700) );
CKINVDCx5p33_ASAP7_75t_R g1007 ( .A(n_135), .Y(n_1007) );
INVx1_ASAP7_75t_L g1146 ( .A(n_136), .Y(n_1146) );
OAI22xp5_ASAP7_75t_SL g1500 ( .A1(n_137), .A2(n_230), .B1(n_458), .B2(n_479), .Y(n_1500) );
INVx1_ASAP7_75t_L g1055 ( .A(n_138), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g1293 ( .A1(n_139), .A2(n_273), .B1(n_1294), .B2(n_1297), .Y(n_1293) );
INVx1_ASAP7_75t_L g911 ( .A(n_140), .Y(n_911) );
INVx1_ASAP7_75t_L g1518 ( .A(n_141), .Y(n_1518) );
INVx1_ASAP7_75t_L g1220 ( .A(n_143), .Y(n_1220) );
AOI22xp5_ASAP7_75t_L g1338 ( .A1(n_144), .A2(n_147), .B1(n_1287), .B2(n_1291), .Y(n_1338) );
INVx1_ASAP7_75t_L g575 ( .A(n_145), .Y(n_575) );
CKINVDCx5p33_ASAP7_75t_R g1016 ( .A(n_146), .Y(n_1016) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_148), .A2(n_246), .B1(n_718), .B2(n_719), .C(n_723), .Y(n_722) );
INVxp67_ASAP7_75t_SL g1110 ( .A(n_149), .Y(n_1110) );
OAI22xp5_ASAP7_75t_L g1130 ( .A1(n_149), .A2(n_204), .B1(n_702), .B2(n_1131), .Y(n_1130) );
INVx1_ASAP7_75t_L g1104 ( .A(n_152), .Y(n_1104) );
XOR2xp5_ASAP7_75t_L g1142 ( .A(n_153), .B(n_1143), .Y(n_1142) );
AOI22xp33_ASAP7_75t_L g1322 ( .A1(n_153), .A2(n_155), .B1(n_1294), .B2(n_1297), .Y(n_1322) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_154), .Y(n_517) );
INVx1_ASAP7_75t_L g1516 ( .A(n_157), .Y(n_1516) );
AOI31xp33_ASAP7_75t_L g712 ( .A1(n_158), .A2(n_713), .A3(n_731), .B(n_742), .Y(n_712) );
NAND2xp33_ASAP7_75t_SL g759 ( .A(n_158), .B(n_760), .Y(n_759) );
INVxp67_ASAP7_75t_SL g775 ( .A(n_158), .Y(n_775) );
INVx1_ASAP7_75t_L g1206 ( .A(n_159), .Y(n_1206) );
BUFx3_ASAP7_75t_L g345 ( .A(n_160), .Y(n_345) );
INVx1_ASAP7_75t_L g1510 ( .A(n_161), .Y(n_1510) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_162), .Y(n_380) );
INVx1_ASAP7_75t_L g895 ( .A(n_163), .Y(n_895) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_164), .Y(n_504) );
CKINVDCx5p33_ASAP7_75t_R g1017 ( .A(n_165), .Y(n_1017) );
AOI22xp5_ASAP7_75t_L g1302 ( .A1(n_166), .A2(n_167), .B1(n_1294), .B2(n_1297), .Y(n_1302) );
INVx1_ASAP7_75t_L g793 ( .A(n_168), .Y(n_793) );
AOI22xp5_ASAP7_75t_L g1309 ( .A1(n_169), .A2(n_255), .B1(n_1287), .B2(n_1291), .Y(n_1309) );
OAI22xp33_ASAP7_75t_L g528 ( .A1(n_170), .A2(n_291), .B1(n_479), .B2(n_480), .Y(n_528) );
CKINVDCx5p33_ASAP7_75t_R g501 ( .A(n_171), .Y(n_501) );
CKINVDCx5p33_ASAP7_75t_R g1019 ( .A(n_172), .Y(n_1019) );
XOR2xp5_ASAP7_75t_L g1039 ( .A(n_173), .B(n_1040), .Y(n_1039) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_174), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_175), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g1156 ( .A1(n_176), .A2(n_234), .B1(n_736), .B2(n_1157), .Y(n_1156) );
AOI22xp33_ASAP7_75t_L g1171 ( .A1(n_176), .A2(n_220), .B1(n_1172), .B2(n_1173), .Y(n_1171) );
OAI211xp5_ASAP7_75t_L g931 ( .A1(n_177), .A2(n_880), .B(n_883), .C(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g945 ( .A(n_177), .Y(n_945) );
INVx1_ASAP7_75t_L g1267 ( .A(n_178), .Y(n_1267) );
INVx1_ASAP7_75t_L g934 ( .A(n_180), .Y(n_934) );
OAI211xp5_ASAP7_75t_L g941 ( .A1(n_180), .A2(n_466), .B(n_942), .C(n_944), .Y(n_941) );
OAI211xp5_ASAP7_75t_L g988 ( .A1(n_181), .A2(n_882), .B(n_989), .C(n_990), .Y(n_988) );
INVx1_ASAP7_75t_L g1002 ( .A(n_181), .Y(n_1002) );
INVx1_ASAP7_75t_L g1204 ( .A(n_182), .Y(n_1204) );
INVx1_ASAP7_75t_L g900 ( .A(n_183), .Y(n_900) );
XOR2x2_ASAP7_75t_L g1490 ( .A(n_184), .B(n_1491), .Y(n_1490) );
AOI22xp33_ASAP7_75t_L g1531 ( .A1(n_184), .A2(n_1532), .B1(n_1535), .B2(n_1538), .Y(n_1531) );
INVx1_ASAP7_75t_L g1197 ( .A(n_185), .Y(n_1197) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_186), .A2(n_241), .B1(n_614), .B2(n_615), .Y(n_613) );
INVx1_ASAP7_75t_L g728 ( .A(n_189), .Y(n_728) );
AOI22xp33_ASAP7_75t_SL g762 ( .A1(n_189), .A2(n_271), .B1(n_604), .B2(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g806 ( .A(n_190), .Y(n_806) );
INVx1_ASAP7_75t_L g875 ( .A(n_191), .Y(n_875) );
INVx1_ASAP7_75t_L g957 ( .A(n_192), .Y(n_957) );
INVx1_ASAP7_75t_L g1096 ( .A(n_194), .Y(n_1096) );
CKINVDCx5p33_ASAP7_75t_R g674 ( .A(n_195), .Y(n_674) );
INVx1_ASAP7_75t_L g993 ( .A(n_196), .Y(n_993) );
OAI211xp5_ASAP7_75t_L g998 ( .A1(n_196), .A2(n_466), .B(n_999), .C(n_1001), .Y(n_998) );
INVxp67_ASAP7_75t_SL g746 ( .A(n_197), .Y(n_746) );
AOI22xp33_ASAP7_75t_SL g620 ( .A1(n_198), .A2(n_284), .B1(n_621), .B2(n_626), .Y(n_620) );
OAI211xp5_ASAP7_75t_L g1067 ( .A1(n_199), .A2(n_882), .B(n_883), .C(n_1068), .Y(n_1067) );
INVx1_ASAP7_75t_L g1079 ( .A(n_199), .Y(n_1079) );
INVx1_ASAP7_75t_L g1070 ( .A(n_200), .Y(n_1070) );
OAI211xp5_ASAP7_75t_L g1077 ( .A1(n_200), .A2(n_466), .B(n_943), .C(n_1078), .Y(n_1077) );
INVx1_ASAP7_75t_L g1255 ( .A(n_201), .Y(n_1255) );
INVx1_ASAP7_75t_L g725 ( .A(n_202), .Y(n_725) );
INVx1_ASAP7_75t_L g645 ( .A(n_203), .Y(n_645) );
INVx1_ASAP7_75t_L g1519 ( .A(n_205), .Y(n_1519) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_206), .B(n_473), .Y(n_1266) );
INVxp67_ASAP7_75t_SL g1273 ( .A(n_206), .Y(n_1273) );
OAI211xp5_ASAP7_75t_SL g873 ( .A1(n_207), .A2(n_662), .B(n_855), .C(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g885 ( .A(n_207), .Y(n_885) );
INVx1_ASAP7_75t_L g1221 ( .A(n_208), .Y(n_1221) );
CKINVDCx5p33_ASAP7_75t_R g682 ( .A(n_209), .Y(n_682) );
INVx1_ASAP7_75t_L g1045 ( .A(n_210), .Y(n_1045) );
CKINVDCx5p33_ASAP7_75t_R g496 ( .A(n_211), .Y(n_496) );
CKINVDCx5p33_ASAP7_75t_R g1009 ( .A(n_212), .Y(n_1009) );
OAI211xp5_ASAP7_75t_L g689 ( .A1(n_213), .A2(n_422), .B(n_690), .C(n_691), .Y(n_689) );
INVx1_ASAP7_75t_L g708 ( .A(n_213), .Y(n_708) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_214), .Y(n_357) );
INVx1_ASAP7_75t_L g1069 ( .A(n_215), .Y(n_1069) );
OAI22xp33_ASAP7_75t_L g877 ( .A1(n_216), .A2(n_282), .B1(n_862), .B2(n_863), .Y(n_877) );
OAI22xp5_ASAP7_75t_L g886 ( .A1(n_216), .A2(n_282), .B1(n_887), .B2(n_888), .Y(n_886) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_217), .Y(n_318) );
INVx1_ASAP7_75t_L g962 ( .A(n_218), .Y(n_962) );
INVx1_ASAP7_75t_L g646 ( .A(n_219), .Y(n_646) );
INVx1_ASAP7_75t_L g968 ( .A(n_221), .Y(n_968) );
INVx1_ASAP7_75t_L g1198 ( .A(n_223), .Y(n_1198) );
INVx1_ASAP7_75t_L g519 ( .A(n_225), .Y(n_519) );
OAI211xp5_ASAP7_75t_L g525 ( .A1(n_225), .A2(n_463), .B(n_466), .C(n_526), .Y(n_525) );
CKINVDCx5p33_ASAP7_75t_R g672 ( .A(n_226), .Y(n_672) );
INVx1_ASAP7_75t_L g1054 ( .A(n_227), .Y(n_1054) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_228), .Y(n_342) );
INVx1_ASAP7_75t_L g1496 ( .A(n_229), .Y(n_1496) );
CKINVDCx5p33_ASAP7_75t_R g1012 ( .A(n_231), .Y(n_1012) );
CKINVDCx5p33_ASAP7_75t_R g1014 ( .A(n_232), .Y(n_1014) );
INVx1_ASAP7_75t_L g1114 ( .A(n_233), .Y(n_1114) );
XOR2xp5_ASAP7_75t_L g1536 ( .A(n_235), .B(n_1537), .Y(n_1536) );
INVx1_ASAP7_75t_L g1099 ( .A(n_237), .Y(n_1099) );
INVx1_ASAP7_75t_L g1251 ( .A(n_238), .Y(n_1251) );
INVx1_ASAP7_75t_L g570 ( .A(n_239), .Y(n_570) );
INVx1_ASAP7_75t_L g1194 ( .A(n_242), .Y(n_1194) );
INVx1_ASAP7_75t_L g842 ( .A(n_243), .Y(n_842) );
OAI211xp5_ASAP7_75t_L g854 ( .A1(n_243), .A2(n_662), .B(n_855), .C(n_857), .Y(n_854) );
INVx1_ASAP7_75t_L g1513 ( .A(n_244), .Y(n_1513) );
INVx1_ASAP7_75t_L g1202 ( .A(n_245), .Y(n_1202) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_246), .A2(n_292), .B1(n_766), .B2(n_768), .Y(n_765) );
INVx1_ASAP7_75t_L g640 ( .A(n_247), .Y(n_640) );
INVxp67_ASAP7_75t_SL g1275 ( .A(n_248), .Y(n_1275) );
CKINVDCx5p33_ASAP7_75t_R g431 ( .A(n_249), .Y(n_431) );
INVx1_ASAP7_75t_L g567 ( .A(n_251), .Y(n_567) );
BUFx3_ASAP7_75t_L g322 ( .A(n_253), .Y(n_322) );
INVx1_ASAP7_75t_L g447 ( .A(n_253), .Y(n_447) );
INVx1_ASAP7_75t_L g839 ( .A(n_254), .Y(n_839) );
XOR2x2_ASAP7_75t_L g868 ( .A(n_257), .B(n_869), .Y(n_868) );
CKINVDCx5p33_ASAP7_75t_R g694 ( .A(n_258), .Y(n_694) );
INVx1_ASAP7_75t_L g1243 ( .A(n_260), .Y(n_1243) );
INVx1_ASAP7_75t_L g1115 ( .A(n_261), .Y(n_1115) );
OAI211xp5_ASAP7_75t_L g515 ( .A1(n_262), .A2(n_421), .B(n_422), .C(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g527 ( .A(n_262), .Y(n_527) );
INVx1_ASAP7_75t_L g561 ( .A(n_263), .Y(n_561) );
INVx1_ASAP7_75t_L g907 ( .A(n_264), .Y(n_907) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_265), .Y(n_373) );
INVx1_ASAP7_75t_L g1223 ( .A(n_267), .Y(n_1223) );
OAI211xp5_ASAP7_75t_L g535 ( .A1(n_269), .A2(n_422), .B(n_536), .C(n_537), .Y(n_535) );
INVx1_ASAP7_75t_L g553 ( .A(n_269), .Y(n_553) );
INVx1_ASAP7_75t_L g337 ( .A(n_270), .Y(n_337) );
INVx2_ASAP7_75t_L g385 ( .A(n_270), .Y(n_385) );
INVx1_ASAP7_75t_L g635 ( .A(n_270), .Y(n_635) );
XOR2x2_ASAP7_75t_L g985 ( .A(n_273), .B(n_986), .Y(n_985) );
INVx1_ASAP7_75t_L g1105 ( .A(n_274), .Y(n_1105) );
CKINVDCx5p33_ASAP7_75t_R g678 ( .A(n_275), .Y(n_678) );
INVx1_ASAP7_75t_L g1254 ( .A(n_276), .Y(n_1254) );
INVx1_ASAP7_75t_L g814 ( .A(n_277), .Y(n_814) );
INVx1_ASAP7_75t_L g975 ( .A(n_278), .Y(n_975) );
INVx1_ASAP7_75t_L g974 ( .A(n_279), .Y(n_974) );
INVx1_ASAP7_75t_L g1059 ( .A(n_280), .Y(n_1059) );
INVx1_ASAP7_75t_L g970 ( .A(n_281), .Y(n_970) );
INVx1_ASAP7_75t_L g910 ( .A(n_283), .Y(n_910) );
XNOR2xp5_ASAP7_75t_L g486 ( .A(n_285), .B(n_487), .Y(n_486) );
OAI22xp33_ASAP7_75t_L g520 ( .A1(n_286), .A2(n_291), .B1(n_439), .B2(n_441), .Y(n_520) );
INVx1_ASAP7_75t_L g876 ( .A(n_287), .Y(n_876) );
OAI211xp5_ASAP7_75t_L g879 ( .A1(n_287), .A2(n_880), .B(n_883), .C(n_884), .Y(n_879) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_288), .Y(n_382) );
INVx1_ASAP7_75t_L g1147 ( .A(n_289), .Y(n_1147) );
INVx1_ASAP7_75t_L g744 ( .A(n_293), .Y(n_744) );
INVx1_ASAP7_75t_L g804 ( .A(n_295), .Y(n_804) );
INVx1_ASAP7_75t_L g437 ( .A(n_296), .Y(n_437) );
OAI211xp5_ASAP7_75t_L g462 ( .A1(n_296), .A2(n_463), .B(n_466), .C(n_470), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_323), .B(n_1280), .Y(n_297) );
INVx2_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_308), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g1530 ( .A(n_302), .B(n_311), .Y(n_1530) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g1534 ( .A(n_304), .B(n_307), .Y(n_1534) );
INVx1_ASAP7_75t_L g1539 ( .A(n_304), .Y(n_1539) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g1542 ( .A(n_307), .B(n_1539), .Y(n_1542) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_313), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x4_ASAP7_75t_L g453 ( .A(n_311), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x4_ASAP7_75t_L g418 ( .A(n_312), .B(n_322), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_313), .A2(n_449), .B1(n_1104), .B2(n_1105), .Y(n_1103) );
AOI22xp33_ASAP7_75t_L g1185 ( .A1(n_313), .A2(n_449), .B1(n_1146), .B2(n_1147), .Y(n_1185) );
AND2x4_ASAP7_75t_SL g1529 ( .A(n_313), .B(n_1530), .Y(n_1529) );
INVx3_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OR2x6_ASAP7_75t_L g314 ( .A(n_315), .B(n_320), .Y(n_314) );
OR2x6_ASAP7_75t_L g445 ( .A(n_315), .B(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g522 ( .A(n_315), .B(n_446), .Y(n_522) );
INVx1_ASAP7_75t_L g587 ( .A(n_315), .Y(n_587) );
BUFx4f_ASAP7_75t_L g956 ( .A(n_315), .Y(n_956) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx4f_ASAP7_75t_L g395 ( .A(n_316), .Y(n_395) );
INVx3_ASAP7_75t_L g440 ( .A(n_316), .Y(n_440) );
INVx3_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx2_ASAP7_75t_L g401 ( .A(n_318), .Y(n_401) );
INVx2_ASAP7_75t_L g406 ( .A(n_318), .Y(n_406) );
NAND2x1_ASAP7_75t_L g410 ( .A(n_318), .B(n_319), .Y(n_410) );
AND2x2_ASAP7_75t_L g427 ( .A(n_318), .B(n_319), .Y(n_427) );
INVx1_ASAP7_75t_L g436 ( .A(n_318), .Y(n_436) );
AND2x2_ASAP7_75t_L g450 ( .A(n_318), .B(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_319), .B(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g405 ( .A(n_319), .B(n_406), .Y(n_405) );
BUFx2_ASAP7_75t_L g430 ( .A(n_319), .Y(n_430) );
INVx2_ASAP7_75t_L g451 ( .A(n_319), .Y(n_451) );
INVx1_ASAP7_75t_L g603 ( .A(n_319), .Y(n_603) );
AND2x2_ASAP7_75t_L g605 ( .A(n_319), .B(n_401), .Y(n_605) );
OR2x6_ASAP7_75t_L g439 ( .A(n_320), .B(n_440), .Y(n_439) );
INVxp67_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g424 ( .A(n_321), .Y(n_424) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x4_ASAP7_75t_L g434 ( .A(n_322), .B(n_435), .Y(n_434) );
BUFx2_ASAP7_75t_L g443 ( .A(n_322), .Y(n_443) );
XNOR2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_780), .Y(n_323) );
OAI22xp33_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_326), .B1(n_529), .B2(n_779), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
XNOR2x1_ASAP7_75t_L g327 ( .A(n_328), .B(n_486), .Y(n_327) );
XNOR2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
AND3x1_ASAP7_75t_L g330 ( .A(n_331), .B(n_419), .C(n_456), .Y(n_330) );
NOR2xp33_ASAP7_75t_SL g331 ( .A(n_332), .B(n_389), .Y(n_331) );
OAI33xp33_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_341), .A3(n_356), .B1(n_368), .B2(n_377), .B3(n_383), .Y(n_332) );
OAI33xp33_ASAP7_75t_L g505 ( .A1(n_333), .A2(n_383), .A3(n_506), .B1(n_508), .B2(n_509), .B3(n_513), .Y(n_505) );
OAI33xp33_ASAP7_75t_L g559 ( .A1(n_333), .A2(n_383), .A3(n_560), .B1(n_563), .B2(n_568), .B3(n_574), .Y(n_559) );
OAI33xp33_ASAP7_75t_L g669 ( .A1(n_333), .A2(n_383), .A3(n_670), .B1(n_673), .B2(n_676), .B3(n_680), .Y(n_669) );
BUFx3_ASAP7_75t_L g1084 ( .A(n_333), .Y(n_1084) );
OAI33xp33_ASAP7_75t_L g1520 ( .A1(n_333), .A2(n_383), .A3(n_1521), .B1(n_1522), .B2(n_1523), .B3(n_1525), .Y(n_1520) );
BUFx4f_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx4f_ASAP7_75t_L g816 ( .A(n_334), .Y(n_816) );
BUFx2_ASAP7_75t_L g893 ( .A(n_334), .Y(n_893) );
BUFx8_ASAP7_75t_L g1022 ( .A(n_334), .Y(n_1022) );
OR2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_338), .Y(n_334) );
AND2x2_ASAP7_75t_SL g417 ( .A(n_335), .B(n_418), .Y(n_417) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_335), .Y(n_485) );
INVx1_ASAP7_75t_L g810 ( .A(n_335), .Y(n_810) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx2_ASAP7_75t_L g455 ( .A(n_336), .Y(n_455) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp33_ASAP7_75t_SL g338 ( .A(n_339), .B(n_340), .Y(n_338) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_339), .Y(n_483) );
AND3x4_ASAP7_75t_L g618 ( .A(n_339), .B(n_473), .C(n_619), .Y(n_618) );
INVx3_ASAP7_75t_L g388 ( .A(n_340), .Y(n_388) );
BUFx3_ASAP7_75t_L g473 ( .A(n_340), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_343), .B1(n_348), .B2(n_349), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_342), .A2(n_380), .B1(n_394), .B2(n_396), .Y(n_393) );
OAI22xp33_ASAP7_75t_L g560 ( .A1(n_343), .A2(n_507), .B1(n_561), .B2(n_562), .Y(n_560) );
OAI22xp33_ASAP7_75t_L g574 ( .A1(n_343), .A2(n_381), .B1(n_575), .B2(n_576), .Y(n_574) );
OAI22xp33_ASAP7_75t_L g670 ( .A1(n_343), .A2(n_507), .B1(n_671), .B2(n_672), .Y(n_670) );
OAI22xp33_ASAP7_75t_L g680 ( .A1(n_343), .A2(n_381), .B1(n_681), .B2(n_682), .Y(n_680) );
OAI22xp33_ASAP7_75t_L g1210 ( .A1(n_343), .A2(n_349), .B1(n_1197), .B2(n_1206), .Y(n_1210) );
OAI22xp33_ASAP7_75t_L g1215 ( .A1(n_343), .A2(n_381), .B1(n_1198), .B2(n_1208), .Y(n_1215) );
OAI22xp33_ASAP7_75t_L g1242 ( .A1(n_343), .A2(n_1243), .B1(n_1244), .B2(n_1245), .Y(n_1242) );
OAI22xp33_ASAP7_75t_L g1253 ( .A1(n_343), .A2(n_507), .B1(n_1254), .B2(n_1255), .Y(n_1253) );
OAI22xp33_ASAP7_75t_L g1525 ( .A1(n_343), .A2(n_1510), .B1(n_1516), .B2(n_1526), .Y(n_1525) );
BUFx4f_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g379 ( .A(n_344), .Y(n_379) );
OR2x4_ASAP7_75t_L g458 ( .A(n_344), .B(n_388), .Y(n_458) );
OR2x4_ASAP7_75t_L g479 ( .A(n_344), .B(n_461), .Y(n_479) );
BUFx3_ASAP7_75t_L g820 ( .A(n_344), .Y(n_820) );
BUFx3_ASAP7_75t_L g896 ( .A(n_344), .Y(n_896) );
OR2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_345), .Y(n_355) );
INVx2_ASAP7_75t_L g362 ( .A(n_345), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_345), .B(n_354), .Y(n_367) );
AND2x4_ASAP7_75t_L g468 ( .A(n_345), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g625 ( .A(n_346), .Y(n_625) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVxp67_ASAP7_75t_L g361 ( .A(n_347), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_348), .A2(n_382), .B1(n_412), .B2(n_413), .Y(n_411) );
INVx3_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g898 ( .A(n_350), .Y(n_898) );
INVx2_ASAP7_75t_L g1026 ( .A(n_350), .Y(n_1026) );
INVx3_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_351), .Y(n_507) );
INVx4_ASAP7_75t_L g856 ( .A(n_351), .Y(n_856) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx3_ASAP7_75t_L g381 ( .A(n_352), .Y(n_381) );
BUFx2_ASAP7_75t_L g465 ( .A(n_352), .Y(n_465) );
NAND2x1p5_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
BUFx2_ASAP7_75t_L g476 ( .A(n_353), .Y(n_476) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g469 ( .A(n_354), .Y(n_469) );
BUFx2_ASAP7_75t_L g474 ( .A(n_355), .Y(n_474) );
AND2x4_ASAP7_75t_L g616 ( .A(n_355), .B(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g707 ( .A(n_355), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_358), .B1(n_363), .B2(n_364), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_357), .A2(n_369), .B1(n_403), .B2(n_407), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_358), .A2(n_364), .B1(n_496), .B2(n_503), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g1523 ( .A1(n_358), .A2(n_1513), .B1(n_1519), .B2(n_1524), .Y(n_1523) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g460 ( .A(n_359), .B(n_461), .Y(n_460) );
AND2x4_ASAP7_75t_L g549 ( .A(n_359), .B(n_461), .Y(n_549) );
BUFx6f_ASAP7_75t_L g718 ( .A(n_359), .Y(n_718) );
INVx2_ASAP7_75t_L g1030 ( .A(n_359), .Y(n_1030) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g372 ( .A(n_360), .Y(n_372) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_360), .Y(n_511) );
BUFx8_ASAP7_75t_L g566 ( .A(n_360), .Y(n_566) );
AND2x4_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
AND2x4_ASAP7_75t_L g624 ( .A(n_362), .B(n_625), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_363), .A2(n_373), .B1(n_394), .B2(n_415), .Y(n_414) );
OAI22xp5_ASAP7_75t_L g1522 ( .A1(n_364), .A2(n_677), .B1(n_1512), .B2(n_1518), .Y(n_1522) );
INVx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx3_ASAP7_75t_L g512 ( .A(n_365), .Y(n_512) );
CKINVDCx8_ASAP7_75t_R g825 ( .A(n_365), .Y(n_825) );
INVx3_ASAP7_75t_L g1524 ( .A(n_365), .Y(n_1524) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g572 ( .A(n_366), .Y(n_572) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx2_ASAP7_75t_L g376 ( .A(n_367), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_370), .B1(n_373), .B2(n_374), .Y(n_368) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx3_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx2_ASAP7_75t_L g1161 ( .A(n_372), .Y(n_1161) );
INVx1_ASAP7_75t_L g1167 ( .A(n_372), .Y(n_1167) );
BUFx2_ASAP7_75t_L g1248 ( .A(n_372), .Y(n_1248) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_374), .A2(n_564), .B1(n_565), .B2(n_567), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_374), .A2(n_569), .B1(n_674), .B2(n_675), .Y(n_673) );
OAI22xp33_ASAP7_75t_SL g1211 ( .A1(n_374), .A2(n_824), .B1(n_1194), .B2(n_1202), .Y(n_1211) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx2_ASAP7_75t_L g982 ( .A(n_375), .Y(n_982) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OR2x6_ASAP7_75t_L g480 ( .A(n_376), .B(n_388), .Y(n_480) );
BUFx3_ASAP7_75t_L g827 ( .A(n_376), .Y(n_827) );
OAI22xp33_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_380), .B1(n_381), .B2(n_382), .Y(n_377) );
OAI22xp33_ASAP7_75t_L g506 ( .A1(n_378), .A2(n_492), .B1(n_499), .B2(n_507), .Y(n_506) );
OAI22xp33_ASAP7_75t_L g513 ( .A1(n_378), .A2(n_381), .B1(n_494), .B2(n_501), .Y(n_513) );
INVx2_ASAP7_75t_SL g1088 ( .A(n_378), .Y(n_1088) );
OAI22xp33_ASAP7_75t_L g1098 ( .A1(n_378), .A2(n_1099), .B1(n_1100), .B2(n_1101), .Y(n_1098) );
OAI22xp33_ASAP7_75t_L g1521 ( .A1(n_378), .A2(n_381), .B1(n_1509), .B2(n_1515), .Y(n_1521) );
INVx2_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
INVx3_ASAP7_75t_L g979 ( .A(n_379), .Y(n_979) );
INVx2_ASAP7_75t_L g822 ( .A(n_381), .Y(n_822) );
BUFx6f_ASAP7_75t_L g1100 ( .A(n_381), .Y(n_1100) );
OR2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_386), .Y(n_383) );
AND2x4_ASAP7_75t_L g391 ( .A(n_384), .B(n_392), .Y(n_391) );
OR2x6_ASAP7_75t_L g730 ( .A(n_384), .B(n_386), .Y(n_730) );
BUFx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g619 ( .A(n_385), .Y(n_619) );
NAND2x1p5_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
NAND3x1_ASAP7_75t_L g633 ( .A(n_387), .B(n_388), .C(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g461 ( .A(n_388), .Y(n_461) );
AND2x4_ASAP7_75t_L g467 ( .A(n_388), .B(n_468), .Y(n_467) );
OAI33xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_393), .A3(n_402), .B1(n_411), .B2(n_414), .B3(n_416), .Y(n_389) );
OAI33xp33_ASAP7_75t_L g577 ( .A1(n_390), .A2(n_578), .A3(n_580), .B1(n_583), .B2(n_584), .B3(n_585), .Y(n_577) );
OAI33xp33_ASAP7_75t_L g683 ( .A1(n_390), .A2(n_584), .A3(n_684), .B1(n_685), .B2(n_686), .B3(n_687), .Y(n_683) );
OAI22xp5_ASAP7_75t_SL g1117 ( .A1(n_390), .A2(n_921), .B1(n_1118), .B2(n_1123), .Y(n_1117) );
OAI33xp33_ASAP7_75t_L g1256 ( .A1(n_390), .A2(n_584), .A3(n_1257), .B1(n_1258), .B2(n_1259), .B3(n_1260), .Y(n_1256) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g490 ( .A(n_391), .Y(n_490) );
INVx4_ASAP7_75t_L g607 ( .A(n_391), .Y(n_607) );
INVx2_ASAP7_75t_L g789 ( .A(n_391), .Y(n_789) );
INVx1_ASAP7_75t_L g1010 ( .A(n_391), .Y(n_1010) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_394), .A2(n_492), .B1(n_493), .B2(n_494), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_394), .A2(n_396), .B1(n_503), .B2(n_504), .Y(n_502) );
OAI22xp33_ASAP7_75t_L g578 ( .A1(n_394), .A2(n_561), .B1(n_575), .B2(n_579), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_394), .A2(n_415), .B1(n_671), .B2(n_681), .Y(n_684) );
OAI22xp33_ASAP7_75t_L g1196 ( .A1(n_394), .A2(n_1197), .B1(n_1198), .B2(n_1199), .Y(n_1196) );
OAI22xp5_ASAP7_75t_L g1508 ( .A1(n_394), .A2(n_396), .B1(n_1509), .B2(n_1510), .Y(n_1508) );
OAI22xp5_ASAP7_75t_L g1517 ( .A1(n_394), .A2(n_493), .B1(n_1518), .B2(n_1519), .Y(n_1517) );
INVx4_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx3_ASAP7_75t_L g792 ( .A(n_395), .Y(n_792) );
BUFx6f_ASAP7_75t_L g973 ( .A(n_395), .Y(n_973) );
OAI22xp5_ASAP7_75t_L g1201 ( .A1(n_396), .A2(n_1202), .B1(n_1203), .B2(n_1204), .Y(n_1201) );
OAI22xp5_ASAP7_75t_L g1260 ( .A1(n_396), .A2(n_1249), .B1(n_1252), .B2(n_1261), .Y(n_1260) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx4_ASAP7_75t_L g415 ( .A(n_398), .Y(n_415) );
INVx2_ASAP7_75t_SL g493 ( .A(n_398), .Y(n_493) );
INVx1_ASAP7_75t_L g579 ( .A(n_398), .Y(n_579) );
BUFx6f_ASAP7_75t_L g795 ( .A(n_398), .Y(n_795) );
INVx1_ASAP7_75t_L g1199 ( .A(n_398), .Y(n_1199) );
INVx8_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
OR2x2_ASAP7_75t_L g442 ( .A(n_399), .B(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g542 ( .A(n_399), .B(n_424), .Y(n_542) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_403), .A2(n_413), .B1(n_496), .B2(n_497), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_403), .A2(n_499), .B1(n_500), .B2(n_501), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g1511 ( .A1(n_403), .A2(n_500), .B1(n_1512), .B2(n_1513), .Y(n_1511) );
OAI22xp5_ASAP7_75t_L g1514 ( .A1(n_403), .A2(n_1207), .B1(n_1515), .B2(n_1516), .Y(n_1514) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g798 ( .A(n_404), .Y(n_798) );
BUFx2_ASAP7_75t_L g918 ( .A(n_404), .Y(n_918) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx2_ASAP7_75t_L g412 ( .A(n_405), .Y(n_412) );
INVx1_ASAP7_75t_L g582 ( .A(n_405), .Y(n_582) );
BUFx2_ASAP7_75t_L g803 ( .A(n_405), .Y(n_803) );
BUFx3_ASAP7_75t_L g967 ( .A(n_405), .Y(n_967) );
AND2x2_ASAP7_75t_L g602 ( .A(n_406), .B(n_603), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_407), .A2(n_564), .B1(n_570), .B2(n_581), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_407), .A2(n_581), .B1(n_674), .B2(n_678), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_407), .A2(n_581), .B1(n_672), .B2(n_682), .Y(n_686) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g421 ( .A(n_408), .Y(n_421) );
INVx2_ASAP7_75t_L g919 ( .A(n_408), .Y(n_919) );
INVx4_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_409), .Y(n_500) );
BUFx4f_ASAP7_75t_L g690 ( .A(n_409), .Y(n_690) );
BUFx4f_ASAP7_75t_L g836 ( .A(n_409), .Y(n_836) );
BUFx4f_ASAP7_75t_L g969 ( .A(n_409), .Y(n_969) );
BUFx4f_ASAP7_75t_L g1207 ( .A(n_409), .Y(n_1207) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx3_ASAP7_75t_L g413 ( .A(n_410), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_413), .A2(n_562), .B1(n_576), .B2(n_581), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_413), .A2(n_797), .B1(n_798), .B2(n_799), .Y(n_796) );
BUFx2_ASAP7_75t_SL g805 ( .A(n_413), .Y(n_805) );
BUFx3_ASAP7_75t_L g882 ( .A(n_413), .Y(n_882) );
INVx2_ASAP7_75t_SL g964 ( .A(n_413), .Y(n_964) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_415), .A2(n_567), .B1(n_573), .B2(n_586), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_415), .A2(n_586), .B1(n_675), .B2(n_679), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g1257 ( .A1(n_415), .A2(n_1203), .B1(n_1243), .B2(n_1254), .Y(n_1257) );
OAI33xp33_ASAP7_75t_L g489 ( .A1(n_416), .A2(n_490), .A3(n_491), .B1(n_495), .B2(n_498), .B3(n_502), .Y(n_489) );
OAI33xp33_ASAP7_75t_L g1192 ( .A1(n_416), .A2(n_1193), .A3(n_1196), .B1(n_1200), .B2(n_1201), .B3(n_1205), .Y(n_1192) );
OAI33xp33_ASAP7_75t_L g1507 ( .A1(n_416), .A2(n_490), .A3(n_1508), .B1(n_1511), .B2(n_1514), .B3(n_1517), .Y(n_1507) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g584 ( .A(n_417), .Y(n_584) );
NAND3xp33_ASAP7_75t_L g608 ( .A(n_417), .B(n_609), .C(n_611), .Y(n_608) );
AOI33xp33_ASAP7_75t_L g760 ( .A1(n_417), .A2(n_761), .A3(n_762), .B1(n_765), .B2(n_769), .B3(n_770), .Y(n_760) );
AND2x4_ASAP7_75t_L g808 ( .A(n_418), .B(n_809), .Y(n_808) );
OAI31xp33_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_438), .A3(n_444), .B(n_452), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_421), .A2(n_897), .B1(n_911), .B2(n_917), .Y(n_920) );
OAI22xp5_ASAP7_75t_L g1011 ( .A1(n_421), .A2(n_1012), .B1(n_1013), .B2(n_1014), .Y(n_1011) );
OAI22xp33_ASAP7_75t_L g1063 ( .A1(n_421), .A2(n_961), .B1(n_1049), .B2(n_1054), .Y(n_1063) );
NAND3xp33_ASAP7_75t_L g638 ( .A(n_422), .B(n_639), .C(n_644), .Y(n_638) );
NAND3xp33_ASAP7_75t_SL g1271 ( .A(n_422), .B(n_1272), .C(n_1274), .Y(n_1271) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g754 ( .A(n_423), .Y(n_754) );
AND2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
AND2x2_ASAP7_75t_L g429 ( .A(n_424), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g844 ( .A(n_424), .B(n_597), .Y(n_844) );
INVx1_ASAP7_75t_L g753 ( .A(n_425), .Y(n_753) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx2_ASAP7_75t_L g1180 ( .A(n_426), .Y(n_1180) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_427), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_431), .B1(n_432), .B2(n_437), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_429), .A2(n_517), .B1(n_518), .B2(n_519), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_429), .A2(n_434), .B1(n_735), .B2(n_738), .Y(n_750) );
AND2x4_ASAP7_75t_L g539 ( .A(n_430), .B(n_443), .Y(n_539) );
AND2x2_ASAP7_75t_L g693 ( .A(n_430), .B(n_443), .Y(n_693) );
AOI22xp33_ASAP7_75t_SL g470 ( .A1(n_431), .A2(n_471), .B1(n_475), .B2(n_477), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_432), .A2(n_692), .B1(n_693), .B2(n_694), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_432), .A2(n_539), .B1(n_1069), .B2(n_1070), .Y(n_1068) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx3_ASAP7_75t_L g518 ( .A(n_434), .Y(n_518) );
INVx2_ASAP7_75t_L g841 ( .A(n_434), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_434), .A2(n_539), .B1(n_933), .B2(n_934), .Y(n_932) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g745 ( .A(n_439), .Y(n_745) );
BUFx3_ASAP7_75t_L g812 ( .A(n_440), .Y(n_812) );
BUFx3_ASAP7_75t_L g1203 ( .A(n_440), .Y(n_1203) );
BUFx6f_ASAP7_75t_L g1261 ( .A(n_440), .Y(n_1261) );
INVx2_ASAP7_75t_SL g889 ( .A(n_441), .Y(n_889) );
BUFx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g643 ( .A(n_442), .Y(n_643) );
INVx1_ASAP7_75t_L g697 ( .A(n_442), .Y(n_697) );
AND2x2_ASAP7_75t_L g641 ( .A(n_443), .B(n_601), .Y(n_641) );
BUFx6f_ASAP7_75t_L g846 ( .A(n_445), .Y(n_846) );
BUFx2_ASAP7_75t_L g887 ( .A(n_445), .Y(n_887) );
AND2x4_ASAP7_75t_L g449 ( .A(n_446), .B(n_450), .Y(n_449) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
CKINVDCx16_ASAP7_75t_R g448 ( .A(n_449), .Y(n_448) );
INVx4_ASAP7_75t_L g544 ( .A(n_449), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_449), .A2(n_744), .B1(n_745), .B2(n_746), .Y(n_743) );
BUFx3_ASAP7_75t_L g595 ( .A(n_450), .Y(n_595) );
BUFx6f_ASAP7_75t_L g767 ( .A(n_450), .Y(n_767) );
INVx2_ASAP7_75t_L g1178 ( .A(n_450), .Y(n_1178) );
OAI31xp33_ASAP7_75t_L g514 ( .A1(n_452), .A2(n_515), .A3(n_520), .B(n_521), .Y(n_514) );
OAI31xp33_ASAP7_75t_L g688 ( .A1(n_452), .A2(n_689), .A3(n_695), .B(n_698), .Y(n_688) );
OAI31xp33_ASAP7_75t_L g1216 ( .A1(n_452), .A2(n_1217), .A3(n_1218), .B(n_1224), .Y(n_1216) );
BUFx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx2_ASAP7_75t_SL g545 ( .A(n_453), .Y(n_545) );
INVx1_ASAP7_75t_L g755 ( .A(n_453), .Y(n_755) );
BUFx3_ASAP7_75t_L g848 ( .A(n_453), .Y(n_848) );
OAI21xp5_ASAP7_75t_L g1270 ( .A1(n_453), .A2(n_1271), .B(n_1278), .Y(n_1270) );
OAI31xp33_ASAP7_75t_L g1492 ( .A1(n_453), .A2(n_1493), .A3(n_1494), .B(n_1498), .Y(n_1492) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OAI31xp33_ASAP7_75t_SL g456 ( .A1(n_457), .A2(n_462), .A3(n_478), .B(n_481), .Y(n_456) );
INVx2_ASAP7_75t_SL g652 ( .A(n_458), .Y(n_652) );
INVx2_ASAP7_75t_SL g852 ( .A(n_458), .Y(n_852) );
INVx1_ASAP7_75t_L g948 ( .A(n_458), .Y(n_948) );
INVx1_ASAP7_75t_L g1076 ( .A(n_458), .Y(n_1076) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OAI22xp33_ASAP7_75t_L g830 ( .A1(n_463), .A2(n_793), .B1(n_806), .B2(n_818), .Y(n_830) );
OAI22xp33_ASAP7_75t_L g909 ( .A1(n_463), .A2(n_896), .B1(n_910), .B2(n_911), .Y(n_909) );
OAI22xp33_ASAP7_75t_L g977 ( .A1(n_463), .A2(n_955), .B1(n_968), .B2(n_978), .Y(n_977) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g1047 ( .A(n_465), .Y(n_1047) );
NAND3xp33_ASAP7_75t_L g550 ( .A(n_466), .B(n_551), .C(n_554), .Y(n_550) );
NAND3xp33_ASAP7_75t_SL g733 ( .A(n_466), .B(n_734), .C(n_737), .Y(n_733) );
NAND3xp33_ASAP7_75t_SL g1501 ( .A(n_466), .B(n_1502), .C(n_1503), .Y(n_1501) );
CKINVDCx8_ASAP7_75t_R g466 ( .A(n_467), .Y(n_466) );
CKINVDCx8_ASAP7_75t_R g662 ( .A(n_467), .Y(n_662) );
AOI211xp5_ASAP7_75t_L g1128 ( .A1(n_467), .A2(n_556), .B(n_1129), .C(n_1130), .Y(n_1128) );
NOR3xp33_ASAP7_75t_L g1148 ( .A(n_467), .B(n_1149), .C(n_1152), .Y(n_1148) );
BUFx3_ASAP7_75t_L g556 ( .A(n_468), .Y(n_556) );
INVx2_ASAP7_75t_L g627 ( .A(n_468), .Y(n_627) );
BUFx2_ASAP7_75t_L g655 ( .A(n_468), .Y(n_655) );
BUFx2_ASAP7_75t_L g1165 ( .A(n_468), .Y(n_1165) );
BUFx2_ASAP7_75t_L g1231 ( .A(n_468), .Y(n_1231) );
BUFx2_ASAP7_75t_L g1265 ( .A(n_468), .Y(n_1265) );
INVx1_ASAP7_75t_L g617 ( .A(n_469), .Y(n_617) );
AOI22xp33_ASAP7_75t_SL g526 ( .A1(n_471), .A2(n_475), .B1(n_517), .B2(n_527), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_471), .A2(n_475), .B1(n_738), .B2(n_739), .Y(n_737) );
AOI222xp33_ASAP7_75t_L g1264 ( .A1(n_471), .A2(n_475), .B1(n_1265), .B2(n_1266), .C1(n_1267), .C2(n_1268), .Y(n_1264) );
AOI22xp33_ASAP7_75t_L g1503 ( .A1(n_471), .A2(n_475), .B1(n_1496), .B2(n_1504), .Y(n_1503) );
AND2x4_ASAP7_75t_L g471 ( .A(n_472), .B(n_474), .Y(n_471) );
AND2x2_ASAP7_75t_L g475 ( .A(n_472), .B(n_476), .Y(n_475) );
AND2x4_ASAP7_75t_L g552 ( .A(n_472), .B(n_474), .Y(n_552) );
AND2x2_ASAP7_75t_L g657 ( .A(n_472), .B(n_474), .Y(n_657) );
AND2x4_ASAP7_75t_L g658 ( .A(n_472), .B(n_476), .Y(n_658) );
INVx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g704 ( .A(n_473), .B(n_705), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_475), .A2(n_538), .B1(n_552), .B2(n_553), .Y(n_551) );
AOI32xp33_ASAP7_75t_L g703 ( .A1(n_475), .A2(n_694), .A3(n_704), .B1(n_706), .B2(n_708), .Y(n_703) );
INVx2_ASAP7_75t_SL g660 ( .A(n_479), .Y(n_660) );
BUFx3_ASAP7_75t_L g862 ( .A(n_479), .Y(n_862) );
BUFx2_ASAP7_75t_L g1150 ( .A(n_479), .Y(n_1150) );
INVx2_ASAP7_75t_L g661 ( .A(n_480), .Y(n_661) );
INVx1_ASAP7_75t_L g864 ( .A(n_480), .Y(n_864) );
INVx1_ASAP7_75t_L g940 ( .A(n_480), .Y(n_940) );
OAI31xp33_ASAP7_75t_SL g523 ( .A1(n_481), .A2(n_524), .A3(n_525), .B(n_528), .Y(n_523) );
OAI31xp33_ASAP7_75t_L g546 ( .A1(n_481), .A2(n_547), .A3(n_550), .B(n_557), .Y(n_546) );
OAI21xp5_ASAP7_75t_L g649 ( .A1(n_481), .A2(n_650), .B(n_653), .Y(n_649) );
OAI31xp33_ASAP7_75t_SL g699 ( .A1(n_481), .A2(n_700), .A3(n_701), .B(n_709), .Y(n_699) );
OAI21xp5_ASAP7_75t_L g1262 ( .A1(n_481), .A2(n_1263), .B(n_1269), .Y(n_1262) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_484), .Y(n_481) );
AND2x2_ASAP7_75t_L g741 ( .A(n_482), .B(n_484), .Y(n_741) );
AND2x2_ASAP7_75t_SL g866 ( .A(n_482), .B(n_484), .Y(n_866) );
AND2x2_ASAP7_75t_L g950 ( .A(n_482), .B(n_484), .Y(n_950) );
AND2x4_ASAP7_75t_L g1135 ( .A(n_482), .B(n_484), .Y(n_1135) );
INVx1_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND3x1_ASAP7_75t_L g487 ( .A(n_488), .B(n_514), .C(n_523), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_489), .B(n_505), .Y(n_488) );
BUFx6f_ASAP7_75t_L g953 ( .A(n_490), .Y(n_953) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_497), .A2(n_504), .B1(n_510), .B2(n_512), .Y(n_509) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_500), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g1193 ( .A1(n_500), .A2(n_581), .B1(n_1194), .B2(n_1195), .Y(n_1193) );
OAI22xp5_ASAP7_75t_L g1259 ( .A1(n_500), .A2(n_1013), .B1(n_1245), .B2(n_1255), .Y(n_1259) );
INVx1_ASAP7_75t_L g1000 ( .A(n_507), .Y(n_1000) );
OAI22xp33_ASAP7_75t_L g1085 ( .A1(n_507), .A2(n_1086), .B1(n_1087), .B2(n_1089), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g826 ( .A1(n_510), .A2(n_799), .B1(n_814), .B2(n_827), .Y(n_826) );
OAI22xp5_ASAP7_75t_L g980 ( .A1(n_510), .A2(n_960), .B1(n_974), .B2(n_981), .Y(n_980) );
INVx2_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_511), .Y(n_614) );
INVx3_ASAP7_75t_L g677 ( .A(n_511), .Y(n_677) );
INVx5_ASAP7_75t_L g824 ( .A(n_511), .Y(n_824) );
INVx2_ASAP7_75t_SL g1092 ( .A(n_511), .Y(n_1092) );
OAI22xp5_ASAP7_75t_L g1090 ( .A1(n_512), .A2(n_1091), .B1(n_1092), .B2(n_1093), .Y(n_1090) );
OAI22xp5_ASAP7_75t_L g1250 ( .A1(n_512), .A2(n_565), .B1(n_1251), .B2(n_1252), .Y(n_1250) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_518), .A2(n_538), .B1(n_539), .B2(n_540), .Y(n_537) );
AOI222xp33_ASAP7_75t_L g644 ( .A1(n_518), .A2(n_539), .B1(n_596), .B2(n_645), .C1(n_646), .C2(n_647), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g1219 ( .A1(n_518), .A2(n_693), .B1(n_1220), .B2(n_1221), .Y(n_1219) );
AOI222xp33_ASAP7_75t_L g1272 ( .A1(n_518), .A2(n_596), .B1(n_693), .B2(n_1267), .C1(n_1268), .C2(n_1273), .Y(n_1272) );
AOI22xp33_ASAP7_75t_L g1495 ( .A1(n_518), .A2(n_539), .B1(n_1496), .B2(n_1497), .Y(n_1495) );
INVx1_ASAP7_75t_L g779 ( .A(n_529), .Y(n_779) );
AO22x1_ASAP7_75t_SL g529 ( .A1(n_530), .A2(n_531), .B1(n_663), .B2(n_778), .Y(n_529) );
INVx2_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
XNOR2x1_ASAP7_75t_L g531 ( .A(n_532), .B(n_588), .Y(n_531) );
NAND3xp33_ASAP7_75t_L g533 ( .A(n_534), .B(n_546), .C(n_558), .Y(n_533) );
OAI31xp33_ASAP7_75t_SL g534 ( .A1(n_535), .A2(n_541), .A3(n_543), .B(n_545), .Y(n_534) );
BUFx3_ASAP7_75t_L g838 ( .A(n_539), .Y(n_838) );
INVx1_ASAP7_75t_L g1112 ( .A(n_539), .Y(n_1112) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_540), .B(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g1277 ( .A(n_542), .Y(n_1277) );
OAI21xp5_ASAP7_75t_L g637 ( .A1(n_545), .A2(n_638), .B(n_648), .Y(n_637) );
OAI31xp33_ASAP7_75t_L g929 ( .A1(n_545), .A2(n_930), .A3(n_931), .B(n_935), .Y(n_929) );
OAI31xp33_ASAP7_75t_L g987 ( .A1(n_545), .A2(n_988), .A3(n_994), .B(n_995), .Y(n_987) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g853 ( .A(n_549), .Y(n_853) );
INVx2_ASAP7_75t_L g872 ( .A(n_549), .Y(n_872) );
INVx1_ASAP7_75t_L g949 ( .A(n_549), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_549), .A2(n_652), .B1(n_1104), .B2(n_1105), .Y(n_1132) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_549), .A2(n_652), .B1(n_1146), .B2(n_1147), .Y(n_1145) );
INVx1_ASAP7_75t_L g702 ( .A(n_552), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_552), .A2(n_658), .B1(n_933), .B2(n_945), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_552), .A2(n_658), .B1(n_991), .B2(n_1002), .Y(n_1001) );
AOI22xp33_ASAP7_75t_SL g1078 ( .A1(n_552), .A2(n_658), .B1(n_1069), .B2(n_1079), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g1229 ( .A1(n_552), .A2(n_658), .B1(n_1220), .B2(n_1223), .Y(n_1229) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g724 ( .A(n_556), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_559), .B(n_577), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g1212 ( .A1(n_565), .A2(n_1195), .B1(n_1204), .B2(n_1213), .Y(n_1212) );
INVx3_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_SL g569 ( .A(n_566), .Y(n_569) );
INVx2_ASAP7_75t_SL g1095 ( .A(n_566), .Y(n_1095) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_570), .B1(n_571), .B2(n_573), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_571), .A2(n_677), .B1(n_678), .B2(n_679), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g1094 ( .A1(n_571), .A2(n_1095), .B1(n_1096), .B2(n_1097), .Y(n_1094) );
OAI22xp5_ASAP7_75t_L g1246 ( .A1(n_571), .A2(n_1247), .B1(n_1248), .B2(n_1249), .Y(n_1246) );
BUFx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g1214 ( .A(n_572), .Y(n_1214) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g1013 ( .A(n_582), .Y(n_1013) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND3xp33_ASAP7_75t_L g589 ( .A(n_590), .B(n_637), .C(n_649), .Y(n_589) );
AND4x1_ASAP7_75t_L g590 ( .A(n_591), .B(n_608), .C(n_612), .D(n_628), .Y(n_590) );
NAND3xp33_ASAP7_75t_L g591 ( .A(n_592), .B(n_598), .C(n_606), .Y(n_591) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g1222 ( .A(n_596), .B(n_1223), .Y(n_1222) );
BUFx3_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
BUFx3_ASAP7_75t_L g768 ( .A(n_597), .Y(n_768) );
BUFx6f_ASAP7_75t_L g1109 ( .A(n_597), .Y(n_1109) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g771 ( .A(n_600), .Y(n_771) );
INVx3_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
BUFx6f_ASAP7_75t_L g610 ( .A(n_601), .Y(n_610) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx3_ASAP7_75t_L g764 ( .A(n_602), .Y(n_764) );
HB1xp67_ASAP7_75t_L g1173 ( .A(n_604), .Y(n_1173) );
BUFx3_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g773 ( .A(n_605), .Y(n_773) );
BUFx6f_ASAP7_75t_L g1122 ( .A(n_605), .Y(n_1122) );
INVx1_ASAP7_75t_L g1200 ( .A(n_606), .Y(n_1200) );
INVx2_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_SL g761 ( .A(n_607), .Y(n_761) );
NAND3xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_618), .C(n_620), .Y(n_612) );
BUFx3_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
BUFx12f_ASAP7_75t_L g630 ( .A(n_616), .Y(n_630) );
INVx5_ASAP7_75t_L g720 ( .A(n_616), .Y(n_720) );
INVx1_ASAP7_75t_L g705 ( .A(n_617), .Y(n_705) );
INVx1_ASAP7_75t_L g721 ( .A(n_618), .Y(n_721) );
BUFx3_ASAP7_75t_L g1155 ( .A(n_618), .Y(n_1155) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
BUFx3_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx8_ASAP7_75t_L g716 ( .A(n_624), .Y(n_716) );
BUFx3_ASAP7_75t_L g727 ( .A(n_624), .Y(n_727) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g736 ( .A(n_627), .Y(n_736) );
NAND3xp33_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .C(n_636), .Y(n_628) );
BUFx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
BUFx2_ASAP7_75t_L g1057 ( .A(n_632), .Y(n_1057) );
INVx3_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx3_ASAP7_75t_L g829 ( .A(n_633), .Y(n_829) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_641), .B1(n_642), .B2(n_643), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_640), .A2(n_642), .B1(n_660), .B2(n_661), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_641), .A2(n_1114), .B1(n_1115), .B2(n_1116), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g1274 ( .A1(n_641), .A2(n_1275), .B1(n_1276), .B2(n_1277), .Y(n_1274) );
INVx2_ASAP7_75t_L g847 ( .A(n_643), .Y(n_847) );
INVx1_ASAP7_75t_L g936 ( .A(n_643), .Y(n_936) );
INVx1_ASAP7_75t_L g1225 ( .A(n_643), .Y(n_1225) );
AOI222xp33_ASAP7_75t_L g654 ( .A1(n_645), .A2(n_646), .B1(n_647), .B2(n_655), .C1(n_656), .C2(n_658), .Y(n_654) );
INVx2_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
NAND3xp33_ASAP7_75t_L g653 ( .A(n_654), .B(n_659), .C(n_662), .Y(n_653) );
BUFx3_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
BUFx3_ASAP7_75t_L g858 ( .A(n_657), .Y(n_858) );
BUFx6f_ASAP7_75t_L g859 ( .A(n_658), .Y(n_859) );
INVx1_ASAP7_75t_L g1131 ( .A(n_658), .Y(n_1131) );
AOI22xp33_ASAP7_75t_L g1133 ( .A1(n_660), .A2(n_661), .B1(n_1114), .B2(n_1115), .Y(n_1133) );
INVx2_ASAP7_75t_L g1151 ( .A(n_661), .Y(n_1151) );
NAND3xp33_ASAP7_75t_L g1228 ( .A(n_662), .B(n_1229), .C(n_1230), .Y(n_1228) );
INVx1_ASAP7_75t_L g778 ( .A(n_663), .Y(n_778) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .B1(n_710), .B2(n_777), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NAND3xp33_ASAP7_75t_L g667 ( .A(n_668), .B(n_688), .C(n_699), .Y(n_667) );
NOR2xp33_ASAP7_75t_SL g668 ( .A(n_669), .B(n_683), .Y(n_668) );
INVx2_ASAP7_75t_L g905 ( .A(n_677), .Y(n_905) );
OAI22xp33_ASAP7_75t_SL g1048 ( .A1(n_677), .A2(n_981), .B1(n_1049), .B2(n_1050), .Y(n_1048) );
OAI22xp5_ASAP7_75t_L g1258 ( .A1(n_690), .A2(n_967), .B1(n_1247), .B2(n_1251), .Y(n_1258) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_693), .A2(n_840), .B1(n_875), .B2(n_885), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_693), .A2(n_991), .B1(n_992), .B2(n_993), .Y(n_990) );
INVx2_ASAP7_75t_L g1116 ( .A(n_696), .Y(n_1116) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx3_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVxp67_ASAP7_75t_SL g777 ( .A(n_710), .Y(n_777) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
OR2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_756), .Y(n_711) );
INVx1_ASAP7_75t_L g758 ( .A(n_713), .Y(n_758) );
AOI21xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_717), .B(n_722), .Y(n_713) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g1028 ( .A(n_718), .Y(n_1028) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g1162 ( .A(n_720), .Y(n_1162) );
OAI221xp5_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_725), .B1(n_726), .B2(n_728), .C(n_729), .Y(n_723) );
INVx2_ASAP7_75t_L g1158 ( .A(n_726), .Y(n_1158) );
INVx2_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OAI33xp33_ASAP7_75t_L g1209 ( .A1(n_730), .A2(n_893), .A3(n_1210), .B1(n_1211), .B2(n_1212), .B3(n_1215), .Y(n_1209) );
OAI33xp33_ASAP7_75t_L g1241 ( .A1(n_730), .A2(n_893), .A3(n_1242), .B1(n_1246), .B2(n_1250), .B3(n_1253), .Y(n_1241) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_731), .B(n_742), .Y(n_757) );
OAI31xp33_ASAP7_75t_SL g731 ( .A1(n_732), .A2(n_733), .A3(n_740), .B(n_741), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_739), .B(n_752), .Y(n_751) );
OAI31xp33_ASAP7_75t_L g1226 ( .A1(n_741), .A2(n_1227), .A3(n_1228), .B(n_1232), .Y(n_1226) );
OAI31xp33_ASAP7_75t_SL g1499 ( .A1(n_741), .A2(n_1500), .A3(n_1501), .B(n_1505), .Y(n_1499) );
AO21x1_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_747), .B(n_755), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
NAND3xp33_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .C(n_754), .Y(n_749) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
AOI31xp33_ASAP7_75t_SL g1102 ( .A1(n_755), .A2(n_1103), .A3(n_1106), .B(n_1113), .Y(n_1102) );
AO21x1_ASAP7_75t_L g1184 ( .A1(n_755), .A2(n_1185), .B(n_1186), .Y(n_1184) );
OAI31xp33_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_758), .A3(n_759), .B(n_774), .Y(n_756) );
INVx1_ASAP7_75t_L g776 ( .A(n_760), .Y(n_776) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx2_ASAP7_75t_L g1120 ( .A(n_764), .Y(n_1120) );
INVx1_ASAP7_75t_L g1172 ( .A(n_764), .Y(n_1172) );
INVx2_ASAP7_75t_SL g1183 ( .A(n_764), .Y(n_1183) );
BUFx6f_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_782), .B1(n_1139), .B2(n_1279), .Y(n_780) );
INVx2_ASAP7_75t_SL g781 ( .A(n_782), .Y(n_781) );
XOR2x2_ASAP7_75t_L g782 ( .A(n_783), .B(n_924), .Y(n_782) );
OA21x2_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_867), .B(n_923), .Y(n_783) );
INVx2_ASAP7_75t_SL g784 ( .A(n_785), .Y(n_784) );
OR2x2_ASAP7_75t_L g923 ( .A(n_785), .B(n_868), .Y(n_923) );
NAND3xp33_ASAP7_75t_L g786 ( .A(n_787), .B(n_831), .C(n_849), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_788), .B(n_815), .Y(n_787) );
OAI33xp33_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_790), .A3(n_796), .B1(n_800), .B2(n_807), .B3(n_811), .Y(n_788) );
OAI33xp33_ASAP7_75t_L g912 ( .A1(n_789), .A2(n_913), .A3(n_916), .B1(n_920), .B2(n_921), .B3(n_922), .Y(n_912) );
OAI22xp5_ASAP7_75t_SL g790 ( .A1(n_791), .A2(n_792), .B1(n_793), .B2(n_794), .Y(n_790) );
OAI22xp33_ASAP7_75t_L g817 ( .A1(n_791), .A2(n_804), .B1(n_818), .B2(n_821), .Y(n_817) );
INVx2_ASAP7_75t_SL g915 ( .A(n_792), .Y(n_915) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_794), .A2(n_812), .B1(n_813), .B2(n_814), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g913 ( .A1(n_794), .A2(n_895), .B1(n_910), .B2(n_914), .Y(n_913) );
OAI22xp5_ASAP7_75t_L g922 ( .A1(n_794), .A2(n_902), .B1(n_907), .B2(n_914), .Y(n_922) );
OAI22xp33_ASAP7_75t_L g1006 ( .A1(n_794), .A2(n_1007), .B1(n_1008), .B2(n_1009), .Y(n_1006) );
OAI22xp33_ASAP7_75t_L g1018 ( .A1(n_794), .A2(n_1008), .B1(n_1019), .B2(n_1020), .Y(n_1018) );
INVx6_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx5_ASAP7_75t_L g958 ( .A(n_795), .Y(n_958) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_797), .A2(n_813), .B1(n_824), .B2(n_825), .Y(n_823) );
OAI221xp5_ASAP7_75t_L g1118 ( .A1(n_798), .A2(n_882), .B1(n_1091), .B2(n_1096), .C(n_1119), .Y(n_1118) );
OAI22xp5_ASAP7_75t_L g800 ( .A1(n_801), .A2(n_804), .B1(n_805), .B2(n_806), .Y(n_800) );
INVx2_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx4_ASAP7_75t_L g961 ( .A(n_802), .Y(n_961) );
INVx4_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
OAI33xp33_ASAP7_75t_L g1061 ( .A1(n_807), .A2(n_953), .A3(n_1062), .B1(n_1063), .B2(n_1064), .B3(n_1065), .Y(n_1061) );
INVx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g921 ( .A(n_808), .Y(n_921) );
AOI33xp33_ASAP7_75t_L g1169 ( .A1(n_808), .A2(n_1170), .A3(n_1171), .B1(n_1174), .B2(n_1181), .B3(n_1182), .Y(n_1169) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
OAI33xp33_ASAP7_75t_L g815 ( .A1(n_816), .A2(n_817), .A3(n_823), .B1(n_826), .B2(n_828), .B3(n_830), .Y(n_815) );
OAI33xp33_ASAP7_75t_L g976 ( .A1(n_816), .A2(n_908), .A3(n_977), .B1(n_980), .B2(n_983), .B3(n_984), .Y(n_976) );
OAI33xp33_ASAP7_75t_L g1042 ( .A1(n_816), .A2(n_1043), .A3(n_1048), .B1(n_1051), .B2(n_1056), .B3(n_1058), .Y(n_1042) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVxp67_ASAP7_75t_SL g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g1025 ( .A(n_820), .Y(n_1025) );
INVx1_ASAP7_75t_L g1034 ( .A(n_820), .Y(n_1034) );
INVx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
BUFx3_ASAP7_75t_L g901 ( .A(n_824), .Y(n_901) );
OAI22xp5_ASAP7_75t_L g983 ( .A1(n_824), .A2(n_825), .B1(n_962), .B2(n_975), .Y(n_983) );
INVx8_ASAP7_75t_L g1053 ( .A(n_824), .Y(n_1053) );
OAI22xp5_ASAP7_75t_L g899 ( .A1(n_825), .A2(n_900), .B1(n_901), .B2(n_902), .Y(n_899) );
OAI22xp5_ASAP7_75t_L g1051 ( .A1(n_825), .A2(n_1052), .B1(n_1054), .B2(n_1055), .Y(n_1051) );
OAI22xp5_ASAP7_75t_L g903 ( .A1(n_827), .A2(n_904), .B1(n_906), .B2(n_907), .Y(n_903) );
INVx2_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
CKINVDCx5p33_ASAP7_75t_R g908 ( .A(n_829), .Y(n_908) );
INVx2_ASAP7_75t_L g1031 ( .A(n_829), .Y(n_1031) );
OAI31xp33_ASAP7_75t_L g831 ( .A1(n_832), .A2(n_833), .A3(n_845), .B(n_848), .Y(n_831) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g1015 ( .A1(n_836), .A2(n_1013), .B1(n_1016), .B2(n_1017), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_838), .A2(n_839), .B1(n_840), .B2(n_842), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_839), .A2(n_858), .B1(n_859), .B2(n_860), .Y(n_857) );
INVx2_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx2_ASAP7_75t_L g992 ( .A(n_841), .Y(n_992) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g883 ( .A(n_844), .Y(n_883) );
INVx3_ASAP7_75t_L g989 ( .A(n_844), .Y(n_989) );
AOI211xp5_ASAP7_75t_L g1106 ( .A1(n_844), .A2(n_1107), .B(n_1110), .C(n_1111), .Y(n_1106) );
NOR3xp33_ASAP7_75t_L g1186 ( .A(n_844), .B(n_1187), .C(n_1188), .Y(n_1186) );
OAI31xp33_ASAP7_75t_L g878 ( .A1(n_848), .A2(n_879), .A3(n_886), .B(n_890), .Y(n_878) );
OAI31xp33_ASAP7_75t_SL g1066 ( .A1(n_848), .A2(n_1067), .A3(n_1071), .B(n_1072), .Y(n_1066) );
OAI31xp33_ASAP7_75t_L g849 ( .A1(n_850), .A2(n_854), .A3(n_861), .B(n_865), .Y(n_849) );
INVx2_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
OAI22xp33_ASAP7_75t_L g1032 ( .A1(n_855), .A2(n_1009), .B1(n_1017), .B2(n_1033), .Y(n_1032) );
OAI22xp33_ASAP7_75t_L g1058 ( .A1(n_855), .A2(n_978), .B1(n_1059), .B2(n_1060), .Y(n_1058) );
INVx2_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g943 ( .A(n_856), .Y(n_943) );
INVx1_ASAP7_75t_L g1153 ( .A(n_856), .Y(n_1153) );
INVx2_ASAP7_75t_L g1244 ( .A(n_856), .Y(n_1244) );
INVx1_ASAP7_75t_L g1526 ( .A(n_856), .Y(n_1526) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_858), .A2(n_859), .B1(n_875), .B2(n_876), .Y(n_874) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
OAI31xp33_ASAP7_75t_L g870 ( .A1(n_865), .A2(n_871), .A3(n_873), .B(n_877), .Y(n_870) );
BUFx2_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
NAND3xp33_ASAP7_75t_L g869 ( .A(n_870), .B(n_878), .C(n_891), .Y(n_869) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
OAI221xp5_ASAP7_75t_L g1123 ( .A1(n_882), .A2(n_1089), .B1(n_1101), .B2(n_1124), .C(n_1126), .Y(n_1123) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
NOR2xp33_ASAP7_75t_L g891 ( .A(n_892), .B(n_912), .Y(n_891) );
OAI33xp33_ASAP7_75t_L g892 ( .A1(n_893), .A2(n_894), .A3(n_899), .B1(n_903), .B2(n_908), .B3(n_909), .Y(n_892) );
OAI22xp33_ASAP7_75t_L g894 ( .A1(n_895), .A2(n_896), .B1(n_897), .B2(n_898), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g916 ( .A1(n_900), .A2(n_906), .B1(n_917), .B2(n_919), .Y(n_916) );
INVx2_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
INVx1_ASAP7_75t_L g1168 ( .A(n_908), .Y(n_1168) );
INVx2_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
INVx4_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
OAI33xp33_ASAP7_75t_L g952 ( .A1(n_921), .A2(n_953), .A3(n_954), .B1(n_959), .B2(n_965), .B3(n_971), .Y(n_952) );
OAI33xp33_ASAP7_75t_L g1005 ( .A1(n_921), .A2(n_1006), .A3(n_1010), .B1(n_1011), .B2(n_1015), .B3(n_1018), .Y(n_1005) );
AOI22xp5_ASAP7_75t_L g924 ( .A1(n_925), .A2(n_1036), .B1(n_1037), .B2(n_1138), .Y(n_924) );
INVx1_ASAP7_75t_L g1138 ( .A(n_925), .Y(n_1138) );
AOI22xp5_ASAP7_75t_L g925 ( .A1(n_926), .A2(n_927), .B1(n_985), .B2(n_1035), .Y(n_925) );
INVx2_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
NAND3xp33_ASAP7_75t_L g928 ( .A(n_929), .B(n_937), .C(n_951), .Y(n_928) );
OAI31xp33_ASAP7_75t_L g937 ( .A1(n_938), .A2(n_941), .A3(n_946), .B(n_950), .Y(n_937) );
INVx1_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
HB1xp67_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
OAI22xp33_ASAP7_75t_L g984 ( .A1(n_943), .A2(n_957), .B1(n_970), .B2(n_978), .Y(n_984) );
INVx1_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
OAI31xp33_ASAP7_75t_L g996 ( .A1(n_950), .A2(n_997), .A3(n_998), .B(n_1003), .Y(n_996) );
OAI31xp33_ASAP7_75t_L g1073 ( .A1(n_950), .A2(n_1074), .A3(n_1077), .B(n_1080), .Y(n_1073) );
NOR2xp33_ASAP7_75t_L g951 ( .A(n_952), .B(n_976), .Y(n_951) );
INVx1_ASAP7_75t_L g1170 ( .A(n_953), .Y(n_1170) );
OAI22xp33_ASAP7_75t_L g954 ( .A1(n_955), .A2(n_956), .B1(n_957), .B2(n_958), .Y(n_954) );
OAI22xp33_ASAP7_75t_L g1062 ( .A1(n_956), .A2(n_958), .B1(n_1044), .B2(n_1059), .Y(n_1062) );
OAI22xp5_ASAP7_75t_L g971 ( .A1(n_958), .A2(n_972), .B1(n_974), .B2(n_975), .Y(n_971) );
OAI22xp5_ASAP7_75t_L g1065 ( .A1(n_958), .A2(n_972), .B1(n_1050), .B2(n_1055), .Y(n_1065) );
OAI22xp5_ASAP7_75t_L g959 ( .A1(n_960), .A2(n_961), .B1(n_962), .B2(n_963), .Y(n_959) );
OAI22xp5_ASAP7_75t_L g1064 ( .A1(n_961), .A2(n_969), .B1(n_1045), .B2(n_1060), .Y(n_1064) );
INVx5_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
OAI22xp33_ASAP7_75t_L g965 ( .A1(n_966), .A2(n_968), .B1(n_969), .B2(n_970), .Y(n_965) );
HB1xp67_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
INVx2_ASAP7_75t_L g1125 ( .A(n_967), .Y(n_1125) );
OAI22xp5_ASAP7_75t_L g1205 ( .A1(n_967), .A2(n_1206), .B1(n_1207), .B2(n_1208), .Y(n_1205) );
INVx2_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
INVx3_ASAP7_75t_L g1008 ( .A(n_973), .Y(n_1008) );
OAI22xp33_ASAP7_75t_L g1043 ( .A1(n_978), .A2(n_1044), .B1(n_1045), .B2(n_1046), .Y(n_1043) );
BUFx4f_ASAP7_75t_SL g978 ( .A(n_979), .Y(n_978) );
OAI22xp5_ASAP7_75t_L g1027 ( .A1(n_981), .A2(n_1012), .B1(n_1019), .B2(n_1028), .Y(n_1027) );
OAI22xp5_ASAP7_75t_L g1029 ( .A1(n_981), .A2(n_1014), .B1(n_1020), .B2(n_1030), .Y(n_1029) );
INVx3_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
INVx1_ASAP7_75t_L g1035 ( .A(n_985), .Y(n_1035) );
NAND3xp33_ASAP7_75t_SL g986 ( .A(n_987), .B(n_996), .C(n_1004), .Y(n_986) );
NAND3xp33_ASAP7_75t_L g1218 ( .A(n_989), .B(n_1219), .C(n_1222), .Y(n_1218) );
INVx2_ASAP7_75t_SL g999 ( .A(n_1000), .Y(n_999) );
NOR2xp33_ASAP7_75t_SL g1004 ( .A(n_1005), .B(n_1021), .Y(n_1004) );
OAI22xp33_ASAP7_75t_L g1023 ( .A1(n_1007), .A2(n_1016), .B1(n_1024), .B2(n_1026), .Y(n_1023) );
OAI33xp33_ASAP7_75t_L g1021 ( .A1(n_1022), .A2(n_1023), .A3(n_1027), .B1(n_1029), .B2(n_1031), .B3(n_1032), .Y(n_1021) );
INVx2_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
INVx2_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
AOI22xp5_ASAP7_75t_L g1037 ( .A1(n_1038), .A2(n_1081), .B1(n_1136), .B2(n_1137), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
HB1xp67_ASAP7_75t_L g1136 ( .A(n_1039), .Y(n_1136) );
NAND3xp33_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1066), .C(n_1073), .Y(n_1040) );
NOR2xp33_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1061), .Y(n_1041) );
INVxp67_ASAP7_75t_SL g1046 ( .A(n_1047), .Y(n_1046) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
OAI33xp33_ASAP7_75t_L g1083 ( .A1(n_1056), .A2(n_1084), .A3(n_1085), .B1(n_1090), .B2(n_1094), .B3(n_1098), .Y(n_1083) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1081), .Y(n_1137) );
NOR4xp25_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1102), .C(n_1117), .D(n_1127), .Y(n_1082) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1088), .Y(n_1087) );
INVx1_ASAP7_75t_L g1107 ( .A(n_1108), .Y(n_1107) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
BUFx2_ASAP7_75t_L g1121 ( .A(n_1122), .Y(n_1121) );
INVx3_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
AOI31xp33_ASAP7_75t_L g1127 ( .A1(n_1128), .A2(n_1132), .A3(n_1133), .B(n_1134), .Y(n_1127) );
AO21x1_ASAP7_75t_L g1144 ( .A1(n_1134), .A2(n_1145), .B(n_1148), .Y(n_1144) );
CKINVDCx14_ASAP7_75t_R g1134 ( .A(n_1135), .Y(n_1134) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1139), .Y(n_1279) );
XOR2xp5_ASAP7_75t_L g1139 ( .A(n_1140), .B(n_1237), .Y(n_1139) );
HB1xp67_ASAP7_75t_L g1140 ( .A(n_1141), .Y(n_1140) );
AOI22xp5_ASAP7_75t_L g1141 ( .A1(n_1142), .A2(n_1189), .B1(n_1235), .B2(n_1236), .Y(n_1141) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1142), .Y(n_1236) );
NAND4xp25_ASAP7_75t_SL g1143 ( .A(n_1144), .B(n_1154), .C(n_1169), .D(n_1184), .Y(n_1143) );
AOI33xp33_ASAP7_75t_L g1154 ( .A1(n_1155), .A2(n_1156), .A3(n_1159), .B1(n_1163), .B2(n_1166), .B3(n_1168), .Y(n_1154) );
BUFx2_ASAP7_75t_SL g1157 ( .A(n_1158), .Y(n_1157) );
INVx2_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
BUFx2_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
INVx2_ASAP7_75t_L g1175 ( .A(n_1176), .Y(n_1175) );
INVx2_ASAP7_75t_L g1176 ( .A(n_1177), .Y(n_1176) );
INVx2_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
INVx3_ASAP7_75t_SL g1235 ( .A(n_1189), .Y(n_1235) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1190), .Y(n_1234) );
NAND3xp33_ASAP7_75t_L g1190 ( .A(n_1191), .B(n_1216), .C(n_1226), .Y(n_1190) );
NOR2xp33_ASAP7_75t_L g1191 ( .A(n_1192), .B(n_1209), .Y(n_1191) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_1221), .B(n_1231), .Y(n_1230) );
NAND2xp5_ASAP7_75t_L g1502 ( .A(n_1231), .B(n_1497), .Y(n_1502) );
HB1xp67_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
NAND3xp33_ASAP7_75t_L g1239 ( .A(n_1240), .B(n_1262), .C(n_1270), .Y(n_1239) );
NOR2xp33_ASAP7_75t_L g1240 ( .A(n_1241), .B(n_1256), .Y(n_1240) );
OAI221xp5_ASAP7_75t_L g1280 ( .A1(n_1281), .A2(n_1488), .B1(n_1490), .B2(n_1527), .C(n_1531), .Y(n_1280) );
AND4x1_ASAP7_75t_L g1281 ( .A(n_1282), .B(n_1443), .C(n_1461), .D(n_1477), .Y(n_1281) );
OAI33xp33_ASAP7_75t_L g1282 ( .A1(n_1283), .A2(n_1375), .A3(n_1393), .B1(n_1399), .B2(n_1411), .B3(n_1422), .Y(n_1282) );
OAI211xp5_ASAP7_75t_SL g1283 ( .A1(n_1284), .A2(n_1303), .B(n_1324), .C(n_1356), .Y(n_1283) );
INVx2_ASAP7_75t_L g1377 ( .A(n_1284), .Y(n_1377) );
AOI331xp33_ASAP7_75t_L g1400 ( .A1(n_1284), .A2(n_1305), .A3(n_1370), .B1(n_1398), .B2(n_1401), .B3(n_1403), .C1(n_1404), .Y(n_1400) );
NOR2xp33_ASAP7_75t_L g1435 ( .A(n_1284), .B(n_1326), .Y(n_1435) );
NOR2xp33_ASAP7_75t_L g1478 ( .A(n_1284), .B(n_1306), .Y(n_1478) );
OR2x2_ASAP7_75t_L g1284 ( .A(n_1285), .B(n_1299), .Y(n_1284) );
NAND2xp5_ASAP7_75t_L g1340 ( .A(n_1285), .B(n_1341), .Y(n_1340) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1285), .Y(n_1348) );
INVx2_ASAP7_75t_SL g1369 ( .A(n_1285), .Y(n_1369) );
AND2x2_ASAP7_75t_L g1434 ( .A(n_1285), .B(n_1306), .Y(n_1434) );
NAND2xp5_ASAP7_75t_L g1480 ( .A(n_1285), .B(n_1481), .Y(n_1480) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1286), .B(n_1293), .Y(n_1285) );
AND2x6_ASAP7_75t_L g1287 ( .A(n_1288), .B(n_1289), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1288), .B(n_1292), .Y(n_1291) );
AND2x4_ASAP7_75t_L g1294 ( .A(n_1288), .B(n_1295), .Y(n_1294) );
AND2x6_ASAP7_75t_L g1297 ( .A(n_1288), .B(n_1298), .Y(n_1297) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1288), .B(n_1292), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1373 ( .A(n_1288), .B(n_1292), .Y(n_1373) );
NAND2xp5_ASAP7_75t_L g1489 ( .A(n_1288), .B(n_1295), .Y(n_1489) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1290), .B(n_1296), .Y(n_1295) );
HB1xp67_ASAP7_75t_L g1540 ( .A(n_1295), .Y(n_1540) );
CKINVDCx5p33_ASAP7_75t_R g1341 ( .A(n_1299), .Y(n_1341) );
NAND2xp5_ASAP7_75t_L g1347 ( .A(n_1299), .B(n_1348), .Y(n_1347) );
NAND2xp5_ASAP7_75t_L g1365 ( .A(n_1299), .B(n_1307), .Y(n_1365) );
NAND2xp5_ASAP7_75t_L g1405 ( .A(n_1299), .B(n_1406), .Y(n_1405) );
AOI22xp5_ASAP7_75t_L g1412 ( .A1(n_1299), .A2(n_1391), .B1(n_1413), .B2(n_1416), .Y(n_1412) );
OAI22xp5_ASAP7_75t_L g1452 ( .A1(n_1299), .A2(n_1385), .B1(n_1453), .B2(n_1459), .Y(n_1452) );
AND2x2_ASAP7_75t_L g1469 ( .A(n_1299), .B(n_1336), .Y(n_1469) );
AND2x2_ASAP7_75t_L g1487 ( .A(n_1299), .B(n_1337), .Y(n_1487) );
AND2x4_ASAP7_75t_L g1299 ( .A(n_1300), .B(n_1302), .Y(n_1299) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1305), .B(n_1310), .Y(n_1304) );
O2A1O1Ixp33_ASAP7_75t_SL g1349 ( .A1(n_1305), .A2(n_1350), .B(n_1351), .C(n_1353), .Y(n_1349) );
NAND2xp5_ASAP7_75t_L g1463 ( .A(n_1305), .B(n_1464), .Y(n_1463) );
CKINVDCx14_ASAP7_75t_R g1305 ( .A(n_1306), .Y(n_1305) );
NAND2xp5_ASAP7_75t_L g1382 ( .A(n_1306), .B(n_1311), .Y(n_1382) );
NOR2xp33_ASAP7_75t_L g1384 ( .A(n_1306), .B(n_1385), .Y(n_1384) );
NAND2xp5_ASAP7_75t_L g1389 ( .A(n_1306), .B(n_1345), .Y(n_1389) );
AND2x2_ASAP7_75t_L g1392 ( .A(n_1306), .B(n_1377), .Y(n_1392) );
NAND2xp5_ASAP7_75t_L g1414 ( .A(n_1306), .B(n_1415), .Y(n_1414) );
AND2x2_ASAP7_75t_L g1418 ( .A(n_1306), .B(n_1310), .Y(n_1418) );
AND2x2_ASAP7_75t_L g1449 ( .A(n_1306), .B(n_1369), .Y(n_1449) );
INVx3_ASAP7_75t_L g1306 ( .A(n_1307), .Y(n_1306) );
CKINVDCx5p33_ASAP7_75t_R g1330 ( .A(n_1307), .Y(n_1330) );
NAND2xp5_ASAP7_75t_L g1351 ( .A(n_1307), .B(n_1352), .Y(n_1351) );
OR2x2_ASAP7_75t_L g1379 ( .A(n_1307), .B(n_1380), .Y(n_1379) );
AND2x2_ASAP7_75t_L g1387 ( .A(n_1307), .B(n_1312), .Y(n_1387) );
NAND2xp5_ASAP7_75t_L g1409 ( .A(n_1307), .B(n_1385), .Y(n_1409) );
AND2x4_ASAP7_75t_SL g1307 ( .A(n_1308), .B(n_1309), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_1311), .B(n_1315), .Y(n_1310) );
NAND2xp5_ASAP7_75t_L g1332 ( .A(n_1311), .B(n_1321), .Y(n_1332) );
OR2x2_ASAP7_75t_L g1343 ( .A(n_1311), .B(n_1344), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1363 ( .A(n_1311), .B(n_1364), .Y(n_1363) );
NAND2xp5_ASAP7_75t_L g1402 ( .A(n_1311), .B(n_1358), .Y(n_1402) );
AND2x2_ASAP7_75t_L g1426 ( .A(n_1311), .B(n_1345), .Y(n_1426) );
OR2x2_ASAP7_75t_L g1431 ( .A(n_1311), .B(n_1316), .Y(n_1431) );
OR2x2_ASAP7_75t_L g1442 ( .A(n_1311), .B(n_1327), .Y(n_1442) );
OR2x2_ASAP7_75t_L g1471 ( .A(n_1311), .B(n_1389), .Y(n_1471) );
INVx2_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
OR2x2_ASAP7_75t_L g1326 ( .A(n_1312), .B(n_1327), .Y(n_1326) );
NAND2xp5_ASAP7_75t_L g1350 ( .A(n_1312), .B(n_1321), .Y(n_1350) );
AND2x2_ASAP7_75t_L g1357 ( .A(n_1312), .B(n_1358), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1367 ( .A(n_1312), .B(n_1328), .Y(n_1367) );
OR2x2_ASAP7_75t_L g1380 ( .A(n_1312), .B(n_1317), .Y(n_1380) );
AND2x2_ASAP7_75t_L g1397 ( .A(n_1312), .B(n_1398), .Y(n_1397) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1312), .B(n_1359), .Y(n_1408) );
NAND2xp5_ASAP7_75t_L g1458 ( .A(n_1312), .B(n_1317), .Y(n_1458) );
NOR2xp33_ASAP7_75t_L g1473 ( .A(n_1312), .B(n_1474), .Y(n_1473) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1313), .B(n_1314), .Y(n_1312) );
NOR2xp33_ASAP7_75t_L g1474 ( .A(n_1315), .B(n_1352), .Y(n_1474) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1316), .Y(n_1315) );
OR2x2_ASAP7_75t_L g1316 ( .A(n_1317), .B(n_1320), .Y(n_1316) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1317), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_1317), .B(n_1321), .Y(n_1345) );
AND2x2_ASAP7_75t_L g1317 ( .A(n_1318), .B(n_1319), .Y(n_1317) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
OR2x2_ASAP7_75t_L g1327 ( .A(n_1321), .B(n_1328), .Y(n_1327) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1321), .Y(n_1359) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1321), .Y(n_1364) );
NAND2x1_ASAP7_75t_L g1321 ( .A(n_1322), .B(n_1323), .Y(n_1321) );
AOI221xp5_ASAP7_75t_L g1324 ( .A1(n_1325), .A2(n_1333), .B1(n_1342), .B2(n_1346), .C(n_1349), .Y(n_1324) );
NAND2xp5_ASAP7_75t_L g1325 ( .A(n_1326), .B(n_1329), .Y(n_1325) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1326), .Y(n_1464) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1327), .Y(n_1352) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1328), .B(n_1359), .Y(n_1358) );
NAND2xp5_ASAP7_75t_L g1329 ( .A(n_1330), .B(n_1331), .Y(n_1329) );
OR2x2_ASAP7_75t_L g1395 ( .A(n_1330), .B(n_1332), .Y(n_1395) );
AND2x2_ASAP7_75t_L g1398 ( .A(n_1330), .B(n_1358), .Y(n_1398) );
AND2x2_ASAP7_75t_L g1416 ( .A(n_1330), .B(n_1367), .Y(n_1416) );
OR2x2_ASAP7_75t_L g1428 ( .A(n_1330), .B(n_1347), .Y(n_1428) );
INVx1_ASAP7_75t_L g1441 ( .A(n_1330), .Y(n_1441) );
AND2x2_ASAP7_75t_L g1468 ( .A(n_1330), .B(n_1408), .Y(n_1468) );
AOI22xp5_ASAP7_75t_L g1419 ( .A1(n_1331), .A2(n_1341), .B1(n_1386), .B2(n_1420), .Y(n_1419) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
NAND2xp5_ASAP7_75t_L g1410 ( .A(n_1333), .B(n_1342), .Y(n_1410) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
OR2x2_ASAP7_75t_L g1334 ( .A(n_1335), .B(n_1340), .Y(n_1334) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1336), .Y(n_1335) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1336), .Y(n_1355) );
AND2x2_ASAP7_75t_L g1360 ( .A(n_1336), .B(n_1354), .Y(n_1360) );
NAND2xp5_ASAP7_75t_L g1475 ( .A(n_1336), .B(n_1476), .Y(n_1475) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1337), .Y(n_1370) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1337), .Y(n_1388) );
AND2x2_ASAP7_75t_L g1403 ( .A(n_1337), .B(n_1341), .Y(n_1403) );
NAND2xp5_ASAP7_75t_L g1433 ( .A(n_1337), .B(n_1434), .Y(n_1433) );
NAND2xp5_ASAP7_75t_L g1448 ( .A(n_1337), .B(n_1449), .Y(n_1448) );
NAND2xp5_ASAP7_75t_L g1337 ( .A(n_1338), .B(n_1339), .Y(n_1337) );
OR2x2_ASAP7_75t_L g1368 ( .A(n_1341), .B(n_1369), .Y(n_1368) );
OAI32xp33_ASAP7_75t_L g1381 ( .A1(n_1341), .A2(n_1350), .A3(n_1358), .B1(n_1382), .B2(n_1383), .Y(n_1381) );
HB1xp67_ASAP7_75t_SL g1394 ( .A(n_1341), .Y(n_1394) );
AND2x2_ASAP7_75t_L g1454 ( .A(n_1341), .B(n_1388), .Y(n_1454) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1343), .Y(n_1342) );
OR2x2_ASAP7_75t_L g1482 ( .A(n_1344), .B(n_1382), .Y(n_1482) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
AND2x2_ASAP7_75t_L g1386 ( .A(n_1345), .B(n_1387), .Y(n_1386) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1347), .Y(n_1346) );
INVx1_ASAP7_75t_L g1476 ( .A(n_1347), .Y(n_1476) );
INVx2_ASAP7_75t_L g1354 ( .A(n_1348), .Y(n_1354) );
AOI31xp33_ASAP7_75t_L g1465 ( .A1(n_1348), .A2(n_1425), .A3(n_1466), .B(n_1467), .Y(n_1465) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1350), .Y(n_1391) );
NAND2xp5_ASAP7_75t_L g1401 ( .A(n_1350), .B(n_1402), .Y(n_1401) );
OAI221xp5_ASAP7_75t_L g1411 ( .A1(n_1353), .A2(n_1370), .B1(n_1412), .B2(n_1417), .C(n_1419), .Y(n_1411) );
OR2x2_ASAP7_75t_L g1353 ( .A(n_1354), .B(n_1355), .Y(n_1353) );
OAI221xp5_ASAP7_75t_SL g1375 ( .A1(n_1354), .A2(n_1376), .B1(n_1388), .B2(n_1389), .C(n_1390), .Y(n_1375) );
AND2x2_ASAP7_75t_L g1460 ( .A(n_1354), .B(n_1386), .Y(n_1460) );
AOI221xp5_ASAP7_75t_L g1356 ( .A1(n_1357), .A2(n_1360), .B1(n_1361), .B2(n_1370), .C(n_1371), .Y(n_1356) );
INVx1_ASAP7_75t_L g1484 ( .A(n_1357), .Y(n_1484) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1358), .Y(n_1427) );
NAND2xp5_ASAP7_75t_L g1456 ( .A(n_1358), .B(n_1387), .Y(n_1456) );
OAI22xp33_ASAP7_75t_L g1361 ( .A1(n_1362), .A2(n_1365), .B1(n_1366), .B2(n_1368), .Y(n_1361) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1363), .Y(n_1362) );
INVxp33_ASAP7_75t_L g1366 ( .A(n_1367), .Y(n_1366) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1368), .Y(n_1415) );
INVx2_ASAP7_75t_L g1385 ( .A(n_1369), .Y(n_1385) );
O2A1O1Ixp33_ASAP7_75t_L g1393 ( .A1(n_1369), .A2(n_1394), .B(n_1395), .C(n_1396), .Y(n_1393) );
AND2x2_ASAP7_75t_L g1445 ( .A(n_1369), .B(n_1386), .Y(n_1445) );
INVx1_ASAP7_75t_L g1444 ( .A(n_1370), .Y(n_1444) );
AOI221xp5_ASAP7_75t_L g1477 ( .A1(n_1370), .A2(n_1464), .B1(n_1478), .B2(n_1479), .C(n_1483), .Y(n_1477) );
INVx3_ASAP7_75t_L g1436 ( .A(n_1371), .Y(n_1436) );
AND2x2_ASAP7_75t_L g1371 ( .A(n_1372), .B(n_1374), .Y(n_1371) );
AOI211xp5_ASAP7_75t_L g1376 ( .A1(n_1377), .A2(n_1378), .B(n_1381), .C(n_1386), .Y(n_1376) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
NAND2xp5_ASAP7_75t_L g1421 ( .A(n_1385), .B(n_1403), .Y(n_1421) );
NAND2xp5_ASAP7_75t_L g1390 ( .A(n_1391), .B(n_1392), .Y(n_1390) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1392), .Y(n_1447) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1397), .Y(n_1396) );
NAND2xp5_ASAP7_75t_L g1399 ( .A(n_1400), .B(n_1410), .Y(n_1399) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1403), .Y(n_1439) );
AOI22xp5_ASAP7_75t_L g1453 ( .A1(n_1403), .A2(n_1454), .B1(n_1455), .B2(n_1457), .Y(n_1453) );
INVx1_ASAP7_75t_L g1404 ( .A(n_1405), .Y(n_1404) );
INVxp33_ASAP7_75t_SL g1485 ( .A(n_1406), .Y(n_1485) );
NOR2xp33_ASAP7_75t_L g1406 ( .A(n_1407), .B(n_1409), .Y(n_1406) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1414), .Y(n_1413) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1416), .Y(n_1466) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1421), .Y(n_1420) );
NAND3xp33_ASAP7_75t_L g1422 ( .A(n_1423), .B(n_1429), .C(n_1437), .Y(n_1422) );
INVxp67_ASAP7_75t_L g1423 ( .A(n_1424), .Y(n_1423) );
AOI21xp33_ASAP7_75t_L g1424 ( .A1(n_1425), .A2(n_1427), .B(n_1428), .Y(n_1424) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1426), .Y(n_1425) );
NOR2xp33_ASAP7_75t_L g1450 ( .A(n_1426), .B(n_1451), .Y(n_1450) );
AOI211xp5_ASAP7_75t_L g1429 ( .A1(n_1430), .A2(n_1432), .B(n_1435), .C(n_1436), .Y(n_1429) );
INVx1_ASAP7_75t_L g1430 ( .A(n_1431), .Y(n_1430) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1433), .Y(n_1432) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
NOR2xp33_ASAP7_75t_L g1438 ( .A(n_1439), .B(n_1440), .Y(n_1438) );
OR2x2_ASAP7_75t_L g1440 ( .A(n_1441), .B(n_1442), .Y(n_1440) );
INVx2_ASAP7_75t_L g1451 ( .A(n_1442), .Y(n_1451) );
AOI211xp5_ASAP7_75t_L g1443 ( .A1(n_1444), .A2(n_1445), .B(n_1446), .C(n_1452), .Y(n_1443) );
AOI21xp33_ASAP7_75t_L g1446 ( .A1(n_1447), .A2(n_1448), .B(n_1450), .Y(n_1446) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1456), .Y(n_1455) );
INVx1_ASAP7_75t_L g1457 ( .A(n_1458), .Y(n_1457) );
INVxp33_ASAP7_75t_L g1459 ( .A(n_1460), .Y(n_1459) );
O2A1O1Ixp33_ASAP7_75t_L g1461 ( .A1(n_1462), .A2(n_1465), .B(n_1469), .C(n_1470), .Y(n_1461) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1463), .Y(n_1462) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
AOI21xp5_ASAP7_75t_L g1470 ( .A1(n_1471), .A2(n_1472), .B(n_1475), .Y(n_1470) );
INVxp33_ASAP7_75t_L g1472 ( .A(n_1473), .Y(n_1472) );
INVxp67_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1482), .Y(n_1481) );
AOI21xp33_ASAP7_75t_L g1483 ( .A1(n_1484), .A2(n_1485), .B(n_1486), .Y(n_1483) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1487), .Y(n_1486) );
BUFx2_ASAP7_75t_L g1488 ( .A(n_1489), .Y(n_1488) );
HB1xp67_ASAP7_75t_L g1537 ( .A(n_1491), .Y(n_1537) );
NAND3xp33_ASAP7_75t_SL g1491 ( .A(n_1492), .B(n_1499), .C(n_1506), .Y(n_1491) );
NOR2xp33_ASAP7_75t_L g1506 ( .A(n_1507), .B(n_1520), .Y(n_1506) );
INVx1_ASAP7_75t_L g1527 ( .A(n_1528), .Y(n_1527) );
BUFx3_ASAP7_75t_L g1528 ( .A(n_1529), .Y(n_1528) );
BUFx3_ASAP7_75t_L g1532 ( .A(n_1533), .Y(n_1532) );
BUFx3_ASAP7_75t_L g1533 ( .A(n_1534), .Y(n_1533) );
INVxp33_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
OAI21xp5_ASAP7_75t_L g1538 ( .A1(n_1539), .A2(n_1540), .B(n_1541), .Y(n_1538) );
INVx1_ASAP7_75t_L g1541 ( .A(n_1542), .Y(n_1541) );
endmodule