module fake_jpeg_788_n_183 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_183);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_183;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_38),
.B(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_15),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_42),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_1),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

NAND2x1_ASAP7_75t_SL g52 ( 
.A(n_46),
.B(n_47),
.Y(n_52)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_25),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_50),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_53),
.B(n_56),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_21),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_54),
.B(n_65),
.Y(n_90)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_24),
.B1(n_13),
.B2(n_25),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_33),
.A2(n_25),
.B1(n_20),
.B2(n_27),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_62),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_35),
.A2(n_13),
.B1(n_27),
.B2(n_20),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_29),
.A2(n_23),
.B1(n_12),
.B2(n_22),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_64),
.A2(n_73),
.B(n_74),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_12),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_36),
.A2(n_12),
.B1(n_22),
.B2(n_19),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_68),
.A2(n_69),
.B1(n_81),
.B2(n_16),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_40),
.A2(n_22),
.B1(n_19),
.B2(n_14),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_34),
.B(n_19),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_70),
.B(n_76),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_41),
.A2(n_46),
.B1(n_44),
.B2(n_14),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_32),
.A2(n_14),
.B1(n_28),
.B2(n_16),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_32),
.B(n_1),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_50),
.A2(n_28),
.B1(n_16),
.B2(n_26),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_1),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_2),
.Y(n_91)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

BUFx24_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_43),
.C(n_30),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_56),
.C(n_59),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_91),
.B(n_92),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_3),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_37),
.B1(n_58),
.B2(n_78),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_95),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_60),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_96),
.B(n_97),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_51),
.B(n_55),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_4),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_104),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_60),
.Y(n_100)
);

NOR3xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_26),
.C(n_7),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_67),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_103),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_4),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_52),
.B(n_4),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_5),
.Y(n_121)
);

NAND2x1_ASAP7_75t_SL g106 ( 
.A(n_104),
.B(n_52),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_106),
.A2(n_117),
.B(n_121),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_99),
.A2(n_59),
.B1(n_67),
.B2(n_64),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_99),
.A2(n_74),
.B1(n_73),
.B2(n_81),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_116),
.B1(n_118),
.B2(n_100),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_88),
.C(n_96),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_99),
.A2(n_58),
.B1(n_79),
.B2(n_56),
.Y(n_113)
);

AO21x1_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_117),
.B(n_105),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_102),
.A2(n_30),
.B(n_77),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_78),
.B1(n_77),
.B2(n_26),
.Y(n_118)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_106),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_115),
.Y(n_126)
);

NOR3xp33_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_131),
.C(n_136),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_135),
.B1(n_140),
.B2(n_124),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_119),
.B(n_94),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_132),
.C(n_133),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_130),
.A2(n_139),
.B(n_106),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_94),
.C(n_97),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_89),
.B1(n_102),
.B2(n_90),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_90),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_125),
.B(n_98),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_107),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_95),
.B1(n_84),
.B2(n_86),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_141),
.A2(n_150),
.B(n_139),
.Y(n_155)
);

OAI32xp33_ASAP7_75t_SL g142 ( 
.A1(n_129),
.A2(n_113),
.A3(n_107),
.B1(n_125),
.B2(n_110),
.Y(n_142)
);

AOI221xp5_ASAP7_75t_L g158 ( 
.A1(n_142),
.A2(n_127),
.B1(n_109),
.B2(n_114),
.C(n_87),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_147),
.C(n_148),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_146),
.A2(n_151),
.B1(n_128),
.B2(n_140),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_115),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_133),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_126),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

OA21x2_ASAP7_75t_L g152 ( 
.A1(n_141),
.A2(n_135),
.B(n_130),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_154),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_144),
.B(n_132),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_158),
.Y(n_163)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

OAI322xp33_ASAP7_75t_L g157 ( 
.A1(n_150),
.A2(n_134),
.A3(n_127),
.B1(n_139),
.B2(n_124),
.C1(n_109),
.C2(n_114),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_159),
.C(n_160),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_83),
.C(n_95),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_142),
.A2(n_85),
.B1(n_7),
.B2(n_8),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_142),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_163),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_156),
.B(n_149),
.Y(n_165)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

XNOR2x1_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_152),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_169),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_159),
.C(n_152),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_170),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_161),
.C(n_166),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_171),
.A2(n_143),
.B(n_151),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_168),
.A2(n_155),
.B(n_143),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_167),
.C(n_120),
.Y(n_177)
);

OAI221xp5_ASAP7_75t_L g178 ( 
.A1(n_175),
.A2(n_120),
.B1(n_7),
.B2(n_8),
.C(n_5),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_172),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_176),
.B(n_177),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_178),
.A2(n_5),
.B(n_8),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_179),
.B(n_120),
.C(n_180),
.Y(n_181)
);

BUFx24_ASAP7_75t_SL g182 ( 
.A(n_181),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_182),
.B(n_120),
.Y(n_183)
);


endmodule