module real_jpeg_10647_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_139;
wire n_33;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_1),
.A2(n_36),
.B1(n_37),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_1),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_77),
.Y(n_100)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_3),
.A2(n_36),
.B1(n_37),
.B2(n_54),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_54),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_4),
.A2(n_58),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_4),
.Y(n_64)
);

AOI21xp33_ASAP7_75t_L g72 ( 
.A1(n_4),
.A2(n_46),
.B(n_60),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_4),
.B(n_66),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_4),
.A2(n_28),
.B(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_4),
.B(n_28),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_4),
.A2(n_78),
.B1(n_83),
.B2(n_139),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_4),
.A2(n_45),
.B(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_4),
.B(n_45),
.Y(n_163)
);

BUFx10_ASAP7_75t_L g80 ( 
.A(n_5),
.Y(n_80)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_SL g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_10),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_11),
.A2(n_47),
.B1(n_58),
.B2(n_65),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_11),
.A2(n_36),
.B1(n_37),
.B2(n_47),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_47),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_12),
.A2(n_30),
.B1(n_45),
.B2(n_46),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_12),
.A2(n_30),
.B1(n_36),
.B2(n_37),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_14),
.A2(n_58),
.B1(n_65),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_14),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_68),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_68),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_14),
.A2(n_36),
.B1(n_37),
.B2(n_68),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_15),
.A2(n_36),
.B1(n_37),
.B2(n_40),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_16),
.A2(n_36),
.B1(n_37),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_16),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_114),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_112),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_92),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_21),
.B(n_92),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_69),
.C(n_84),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_22),
.B(n_189),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_55),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_42),
.B2(n_43),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_25),
.B(n_42),
.C(n_55),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_39),
.B2(n_41),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_27),
.A2(n_32),
.B1(n_35),
.B2(n_160),
.Y(n_182)
);

A2O1A1Ixp33_ASAP7_75t_SL g32 ( 
.A1(n_28),
.A2(n_33),
.B(n_34),
.C(n_35),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_33),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_28),
.A2(n_29),
.B1(n_49),
.B2(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_28),
.B(n_52),
.Y(n_167)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_29),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_32),
.A2(n_35),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_32),
.A2(n_35),
.B1(n_128),
.B2(n_130),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_32),
.A2(n_35),
.B1(n_130),
.B2(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_32),
.A2(n_35),
.B1(n_153),
.B2(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_33),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_34),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_35),
.B(n_64),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_36),
.B(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_36),
.B(n_38),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_36),
.B(n_144),
.Y(n_143)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_37),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_39),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_48),
.B1(n_51),
.B2(n_53),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_44),
.A2(n_48),
.B1(n_51),
.B2(n_88),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_49),
.B(n_50),
.C(n_51),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_49),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_45),
.A2(n_46),
.B1(n_59),
.B2(n_60),
.Y(n_62)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_48),
.A2(n_51),
.B1(n_53),
.B2(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_48),
.A2(n_51),
.B1(n_88),
.B2(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_49),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_50),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_51),
.B(n_64),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_63),
.B1(n_66),
.B2(n_67),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_57),
.A2(n_62),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B(n_61),
.C(n_62),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_59),
.Y(n_61)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_59),
.B(n_64),
.C(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_64),
.B(n_83),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_67),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_69),
.A2(n_84),
.B1(n_85),
.B2(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_69),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_74),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_78),
.B1(n_81),
.B2(n_83),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_79),
.B1(n_80),
.B2(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_81),
.B1(n_83),
.B2(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_78),
.A2(n_83),
.B1(n_122),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_78),
.A2(n_83),
.B1(n_124),
.B2(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_78),
.A2(n_83),
.B1(n_155),
.B2(n_170),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_79),
.A2(n_80),
.B1(n_121),
.B2(n_123),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_80),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_89),
.C(n_90),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_86),
.A2(n_87),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_89),
.B(n_90),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_91),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_102),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_101),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_111),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_106),
.B1(n_107),
.B2(n_110),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_104),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_186),
.B(n_191),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_172),
.B(n_185),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_157),
.B(n_171),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_147),
.B(n_156),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_136),
.B(n_146),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_125),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_120),
.B(n_125),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_131),
.B2(n_135),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_126),
.B(n_135),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_129),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_131),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_141),
.B(n_145),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_140),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_148),
.B(n_149),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_150),
.B(n_158),
.Y(n_171)
);

FAx1_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_152),
.CI(n_154),
.CON(n_150),
.SN(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_158),
.Y(n_173)
);

FAx1_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_161),
.CI(n_164),
.CON(n_158),
.SN(n_158)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_163),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_169),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_169),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_173),
.B(n_174),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_179),
.B2(n_180),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_182),
.C(n_183),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_181),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_182),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_187),
.B(n_188),
.Y(n_191)
);


endmodule