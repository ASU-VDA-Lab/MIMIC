module fake_ariane_2606_n_2180 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_499, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_387, n_406, n_117, n_139, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_2, n_462, n_32, n_410, n_379, n_445, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_502, n_166, n_253, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_439, n_222, n_478, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_297, n_503, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_384, n_468, n_61, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_231, n_366, n_234, n_492, n_280, n_215, n_252, n_161, n_454, n_298, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_418, n_223, n_403, n_25, n_83, n_389, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_496, n_76, n_342, n_26, n_246, n_0, n_428, n_159, n_358, n_105, n_30, n_494, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_127, n_2180);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_499;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_387;
input n_406;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_502;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_439;
input n_222;
input n_478;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_297;
input n_503;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_384;
input n_468;
input n_61;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_492;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_418;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_127;

output n_2180;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_1383;
wire n_603;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_690;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_813;
wire n_1985;
wire n_995;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_559;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_661;
wire n_2098;
wire n_1751;
wire n_533;
wire n_1917;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2116;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_1432;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_696;
wire n_1442;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_2087;
wire n_931;
wire n_669;
wire n_1491;
wire n_619;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_1340;
wire n_1240;
wire n_1087;
wire n_632;
wire n_650;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_1578;
wire n_1455;
wire n_836;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_706;
wire n_2120;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2168;
wire n_552;
wire n_670;
wire n_1826;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_677;
wire n_604;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_1156;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_957;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_1708;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2143;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_2173;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_1038;
wire n_1978;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_519;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_2014;
wire n_975;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_1775;
wire n_908;
wire n_788;
wire n_1036;
wire n_2169;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_917;
wire n_1271;
wire n_2096;
wire n_1530;
wire n_631;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_2012;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_1813;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_1003;
wire n_701;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_1344;
wire n_1390;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_1136;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_2148;
wire n_1946;
wire n_933;
wire n_1779;
wire n_954;
wire n_596;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_574;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_937;
wire n_1474;
wire n_2081;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_548;
wire n_523;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_849;
wire n_2095;
wire n_1820;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_311),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_491),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_508),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_106),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_505),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_164),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_479),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_187),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_299),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_319),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_276),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_481),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_90),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_377),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_498),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_303),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_439),
.Y(n_526)
);

BUFx2_ASAP7_75t_SL g527 ( 
.A(n_54),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_97),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_240),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_417),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_392),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_340),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_279),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_291),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_83),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_193),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_212),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_496),
.Y(n_538)
);

BUFx2_ASAP7_75t_SL g539 ( 
.A(n_448),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_11),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_193),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_134),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_434),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_502),
.Y(n_544)
);

CKINVDCx11_ASAP7_75t_R g545 ( 
.A(n_253),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_51),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_396),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_118),
.Y(n_548)
);

CKINVDCx14_ASAP7_75t_R g549 ( 
.A(n_440),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_160),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_56),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_212),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_499),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_395),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_385),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_138),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_501),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_473),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_431),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_472),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_259),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_493),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_318),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_101),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_368),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_23),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_359),
.Y(n_567)
);

CKINVDCx16_ASAP7_75t_R g568 ( 
.A(n_495),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_20),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_258),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_282),
.Y(n_571)
);

INVx1_ASAP7_75t_SL g572 ( 
.A(n_411),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_188),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_437),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_22),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_132),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_363),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_256),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_184),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_485),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_327),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_284),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_217),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_240),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_354),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_129),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_242),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_280),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_145),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_123),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_135),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_88),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_209),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_356),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_140),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_27),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_164),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_190),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_248),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_353),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_160),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_112),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_149),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_321),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_488),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_122),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_326),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_312),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_129),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_390),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_415),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_313),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_370),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_250),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_384),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_477),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_346),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_108),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_208),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_503),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_4),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_92),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_490),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_96),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_198),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_67),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_215),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_252),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_320),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_102),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_500),
.Y(n_631)
);

BUFx10_ASAP7_75t_L g632 ( 
.A(n_123),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_169),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_61),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_143),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_161),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_489),
.Y(n_637)
);

CKINVDCx20_ASAP7_75t_R g638 ( 
.A(n_1),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_494),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_71),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_118),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_215),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_402),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_497),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_3),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_44),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_81),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_0),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_46),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_8),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_165),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_48),
.Y(n_652)
);

CKINVDCx14_ASAP7_75t_R g653 ( 
.A(n_425),
.Y(n_653)
);

CKINVDCx16_ASAP7_75t_R g654 ( 
.A(n_36),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_337),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_372),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_239),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_360),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_170),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_105),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_77),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_350),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_184),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_9),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_29),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_59),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_379),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_339),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_443),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_70),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_176),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_466),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_480),
.Y(n_673)
);

BUFx10_ASAP7_75t_L g674 ( 
.A(n_445),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_4),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_460),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_3),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_241),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_487),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_484),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_409),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_124),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_414),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_30),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_476),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_231),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_272),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_463),
.Y(n_688)
);

BUFx10_ASAP7_75t_L g689 ( 
.A(n_33),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_109),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_482),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_239),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_125),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_206),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_325),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_0),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_128),
.Y(n_697)
);

BUFx10_ASAP7_75t_L g698 ( 
.A(n_478),
.Y(n_698)
);

CKINVDCx16_ASAP7_75t_R g699 ( 
.A(n_307),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_86),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_266),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_133),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_217),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_75),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_171),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_330),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_348),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_113),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_432),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_352),
.Y(n_710)
);

CKINVDCx16_ASAP7_75t_R g711 ( 
.A(n_198),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_86),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_331),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_483),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_122),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_263),
.Y(n_716)
);

INVx1_ASAP7_75t_SL g717 ( 
.A(n_182),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_492),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_486),
.Y(n_719)
);

INVx2_ASAP7_75t_SL g720 ( 
.A(n_450),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_41),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_504),
.Y(n_722)
);

INVx1_ASAP7_75t_SL g723 ( 
.A(n_135),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_545),
.Y(n_724)
);

CKINVDCx16_ASAP7_75t_R g725 ( 
.A(n_654),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_650),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_555),
.Y(n_727)
);

INVxp67_ASAP7_75t_SL g728 ( 
.A(n_624),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_624),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_657),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_657),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_666),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_666),
.Y(n_733)
);

INVxp67_ASAP7_75t_SL g734 ( 
.A(n_690),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_690),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_693),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_650),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_650),
.Y(n_738)
);

CKINVDCx20_ASAP7_75t_R g739 ( 
.A(n_621),
.Y(n_739)
);

CKINVDCx16_ASAP7_75t_R g740 ( 
.A(n_711),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_650),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_546),
.Y(n_742)
);

INVxp67_ASAP7_75t_SL g743 ( 
.A(n_693),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_546),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_550),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_550),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_545),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_621),
.Y(n_748)
);

INVxp67_ASAP7_75t_L g749 ( 
.A(n_601),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_561),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_568),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_515),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_664),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_522),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_528),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_528),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_555),
.Y(n_757)
);

CKINVDCx16_ASAP7_75t_R g758 ( 
.A(n_699),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_600),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_529),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_638),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_549),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_536),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_537),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_551),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_552),
.Y(n_766)
);

INVxp67_ASAP7_75t_SL g767 ( 
.A(n_561),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_570),
.Y(n_768)
);

INVxp67_ASAP7_75t_SL g769 ( 
.A(n_579),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_579),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_575),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_576),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_638),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_578),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_631),
.B(n_1),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_639),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_583),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_586),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_590),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_549),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_598),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_603),
.Y(n_782)
);

CKINVDCx16_ASAP7_75t_R g783 ( 
.A(n_632),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_606),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_527),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_625),
.Y(n_786)
);

CKINVDCx16_ASAP7_75t_R g787 ( 
.A(n_632),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_633),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_635),
.Y(n_789)
);

INVxp67_ASAP7_75t_SL g790 ( 
.A(n_609),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_653),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_653),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_640),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_661),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_532),
.Y(n_795)
);

INVxp67_ASAP7_75t_SL g796 ( 
.A(n_609),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_677),
.Y(n_797)
);

CKINVDCx14_ASAP7_75t_R g798 ( 
.A(n_674),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_682),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_684),
.Y(n_800)
);

INVxp67_ASAP7_75t_SL g801 ( 
.A(n_619),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_626),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_702),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_626),
.Y(n_804)
);

BUFx2_ASAP7_75t_L g805 ( 
.A(n_540),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_540),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_619),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_532),
.Y(n_808)
);

INVxp67_ASAP7_75t_SL g809 ( 
.A(n_670),
.Y(n_809)
);

INVxp67_ASAP7_75t_SL g810 ( 
.A(n_670),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_563),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_671),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_562),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_562),
.Y(n_814)
);

INVxp67_ASAP7_75t_SL g815 ( 
.A(n_671),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_726),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_726),
.Y(n_817)
);

BUFx8_ASAP7_75t_L g818 ( 
.A(n_805),
.Y(n_818)
);

BUFx2_ASAP7_75t_L g819 ( 
.A(n_724),
.Y(n_819)
);

HB1xp67_ASAP7_75t_L g820 ( 
.A(n_724),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_727),
.B(n_712),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_727),
.B(n_712),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_813),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_762),
.B(n_672),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_815),
.B(n_632),
.Y(n_825)
);

OA21x2_ASAP7_75t_L g826 ( 
.A1(n_813),
.A2(n_516),
.B(n_511),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_814),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_737),
.Y(n_828)
);

NOR2x1_ASAP7_75t_L g829 ( 
.A(n_814),
.B(n_639),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_737),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_738),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_757),
.B(n_776),
.Y(n_832)
);

INVx4_ASAP7_75t_L g833 ( 
.A(n_757),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_767),
.B(n_689),
.Y(n_834)
);

NOR2x1_ASAP7_75t_L g835 ( 
.A(n_776),
.B(n_644),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_795),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_769),
.B(n_689),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_728),
.B(n_519),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_SL g839 ( 
.A1(n_739),
.A2(n_692),
.B1(n_567),
.B2(n_594),
.Y(n_839)
);

INVxp67_ASAP7_75t_L g840 ( 
.A(n_755),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_738),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_734),
.B(n_719),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_790),
.B(n_689),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_741),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_741),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_742),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_742),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_744),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_744),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_796),
.B(n_674),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_743),
.B(n_531),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_745),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_801),
.B(n_674),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_745),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_762),
.B(n_698),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_746),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_746),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_780),
.B(n_672),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_750),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_750),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_798),
.B(n_533),
.Y(n_861)
);

AND2x2_ASAP7_75t_SL g862 ( 
.A(n_775),
.B(n_605),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_729),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_770),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_780),
.B(n_534),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_791),
.B(n_710),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_805),
.B(n_809),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_770),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_807),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_730),
.Y(n_870)
);

INVx4_ASAP7_75t_L g871 ( 
.A(n_791),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_752),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_754),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_760),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_830),
.Y(n_875)
);

BUFx2_ASAP7_75t_L g876 ( 
.A(n_818),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_849),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_849),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_830),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_849),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_832),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_862),
.A2(n_759),
.B1(n_751),
.B2(n_758),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_824),
.B(n_792),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_832),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_849),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_862),
.A2(n_759),
.B1(n_751),
.B2(n_567),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_828),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_832),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_828),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_828),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_831),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_831),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_862),
.B(n_792),
.Y(n_893)
);

BUFx6f_ASAP7_75t_SL g894 ( 
.A(n_871),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_841),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_832),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_SL g897 ( 
.A1(n_839),
.A2(n_739),
.B1(n_761),
.B2(n_748),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_831),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_858),
.B(n_785),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_874),
.Y(n_900)
);

BUFx2_ASAP7_75t_L g901 ( 
.A(n_818),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_849),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_863),
.B(n_810),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_866),
.B(n_731),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_874),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_863),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_849),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_850),
.B(n_732),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_850),
.B(n_733),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_853),
.B(n_735),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_844),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_863),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_870),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_844),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_SL g915 ( 
.A(n_818),
.B(n_563),
.Y(n_915)
);

BUFx2_ASAP7_75t_L g916 ( 
.A(n_818),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_870),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_870),
.Y(n_918)
);

NAND2xp33_ASAP7_75t_SL g919 ( 
.A(n_871),
.B(n_594),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_872),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_872),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_844),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_817),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_872),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_845),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_845),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_845),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_872),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_872),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_872),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_873),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_867),
.B(n_736),
.Y(n_932)
);

BUFx2_ASAP7_75t_L g933 ( 
.A(n_819),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_816),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_873),
.Y(n_935)
);

INVx1_ASAP7_75t_SL g936 ( 
.A(n_836),
.Y(n_936)
);

INVxp67_ASAP7_75t_L g937 ( 
.A(n_819),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_840),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_873),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_873),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_816),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_873),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_865),
.B(n_725),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_873),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_867),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_869),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_816),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_841),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_869),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_846),
.Y(n_950)
);

NAND2xp33_ASAP7_75t_SL g951 ( 
.A(n_871),
.B(n_623),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_846),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_823),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_823),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_827),
.Y(n_955)
);

CKINVDCx8_ASAP7_75t_R g956 ( 
.A(n_867),
.Y(n_956)
);

HB1xp67_ASAP7_75t_L g957 ( 
.A(n_867),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_956),
.B(n_871),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_899),
.B(n_853),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_950),
.B(n_834),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_875),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_956),
.B(n_740),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_950),
.B(n_834),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_877),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_877),
.Y(n_965)
);

NOR2xp67_ASAP7_75t_L g966 ( 
.A(n_937),
.B(n_938),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_945),
.B(n_957),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_882),
.B(n_943),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_875),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_933),
.B(n_795),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_934),
.Y(n_971)
);

INVx2_ASAP7_75t_SL g972 ( 
.A(n_933),
.Y(n_972)
);

NOR3xp33_ASAP7_75t_L g973 ( 
.A(n_936),
.B(n_839),
.C(n_811),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_879),
.Y(n_974)
);

NAND3xp33_ASAP7_75t_L g975 ( 
.A(n_893),
.B(n_833),
.C(n_842),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_879),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_893),
.B(n_855),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_895),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_883),
.B(n_825),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_904),
.B(n_825),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_932),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_919),
.B(n_861),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_932),
.B(n_837),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_919),
.B(n_783),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_951),
.B(n_787),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_934),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_951),
.B(n_821),
.Y(n_987)
);

HB1xp67_ASAP7_75t_L g988 ( 
.A(n_903),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_886),
.B(n_808),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_895),
.Y(n_990)
);

NAND2xp33_ASAP7_75t_L g991 ( 
.A(n_877),
.B(n_820),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_952),
.B(n_843),
.Y(n_992)
);

NOR2xp67_ASAP7_75t_L g993 ( 
.A(n_908),
.B(n_747),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_909),
.B(n_808),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_903),
.B(n_837),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_903),
.B(n_843),
.Y(n_996)
);

OR2x6_ASAP7_75t_L g997 ( 
.A(n_876),
.B(n_821),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_948),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_910),
.B(n_811),
.Y(n_999)
);

INVx2_ASAP7_75t_SL g1000 ( 
.A(n_876),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_901),
.B(n_756),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_900),
.B(n_821),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_905),
.B(n_747),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_948),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_901),
.B(n_802),
.Y(n_1005)
);

NOR3xp33_ASAP7_75t_L g1006 ( 
.A(n_897),
.B(n_804),
.C(n_723),
.Y(n_1006)
);

BUFx5_ASAP7_75t_L g1007 ( 
.A(n_920),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_881),
.Y(n_1008)
);

XOR2x2_ASAP7_75t_L g1009 ( 
.A(n_915),
.B(n_748),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_884),
.B(n_888),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_877),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_896),
.B(n_833),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_946),
.B(n_833),
.Y(n_1013)
);

NOR2xp67_ASAP7_75t_L g1014 ( 
.A(n_949),
.B(n_833),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_941),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_953),
.B(n_842),
.Y(n_1016)
);

NAND2xp33_ASAP7_75t_L g1017 ( 
.A(n_877),
.B(n_513),
.Y(n_1017)
);

INVx2_ASAP7_75t_SL g1018 ( 
.A(n_916),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_906),
.B(n_912),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_954),
.B(n_955),
.Y(n_1020)
);

INVxp33_ASAP7_75t_L g1021 ( 
.A(n_916),
.Y(n_1021)
);

NAND2xp33_ASAP7_75t_SL g1022 ( 
.A(n_894),
.B(n_623),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_952),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_941),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_913),
.B(n_821),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_917),
.B(n_838),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_918),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_878),
.B(n_822),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_887),
.Y(n_1029)
);

INVxp67_ASAP7_75t_L g1030 ( 
.A(n_880),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_880),
.B(n_851),
.Y(n_1031)
);

CKINVDCx11_ASAP7_75t_R g1032 ( 
.A(n_878),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_887),
.B(n_826),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_880),
.B(n_822),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_889),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_889),
.B(n_822),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_890),
.B(n_749),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_890),
.B(n_822),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_891),
.B(n_753),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_947),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_891),
.Y(n_1041)
);

AOI221x1_ASAP7_75t_L g1042 ( 
.A1(n_921),
.A2(n_827),
.B1(n_560),
.B2(n_585),
.C(n_580),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_SL g1043 ( 
.A(n_924),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_894),
.B(n_761),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_894),
.B(n_773),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_892),
.B(n_854),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_892),
.Y(n_1047)
);

NAND3xp33_ASAP7_75t_L g1048 ( 
.A(n_928),
.B(n_860),
.C(n_856),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_898),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_898),
.B(n_854),
.Y(n_1050)
);

AO21x1_ASAP7_75t_L g1051 ( 
.A1(n_929),
.A2(n_612),
.B(n_605),
.Y(n_1051)
);

AOI221xp5_ASAP7_75t_L g1052 ( 
.A1(n_930),
.A2(n_692),
.B1(n_806),
.B2(n_717),
.C(n_764),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_878),
.B(n_885),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_911),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_911),
.Y(n_1055)
);

NAND2xp33_ASAP7_75t_L g1056 ( 
.A(n_878),
.B(n_517),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_914),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_914),
.B(n_854),
.Y(n_1058)
);

AND2x2_ASAP7_75t_SL g1059 ( 
.A(n_878),
.B(n_676),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_931),
.B(n_773),
.Y(n_1060)
);

INVxp67_ASAP7_75t_L g1061 ( 
.A(n_935),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_922),
.B(n_854),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_885),
.B(n_676),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_922),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_947),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_925),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_925),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_926),
.B(n_857),
.Y(n_1068)
);

OR2x6_ASAP7_75t_L g1069 ( 
.A(n_926),
.B(n_847),
.Y(n_1069)
);

NAND2xp33_ASAP7_75t_L g1070 ( 
.A(n_885),
.B(n_535),
.Y(n_1070)
);

INVx2_ASAP7_75t_SL g1071 ( 
.A(n_927),
.Y(n_1071)
);

INVxp67_ASAP7_75t_L g1072 ( 
.A(n_939),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_885),
.B(n_902),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_940),
.B(n_857),
.Y(n_1074)
);

OR2x2_ASAP7_75t_SL g1075 ( 
.A(n_942),
.B(n_763),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_927),
.Y(n_1076)
);

INVxp33_ASAP7_75t_L g1077 ( 
.A(n_944),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_885),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_902),
.Y(n_1079)
);

INVxp67_ASAP7_75t_L g1080 ( 
.A(n_902),
.Y(n_1080)
);

NOR3xp33_ASAP7_75t_L g1081 ( 
.A(n_902),
.B(n_542),
.C(n_541),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_SL g1082 ( 
.A(n_902),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_907),
.B(n_857),
.Y(n_1083)
);

CKINVDCx20_ASAP7_75t_R g1084 ( 
.A(n_907),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_907),
.B(n_857),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_907),
.B(n_864),
.Y(n_1086)
);

A2O1A1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_907),
.A2(n_864),
.B(n_852),
.C(n_856),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_923),
.B(n_826),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_923),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_923),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_959),
.B(n_864),
.Y(n_1091)
);

AOI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_968),
.A2(n_720),
.B1(n_710),
.B2(n_864),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_988),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_983),
.B(n_847),
.Y(n_1094)
);

INVxp67_ASAP7_75t_L g1095 ( 
.A(n_972),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_989),
.B(n_548),
.Y(n_1096)
);

AO22x2_ASAP7_75t_L g1097 ( 
.A1(n_973),
.A2(n_1063),
.B1(n_1009),
.B2(n_1059),
.Y(n_1097)
);

NAND2x1p5_ASAP7_75t_L g1098 ( 
.A(n_1000),
.B(n_852),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_961),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_980),
.B(n_995),
.Y(n_1100)
);

AO22x2_ASAP7_75t_L g1101 ( 
.A1(n_1006),
.A2(n_812),
.B1(n_868),
.B2(n_860),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_996),
.B(n_868),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_986),
.Y(n_1103)
);

OAI221xp5_ASAP7_75t_L g1104 ( 
.A1(n_1052),
.A2(n_556),
.B1(n_569),
.B2(n_566),
.C(n_564),
.Y(n_1104)
);

INVxp67_ASAP7_75t_L g1105 ( 
.A(n_970),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_997),
.Y(n_1106)
);

NAND2x1p5_ASAP7_75t_L g1107 ( 
.A(n_1018),
.B(n_846),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_969),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_974),
.Y(n_1109)
);

AO22x2_ASAP7_75t_L g1110 ( 
.A1(n_987),
.A2(n_797),
.B1(n_799),
.B2(n_794),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_977),
.A2(n_553),
.B(n_607),
.C(n_604),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_976),
.Y(n_1112)
);

OR2x6_ASAP7_75t_SL g1113 ( 
.A(n_1001),
.B(n_599),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1016),
.B(n_848),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_978),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_990),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_998),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1004),
.Y(n_1118)
);

AO22x2_ASAP7_75t_L g1119 ( 
.A1(n_984),
.A2(n_766),
.B1(n_768),
.B2(n_765),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_960),
.B(n_848),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1008),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_1032),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_981),
.B(n_771),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1020),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1015),
.Y(n_1125)
);

NAND2x1p5_ASAP7_75t_L g1126 ( 
.A(n_967),
.B(n_848),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1027),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1024),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1036),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_960),
.B(n_859),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1038),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1040),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1034),
.Y(n_1133)
);

OR2x6_ASAP7_75t_SL g1134 ( 
.A(n_1005),
.B(n_602),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_994),
.B(n_772),
.Y(n_1135)
);

CKINVDCx20_ASAP7_75t_R g1136 ( 
.A(n_1084),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_1043),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1065),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1012),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1013),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1010),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_975),
.A2(n_979),
.B1(n_1069),
.B2(n_1014),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1023),
.Y(n_1143)
);

AO22x2_ASAP7_75t_L g1144 ( 
.A1(n_985),
.A2(n_784),
.B1(n_786),
.B2(n_782),
.Y(n_1144)
);

AO22x2_ASAP7_75t_L g1145 ( 
.A1(n_1042),
.A2(n_789),
.B1(n_793),
.B2(n_788),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1029),
.Y(n_1146)
);

INVx1_ASAP7_75t_SL g1147 ( 
.A(n_1039),
.Y(n_1147)
);

OAI221xp5_ASAP7_75t_L g1148 ( 
.A1(n_999),
.A2(n_573),
.B1(n_589),
.B2(n_587),
.C(n_584),
.Y(n_1148)
);

BUFx4f_ASAP7_75t_L g1149 ( 
.A(n_997),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1035),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1041),
.Y(n_1151)
);

AND3x1_ASAP7_75t_L g1152 ( 
.A(n_1044),
.B(n_777),
.C(n_774),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1047),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_966),
.A2(n_720),
.B1(n_615),
.B2(n_658),
.Y(n_1154)
);

CKINVDCx20_ASAP7_75t_R g1155 ( 
.A(n_1045),
.Y(n_1155)
);

BUFx8_ASAP7_75t_L g1156 ( 
.A(n_1043),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1049),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1055),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1057),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_997),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1064),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1066),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_962),
.Y(n_1163)
);

AOI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1003),
.A2(n_681),
.B1(n_683),
.B2(n_611),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1046),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1050),
.Y(n_1166)
);

AO22x2_ASAP7_75t_L g1167 ( 
.A1(n_982),
.A2(n_779),
.B1(n_781),
.B2(n_778),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1058),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_963),
.B(n_923),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_963),
.B(n_859),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1062),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1068),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1019),
.Y(n_1173)
);

OAI221xp5_ASAP7_75t_L g1174 ( 
.A1(n_1060),
.A2(n_591),
.B1(n_595),
.B2(n_593),
.C(n_592),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1069),
.Y(n_1175)
);

AO22x2_ASAP7_75t_L g1176 ( 
.A1(n_975),
.A2(n_803),
.B1(n_800),
.B2(n_859),
.Y(n_1176)
);

OAI221xp5_ASAP7_75t_L g1177 ( 
.A1(n_993),
.A2(n_596),
.B1(n_618),
.B2(n_614),
.C(n_597),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_992),
.B(n_835),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1067),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1037),
.B(n_835),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1021),
.B(n_829),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_992),
.B(n_622),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1069),
.Y(n_1183)
);

OAI221xp5_ASAP7_75t_L g1184 ( 
.A1(n_1002),
.A2(n_627),
.B1(n_634),
.B2(n_630),
.C(n_628),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1076),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_1026),
.B(n_636),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1054),
.Y(n_1187)
);

OR2x2_ASAP7_75t_L g1188 ( 
.A(n_1075),
.B(n_641),
.Y(n_1188)
);

NAND2x1p5_ASAP7_75t_L g1189 ( 
.A(n_964),
.B(n_829),
.Y(n_1189)
);

OAI221xp5_ASAP7_75t_L g1190 ( 
.A1(n_1022),
.A2(n_642),
.B1(n_647),
.B2(n_646),
.C(n_645),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1071),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1077),
.B(n_648),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1025),
.Y(n_1193)
);

AOI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_958),
.A2(n_706),
.B1(n_685),
.B2(n_923),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1028),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_991),
.A2(n_649),
.B1(n_652),
.B2(n_651),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1048),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1090),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1031),
.B(n_826),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1030),
.B(n_659),
.Y(n_1200)
);

BUFx8_ASAP7_75t_L g1201 ( 
.A(n_1082),
.Y(n_1201)
);

AO22x2_ASAP7_75t_L g1202 ( 
.A1(n_1088),
.A2(n_612),
.B1(n_539),
.B2(n_572),
.Y(n_1202)
);

AOI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1081),
.A2(n_663),
.B1(n_665),
.B2(n_660),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1048),
.Y(n_1204)
);

OR2x6_ASAP7_75t_L g1205 ( 
.A(n_1078),
.B(n_826),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1074),
.Y(n_1206)
);

AO22x2_ASAP7_75t_L g1207 ( 
.A1(n_1088),
.A2(n_668),
.B1(n_707),
.B2(n_644),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1083),
.B(n_675),
.Y(n_1208)
);

HB1xp67_ASAP7_75t_L g1209 ( 
.A(n_1082),
.Y(n_1209)
);

AO22x2_ASAP7_75t_L g1210 ( 
.A1(n_1033),
.A2(n_707),
.B1(n_714),
.B2(n_668),
.Y(n_1210)
);

NAND2x1p5_ASAP7_75t_L g1211 ( 
.A(n_964),
.B(n_817),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1086),
.B(n_678),
.Y(n_1212)
);

AO22x2_ASAP7_75t_L g1213 ( 
.A1(n_1033),
.A2(n_714),
.B1(n_718),
.B2(n_698),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_964),
.B(n_718),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1061),
.B(n_686),
.Y(n_1215)
);

OAI221xp5_ASAP7_75t_L g1216 ( 
.A1(n_1072),
.A2(n_697),
.B1(n_700),
.B2(n_696),
.C(n_694),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1080),
.B(n_703),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1085),
.B(n_704),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1079),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1087),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1051),
.Y(n_1221)
);

OAI221xp5_ASAP7_75t_L g1222 ( 
.A1(n_1017),
.A2(n_715),
.B1(n_716),
.B2(n_708),
.C(n_705),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1007),
.Y(n_1223)
);

NAND2x1p5_ASAP7_75t_L g1224 ( 
.A(n_965),
.B(n_817),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1007),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_965),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1007),
.Y(n_1227)
);

OR2x6_ASAP7_75t_L g1228 ( 
.A(n_965),
.B(n_1011),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1011),
.B(n_721),
.Y(n_1229)
);

INVxp67_ASAP7_75t_L g1230 ( 
.A(n_1056),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1011),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1007),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_1089),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1053),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1089),
.B(n_817),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1089),
.B(n_817),
.Y(n_1236)
);

NAND2x1p5_ASAP7_75t_L g1237 ( 
.A(n_1073),
.B(n_817),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1070),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_989),
.B(n_722),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_988),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_959),
.B(n_510),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_988),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_989),
.B(n_713),
.Y(n_1243)
);

AO22x2_ASAP7_75t_L g1244 ( 
.A1(n_973),
.A2(n_6),
.B1(n_2),
.B2(n_5),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_988),
.Y(n_1245)
);

AO22x2_ASAP7_75t_L g1246 ( 
.A1(n_973),
.A2(n_6),
.B1(n_2),
.B2(n_5),
.Y(n_1246)
);

AO22x2_ASAP7_75t_L g1247 ( 
.A1(n_973),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_1247)
);

NOR2xp67_ASAP7_75t_L g1248 ( 
.A(n_962),
.B(n_512),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_988),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_971),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_988),
.Y(n_1251)
);

NAND2x1p5_ASAP7_75t_L g1252 ( 
.A(n_972),
.B(n_565),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_959),
.B(n_514),
.Y(n_1253)
);

OAI221xp5_ASAP7_75t_L g1254 ( 
.A1(n_989),
.A2(n_521),
.B1(n_523),
.B2(n_520),
.C(n_518),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_971),
.Y(n_1255)
);

INVxp67_ASAP7_75t_L g1256 ( 
.A(n_972),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_988),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_989),
.B(n_709),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1032),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_988),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_988),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_988),
.Y(n_1262)
);

BUFx8_ASAP7_75t_L g1263 ( 
.A(n_972),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_988),
.Y(n_1264)
);

AND2x6_ASAP7_75t_L g1265 ( 
.A(n_961),
.B(n_565),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_988),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_983),
.B(n_7),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_972),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_959),
.B(n_524),
.Y(n_1269)
);

HB1xp67_ASAP7_75t_L g1270 ( 
.A(n_972),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_989),
.B(n_525),
.Y(n_1271)
);

AO22x2_ASAP7_75t_L g1272 ( 
.A1(n_973),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_988),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_959),
.B(n_526),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_959),
.B(n_530),
.Y(n_1275)
);

AO22x2_ASAP7_75t_L g1276 ( 
.A1(n_973),
.A2(n_13),
.B1(n_10),
.B2(n_12),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_988),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_972),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_971),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_988),
.Y(n_1280)
);

AO22x2_ASAP7_75t_L g1281 ( 
.A1(n_973),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_1281)
);

AO22x2_ASAP7_75t_L g1282 ( 
.A1(n_973),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1032),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_988),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1096),
.B(n_538),
.Y(n_1285)
);

NOR2xp67_ASAP7_75t_L g1286 ( 
.A(n_1095),
.B(n_543),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1147),
.B(n_16),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1100),
.B(n_17),
.Y(n_1288)
);

INVx11_ASAP7_75t_L g1289 ( 
.A(n_1201),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1199),
.A2(n_547),
.B(n_544),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1124),
.B(n_17),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1197),
.A2(n_557),
.B(n_554),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1114),
.A2(n_559),
.B(n_558),
.Y(n_1293)
);

AOI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1221),
.A2(n_637),
.B(n_565),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_SL g1295 ( 
.A(n_1163),
.B(n_571),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1160),
.B(n_18),
.Y(n_1296)
);

AOI21xp33_ASAP7_75t_L g1297 ( 
.A1(n_1239),
.A2(n_577),
.B(n_574),
.Y(n_1297)
);

BUFx4f_ASAP7_75t_L g1298 ( 
.A(n_1283),
.Y(n_1298)
);

NOR2xp67_ASAP7_75t_L g1299 ( 
.A(n_1256),
.B(n_581),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1169),
.A2(n_265),
.B(n_264),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1204),
.A2(n_588),
.B(n_582),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_L g1302 ( 
.A(n_1270),
.Y(n_1302)
);

AOI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1176),
.A2(n_1220),
.B(n_1130),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1173),
.A2(n_610),
.B(n_608),
.Y(n_1304)
);

OA22x2_ASAP7_75t_L g1305 ( 
.A1(n_1105),
.A2(n_1164),
.B1(n_1240),
.B2(n_1093),
.Y(n_1305)
);

NAND3xp33_ASAP7_75t_L g1306 ( 
.A(n_1243),
.B(n_616),
.C(n_613),
.Y(n_1306)
);

A2O1A1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1258),
.A2(n_617),
.B(n_629),
.C(n_620),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1135),
.B(n_18),
.Y(n_1308)
);

NAND2x1p5_ASAP7_75t_L g1309 ( 
.A(n_1149),
.B(n_565),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1121),
.Y(n_1310)
);

OAI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1133),
.A2(n_655),
.B(n_643),
.Y(n_1311)
);

AOI22x1_ASAP7_75t_L g1312 ( 
.A1(n_1206),
.A2(n_656),
.B1(n_669),
.B2(n_667),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1140),
.A2(n_1225),
.B(n_1223),
.Y(n_1313)
);

OAI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1091),
.A2(n_679),
.B(n_673),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1271),
.B(n_19),
.Y(n_1315)
);

BUFx6f_ASAP7_75t_L g1316 ( 
.A(n_1228),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1141),
.B(n_19),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1186),
.B(n_20),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1227),
.A2(n_687),
.B(n_680),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1232),
.A2(n_691),
.B(n_688),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1120),
.A2(n_701),
.B(n_695),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1137),
.B(n_21),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1170),
.A2(n_662),
.B(n_637),
.Y(n_1323)
);

O2A1O1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1148),
.A2(n_1174),
.B(n_1111),
.C(n_1241),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1103),
.Y(n_1325)
);

CKINVDCx10_ASAP7_75t_R g1326 ( 
.A(n_1113),
.Y(n_1326)
);

OAI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1129),
.A2(n_21),
.B(n_22),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1139),
.A2(n_662),
.B(n_637),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1278),
.B(n_23),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1099),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_1268),
.B(n_24),
.Y(n_1331)
);

O2A1O1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1253),
.A2(n_26),
.B(n_24),
.C(n_25),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_SL g1333 ( 
.A(n_1226),
.B(n_637),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_SL g1334 ( 
.A(n_1231),
.B(n_662),
.Y(n_1334)
);

BUFx8_ASAP7_75t_L g1335 ( 
.A(n_1283),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1228),
.Y(n_1336)
);

OAI21xp33_ASAP7_75t_L g1337 ( 
.A1(n_1182),
.A2(n_662),
.B(n_25),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1155),
.B(n_26),
.Y(n_1338)
);

AOI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1176),
.A2(n_268),
.B(n_267),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1131),
.A2(n_1166),
.B(n_1165),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1125),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1136),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1168),
.A2(n_270),
.B(n_269),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1254),
.B(n_27),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_1106),
.B(n_28),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1094),
.B(n_28),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1180),
.B(n_29),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1128),
.Y(n_1348)
);

INVx4_ASAP7_75t_L g1349 ( 
.A(n_1283),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1171),
.A2(n_273),
.B(n_271),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1132),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1172),
.A2(n_275),
.B(n_274),
.Y(n_1352)
);

INVxp67_ASAP7_75t_SL g1353 ( 
.A(n_1201),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1237),
.A2(n_278),
.B(n_277),
.Y(n_1354)
);

AOI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1152),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1142),
.A2(n_283),
.B(n_281),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1123),
.B(n_31),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1269),
.A2(n_286),
.B(n_285),
.Y(n_1358)
);

AOI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1167),
.A2(n_288),
.B(n_287),
.Y(n_1359)
);

INVx3_ASAP7_75t_L g1360 ( 
.A(n_1233),
.Y(n_1360)
);

OR2x2_ASAP7_75t_L g1361 ( 
.A(n_1242),
.B(n_32),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1275),
.A2(n_290),
.B(n_289),
.Y(n_1362)
);

O2A1O1Ixp33_ASAP7_75t_L g1363 ( 
.A1(n_1274),
.A2(n_35),
.B(n_33),
.C(n_34),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1108),
.Y(n_1364)
);

OAI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1219),
.A2(n_34),
.B(n_35),
.Y(n_1365)
);

BUFx2_ASAP7_75t_SL g1366 ( 
.A(n_1259),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1208),
.A2(n_293),
.B(n_292),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1212),
.A2(n_295),
.B(n_294),
.Y(n_1368)
);

A2O1A1Ixp33_ASAP7_75t_L g1369 ( 
.A1(n_1092),
.A2(n_38),
.B(n_36),
.C(n_37),
.Y(n_1369)
);

INVx4_ASAP7_75t_L g1370 ( 
.A(n_1122),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1216),
.B(n_37),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_SL g1372 ( 
.A(n_1263),
.B(n_38),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1123),
.B(n_39),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1218),
.A2(n_297),
.B(n_296),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1102),
.A2(n_300),
.B(n_298),
.Y(n_1375)
);

INVx1_ASAP7_75t_SL g1376 ( 
.A(n_1229),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1109),
.B(n_39),
.Y(n_1377)
);

INVx2_ASAP7_75t_SL g1378 ( 
.A(n_1263),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1112),
.B(n_40),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1178),
.A2(n_302),
.B(n_301),
.Y(n_1380)
);

INVx2_ASAP7_75t_SL g1381 ( 
.A(n_1156),
.Y(n_1381)
);

BUFx8_ASAP7_75t_L g1382 ( 
.A(n_1267),
.Y(n_1382)
);

AND2x4_ASAP7_75t_L g1383 ( 
.A(n_1209),
.B(n_40),
.Y(n_1383)
);

INVxp67_ASAP7_75t_SL g1384 ( 
.A(n_1098),
.Y(n_1384)
);

O2A1O1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1222),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_1385)
);

BUFx4f_ASAP7_75t_L g1386 ( 
.A(n_1126),
.Y(n_1386)
);

AOI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1192),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_SL g1388 ( 
.A(n_1156),
.B(n_45),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_SL g1389 ( 
.A(n_1248),
.B(n_45),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_L g1390 ( 
.A(n_1134),
.B(n_46),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1189),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1115),
.B(n_47),
.Y(n_1392)
);

OAI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1195),
.A2(n_49),
.B(n_50),
.Y(n_1393)
);

INVx4_ASAP7_75t_L g1394 ( 
.A(n_1214),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1116),
.B(n_1117),
.Y(n_1395)
);

INVx4_ASAP7_75t_L g1396 ( 
.A(n_1214),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1245),
.B(n_50),
.Y(n_1397)
);

A2O1A1Ixp33_ASAP7_75t_L g1398 ( 
.A1(n_1154),
.A2(n_53),
.B(n_51),
.C(n_52),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1118),
.B(n_52),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1249),
.B(n_53),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1251),
.B(n_54),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1257),
.B(n_55),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1260),
.B(n_55),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1127),
.A2(n_1215),
.B1(n_1193),
.B2(n_1217),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1261),
.B(n_56),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1097),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1238),
.A2(n_305),
.B(n_304),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1230),
.A2(n_308),
.B(n_306),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1138),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1179),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1262),
.B(n_57),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1234),
.A2(n_310),
.B(n_309),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_SL g1413 ( 
.A(n_1107),
.B(n_58),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_SL g1414 ( 
.A(n_1188),
.B(n_1175),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1250),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1235),
.A2(n_315),
.B(n_314),
.Y(n_1416)
);

NOR3xp33_ASAP7_75t_SL g1417 ( 
.A(n_1177),
.B(n_60),
.C(n_61),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1264),
.B(n_60),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1200),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1266),
.B(n_62),
.Y(n_1420)
);

AOI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1101),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_1421)
);

AOI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1236),
.A2(n_317),
.B(n_316),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1143),
.A2(n_323),
.B(n_322),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1146),
.A2(n_328),
.B(n_324),
.Y(n_1424)
);

O2A1O1Ixp33_ASAP7_75t_L g1425 ( 
.A1(n_1104),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1150),
.A2(n_332),
.B(n_329),
.Y(n_1426)
);

A2O1A1Ixp33_ASAP7_75t_L g1427 ( 
.A1(n_1184),
.A2(n_69),
.B(n_66),
.C(n_68),
.Y(n_1427)
);

AOI21xp33_ASAP7_75t_L g1428 ( 
.A1(n_1097),
.A2(n_68),
.B(n_69),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1151),
.Y(n_1429)
);

INVx1_ASAP7_75t_SL g1430 ( 
.A(n_1181),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1273),
.B(n_70),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1153),
.A2(n_1158),
.B(n_1157),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_SL g1433 ( 
.A(n_1183),
.B(n_71),
.Y(n_1433)
);

NAND3xp33_ASAP7_75t_SL g1434 ( 
.A(n_1203),
.B(n_72),
.C(n_73),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1277),
.B(n_72),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1159),
.A2(n_334),
.B(n_333),
.Y(n_1436)
);

AOI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1161),
.A2(n_336),
.B(n_335),
.Y(n_1437)
);

AND2x6_ASAP7_75t_SL g1438 ( 
.A(n_1280),
.B(n_73),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1187),
.A2(n_1191),
.B1(n_1196),
.B2(n_1167),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1162),
.A2(n_341),
.B(n_338),
.Y(n_1440)
);

AOI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1101),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1284),
.B(n_74),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1119),
.B(n_76),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1119),
.B(n_77),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1198),
.A2(n_343),
.B(n_342),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1185),
.B(n_78),
.Y(n_1446)
);

AOI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1144),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_1447)
);

NOR2x1_ASAP7_75t_R g1448 ( 
.A(n_1244),
.B(n_79),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1255),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1144),
.B(n_80),
.Y(n_1450)
);

NOR2x1_ASAP7_75t_L g1451 ( 
.A(n_1190),
.B(n_509),
.Y(n_1451)
);

A2O1A1Ixp33_ASAP7_75t_L g1452 ( 
.A1(n_1194),
.A2(n_83),
.B(n_81),
.C(n_82),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1205),
.A2(n_345),
.B(n_344),
.Y(n_1453)
);

A2O1A1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1279),
.A2(n_85),
.B(n_82),
.C(n_84),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1110),
.B(n_1145),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1110),
.A2(n_87),
.B1(n_84),
.B2(n_85),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1205),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1252),
.B(n_1211),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1224),
.A2(n_349),
.B(n_347),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1244),
.B(n_87),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_1246),
.Y(n_1461)
);

CKINVDCx20_ASAP7_75t_R g1462 ( 
.A(n_1246),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1202),
.B(n_1213),
.Y(n_1463)
);

CKINVDCx14_ASAP7_75t_R g1464 ( 
.A(n_1265),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1202),
.B(n_88),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1265),
.B(n_89),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1247),
.B(n_89),
.Y(n_1467)
);

AOI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1213),
.A2(n_355),
.B(n_351),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1207),
.A2(n_358),
.B(n_357),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1247),
.B(n_90),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1272),
.B(n_91),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1207),
.A2(n_362),
.B(n_361),
.Y(n_1472)
);

OAI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1265),
.A2(n_91),
.B(n_92),
.Y(n_1473)
);

AOI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1272),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1276),
.B(n_93),
.Y(n_1475)
);

A2O1A1Ixp33_ASAP7_75t_L g1476 ( 
.A1(n_1276),
.A2(n_96),
.B(n_94),
.C(n_95),
.Y(n_1476)
);

AOI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1210),
.A2(n_365),
.B(n_364),
.Y(n_1477)
);

OR2x6_ASAP7_75t_L g1478 ( 
.A(n_1281),
.B(n_97),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1281),
.B(n_98),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1282),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_1480)
);

INVx4_ASAP7_75t_L g1481 ( 
.A(n_1282),
.Y(n_1481)
);

OAI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1197),
.A2(n_99),
.B(n_100),
.Y(n_1482)
);

AOI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1199),
.A2(n_367),
.B(n_366),
.Y(n_1483)
);

OAI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1173),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.Y(n_1484)
);

A2O1A1Ixp33_ASAP7_75t_L g1485 ( 
.A1(n_1096),
.A2(n_105),
.B(n_103),
.C(n_104),
.Y(n_1485)
);

CKINVDCx8_ASAP7_75t_R g1486 ( 
.A(n_1283),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1285),
.A2(n_107),
.B1(n_104),
.B2(n_106),
.Y(n_1487)
);

CKINVDCx20_ASAP7_75t_R g1488 ( 
.A(n_1335),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1430),
.B(n_107),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1310),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1298),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1376),
.B(n_108),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1302),
.B(n_109),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1342),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1338),
.B(n_110),
.Y(n_1495)
);

NAND2x1p5_ASAP7_75t_L g1496 ( 
.A(n_1316),
.B(n_369),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1384),
.B(n_110),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1287),
.B(n_111),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1345),
.B(n_111),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1382),
.Y(n_1500)
);

AND2x2_ASAP7_75t_SL g1501 ( 
.A(n_1475),
.B(n_112),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_SL g1502 ( 
.A(n_1315),
.B(n_1386),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_1289),
.Y(n_1503)
);

AOI221x1_ASAP7_75t_L g1504 ( 
.A1(n_1337),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.C(n_116),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1294),
.A2(n_373),
.B(n_371),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_SL g1506 ( 
.A(n_1386),
.B(n_114),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1298),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1382),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1345),
.B(n_115),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1395),
.B(n_116),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1383),
.B(n_117),
.Y(n_1511)
);

BUFx2_ASAP7_75t_L g1512 ( 
.A(n_1394),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1295),
.B(n_117),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1330),
.Y(n_1514)
);

BUFx6f_ASAP7_75t_L g1515 ( 
.A(n_1316),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1364),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_SL g1517 ( 
.A1(n_1390),
.A2(n_1462),
.B1(n_1478),
.B2(n_1480),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1383),
.B(n_1403),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_1335),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1308),
.B(n_119),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_1326),
.Y(n_1521)
);

CKINVDCx20_ASAP7_75t_R g1522 ( 
.A(n_1486),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_SL g1523 ( 
.A(n_1404),
.B(n_119),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1394),
.B(n_374),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1396),
.B(n_120),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1429),
.Y(n_1526)
);

AND3x1_ASAP7_75t_SL g1527 ( 
.A(n_1388),
.B(n_120),
.C(n_121),
.Y(n_1527)
);

BUFx6f_ASAP7_75t_L g1528 ( 
.A(n_1316),
.Y(n_1528)
);

AOI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1344),
.A2(n_125),
.B1(n_121),
.B2(n_124),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1418),
.B(n_126),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1396),
.B(n_1340),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1366),
.Y(n_1532)
);

NAND2x1p5_ASAP7_75t_L g1533 ( 
.A(n_1336),
.B(n_375),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1288),
.B(n_126),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_1481),
.B(n_127),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1318),
.B(n_127),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1449),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1325),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1291),
.B(n_128),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1341),
.Y(n_1540)
);

NOR2xp67_ASAP7_75t_L g1541 ( 
.A(n_1391),
.B(n_1432),
.Y(n_1541)
);

AOI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1371),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1336),
.B(n_376),
.Y(n_1543)
);

CKINVDCx16_ASAP7_75t_R g1544 ( 
.A(n_1370),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_SL g1545 ( 
.A(n_1336),
.B(n_130),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1317),
.B(n_1346),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1360),
.B(n_378),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1348),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1351),
.Y(n_1549)
);

INVxp67_ASAP7_75t_SL g1550 ( 
.A(n_1360),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1409),
.Y(n_1551)
);

NOR2xp33_ASAP7_75t_L g1552 ( 
.A(n_1481),
.B(n_131),
.Y(n_1552)
);

INVx4_ASAP7_75t_L g1553 ( 
.A(n_1349),
.Y(n_1553)
);

AND2x4_ASAP7_75t_L g1554 ( 
.A(n_1391),
.B(n_380),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1347),
.B(n_133),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1446),
.B(n_134),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1410),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1415),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1377),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1461),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1349),
.Y(n_1561)
);

BUFx6f_ASAP7_75t_L g1562 ( 
.A(n_1457),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1379),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1446),
.B(n_1357),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1370),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1435),
.B(n_136),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1475),
.A2(n_140),
.B1(n_137),
.B2(n_139),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1373),
.B(n_139),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1309),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1439),
.B(n_141),
.Y(n_1570)
);

NAND2x1p5_ASAP7_75t_L g1571 ( 
.A(n_1333),
.B(n_381),
.Y(n_1571)
);

INVx3_ASAP7_75t_L g1572 ( 
.A(n_1296),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1455),
.B(n_141),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1296),
.B(n_142),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1303),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1292),
.B(n_142),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1381),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1478),
.A2(n_145),
.B1(n_143),
.B2(n_144),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_1438),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1392),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1399),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1460),
.B(n_144),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1397),
.B(n_1420),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1428),
.A2(n_148),
.B1(n_146),
.B2(n_147),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1400),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1305),
.B(n_146),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1329),
.B(n_147),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_SL g1588 ( 
.A(n_1301),
.B(n_148),
.Y(n_1588)
);

NAND2x1_ASAP7_75t_L g1589 ( 
.A(n_1313),
.B(n_382),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_SL g1590 ( 
.A(n_1311),
.B(n_149),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1401),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1402),
.Y(n_1592)
);

AOI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1434),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1405),
.Y(n_1594)
);

AOI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1467),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1414),
.B(n_153),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1324),
.B(n_153),
.Y(n_1597)
);

NAND2x1_ASAP7_75t_L g1598 ( 
.A(n_1451),
.B(n_383),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1411),
.Y(n_1599)
);

AOI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1471),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_1600)
);

NAND2x1_ASAP7_75t_L g1601 ( 
.A(n_1458),
.B(n_1356),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1322),
.B(n_154),
.Y(n_1602)
);

INVxp67_ASAP7_75t_L g1603 ( 
.A(n_1331),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1361),
.B(n_155),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_SL g1605 ( 
.A(n_1314),
.B(n_156),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1431),
.B(n_1442),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_1378),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1297),
.B(n_157),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1353),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1322),
.B(n_157),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1286),
.B(n_386),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1406),
.B(n_158),
.Y(n_1612)
);

CKINVDCx20_ASAP7_75t_R g1613 ( 
.A(n_1464),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_1417),
.Y(n_1614)
);

BUFx6f_ASAP7_75t_L g1615 ( 
.A(n_1354),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1443),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1299),
.B(n_158),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1444),
.B(n_159),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1483),
.Y(n_1619)
);

NAND2x1_ASAP7_75t_L g1620 ( 
.A(n_1453),
.B(n_387),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1355),
.A2(n_162),
.B1(n_159),
.B2(n_161),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1372),
.B(n_162),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1450),
.B(n_163),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1447),
.B(n_163),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1304),
.B(n_165),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1421),
.B(n_166),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1465),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_SL g1628 ( 
.A(n_1306),
.B(n_166),
.Y(n_1628)
);

AND2x4_ASAP7_75t_L g1629 ( 
.A(n_1334),
.B(n_507),
.Y(n_1629)
);

BUFx12f_ASAP7_75t_L g1630 ( 
.A(n_1448),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1441),
.B(n_167),
.Y(n_1631)
);

AOI22x1_ASAP7_75t_L g1632 ( 
.A1(n_1327),
.A2(n_1365),
.B1(n_1482),
.B2(n_1321),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1307),
.B(n_1463),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1359),
.Y(n_1634)
);

AND3x1_ASAP7_75t_SL g1635 ( 
.A(n_1448),
.B(n_167),
.C(n_168),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1300),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1433),
.B(n_168),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1393),
.B(n_169),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1470),
.B(n_170),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1456),
.A2(n_173),
.B1(n_171),
.B2(n_172),
.Y(n_1640)
);

INVx5_ASAP7_75t_L g1641 ( 
.A(n_1339),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1479),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1413),
.B(n_506),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1474),
.B(n_174),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1425),
.B(n_175),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1385),
.B(n_175),
.Y(n_1646)
);

AOI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1387),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1332),
.Y(n_1648)
);

BUFx12f_ASAP7_75t_L g1649 ( 
.A(n_1484),
.Y(n_1649)
);

INVx8_ASAP7_75t_L g1650 ( 
.A(n_1389),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1485),
.B(n_177),
.Y(n_1651)
);

A2O1A1Ixp33_ASAP7_75t_L g1652 ( 
.A1(n_1363),
.A2(n_180),
.B(n_178),
.C(n_179),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1398),
.B(n_1476),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1419),
.B(n_179),
.Y(n_1654)
);

NAND2x1p5_ASAP7_75t_L g1655 ( 
.A(n_1459),
.B(n_388),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1454),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1369),
.B(n_180),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1452),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1466),
.B(n_1293),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1427),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1312),
.B(n_181),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1319),
.B(n_181),
.Y(n_1662)
);

NAND2x1p5_ASAP7_75t_L g1663 ( 
.A(n_1358),
.B(n_389),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1473),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_1362),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1477),
.B(n_182),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_1320),
.Y(n_1667)
);

AOI22x1_ASAP7_75t_L g1668 ( 
.A1(n_1290),
.A2(n_186),
.B1(n_183),
.B2(n_185),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1468),
.B(n_183),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1375),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1572),
.B(n_1472),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1490),
.Y(n_1672)
);

AOI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1665),
.A2(n_1601),
.B(n_1670),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1518),
.B(n_185),
.Y(n_1674)
);

BUFx12f_ASAP7_75t_L g1675 ( 
.A(n_1519),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1665),
.A2(n_1368),
.B(n_1367),
.Y(n_1676)
);

AND2x4_ASAP7_75t_L g1677 ( 
.A(n_1572),
.B(n_1469),
.Y(n_1677)
);

INVx1_ASAP7_75t_SL g1678 ( 
.A(n_1522),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1583),
.B(n_1603),
.Y(n_1679)
);

AND2x4_ASAP7_75t_L g1680 ( 
.A(n_1515),
.B(n_1416),
.Y(n_1680)
);

AOI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1589),
.A2(n_1408),
.B(n_1374),
.Y(n_1681)
);

NOR2x1_ASAP7_75t_SL g1682 ( 
.A(n_1531),
.B(n_1422),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1514),
.Y(n_1683)
);

AOI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1659),
.A2(n_1323),
.B(n_1343),
.Y(n_1684)
);

INVx2_ASAP7_75t_SL g1685 ( 
.A(n_1491),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1516),
.Y(n_1686)
);

CKINVDCx20_ASAP7_75t_R g1687 ( 
.A(n_1488),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1538),
.Y(n_1688)
);

BUFx12f_ASAP7_75t_L g1689 ( 
.A(n_1503),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_SL g1690 ( 
.A(n_1667),
.B(n_1350),
.Y(n_1690)
);

INVx3_ASAP7_75t_L g1691 ( 
.A(n_1507),
.Y(n_1691)
);

AOI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1641),
.A2(n_1352),
.B(n_1407),
.Y(n_1692)
);

NOR2xp67_ASAP7_75t_SL g1693 ( 
.A(n_1630),
.B(n_1423),
.Y(n_1693)
);

INVxp67_ASAP7_75t_SL g1694 ( 
.A(n_1550),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1526),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1614),
.B(n_186),
.Y(n_1696)
);

INVxp67_ASAP7_75t_L g1697 ( 
.A(n_1494),
.Y(n_1697)
);

A2O1A1Ixp33_ASAP7_75t_L g1698 ( 
.A1(n_1529),
.A2(n_1412),
.B(n_1426),
.C(n_1424),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1501),
.B(n_187),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1537),
.Y(n_1700)
);

CKINVDCx11_ASAP7_75t_R g1701 ( 
.A(n_1613),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1558),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1540),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1548),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1549),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1546),
.B(n_1380),
.Y(n_1706)
);

A2O1A1Ixp33_ASAP7_75t_L g1707 ( 
.A1(n_1529),
.A2(n_1436),
.B(n_1440),
.C(n_1437),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1551),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1495),
.B(n_188),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1557),
.Y(n_1710)
);

INVxp67_ASAP7_75t_L g1711 ( 
.A(n_1489),
.Y(n_1711)
);

BUFx6f_ASAP7_75t_L g1712 ( 
.A(n_1515),
.Y(n_1712)
);

BUFx2_ASAP7_75t_L g1713 ( 
.A(n_1561),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1562),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1606),
.B(n_189),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1562),
.Y(n_1716)
);

NAND2x1p5_ASAP7_75t_L g1717 ( 
.A(n_1553),
.B(n_1515),
.Y(n_1717)
);

A2O1A1Ixp33_ASAP7_75t_SL g1718 ( 
.A1(n_1648),
.A2(n_1445),
.B(n_1328),
.C(n_191),
.Y(n_1718)
);

AOI222xp33_ASAP7_75t_L g1719 ( 
.A1(n_1517),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.C1(n_192),
.C2(n_194),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1517),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1573),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1492),
.B(n_1499),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1580),
.B(n_195),
.Y(n_1723)
);

BUFx2_ASAP7_75t_L g1724 ( 
.A(n_1512),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1573),
.B(n_196),
.Y(n_1725)
);

AOI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1641),
.A2(n_196),
.B(n_197),
.Y(n_1726)
);

OR2x6_ASAP7_75t_L g1727 ( 
.A(n_1650),
.B(n_391),
.Y(n_1727)
);

BUFx6f_ASAP7_75t_L g1728 ( 
.A(n_1528),
.Y(n_1728)
);

NAND2x1p5_ASAP7_75t_L g1729 ( 
.A(n_1553),
.B(n_1528),
.Y(n_1729)
);

O2A1O1Ixp5_ASAP7_75t_L g1730 ( 
.A1(n_1523),
.A2(n_197),
.B(n_199),
.C(n_200),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1585),
.B(n_199),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1649),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1528),
.B(n_201),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1564),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1591),
.B(n_202),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_1521),
.Y(n_1736)
);

OAI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1597),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_1737)
);

INVx2_ASAP7_75t_SL g1738 ( 
.A(n_1532),
.Y(n_1738)
);

BUFx3_ASAP7_75t_L g1739 ( 
.A(n_1565),
.Y(n_1739)
);

BUFx3_ASAP7_75t_L g1740 ( 
.A(n_1500),
.Y(n_1740)
);

OAI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1597),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1616),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1627),
.Y(n_1743)
);

INVxp67_ASAP7_75t_SL g1744 ( 
.A(n_1541),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1592),
.B(n_206),
.Y(n_1745)
);

AOI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1641),
.A2(n_1632),
.B(n_1664),
.Y(n_1746)
);

AND2x6_ASAP7_75t_L g1747 ( 
.A(n_1629),
.B(n_393),
.Y(n_1747)
);

NOR2xp67_ASAP7_75t_L g1748 ( 
.A(n_1497),
.B(n_394),
.Y(n_1748)
);

OR2x6_ASAP7_75t_L g1749 ( 
.A(n_1650),
.B(n_397),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1609),
.B(n_207),
.Y(n_1750)
);

A2O1A1Ixp33_ASAP7_75t_L g1751 ( 
.A1(n_1542),
.A2(n_207),
.B(n_208),
.C(n_209),
.Y(n_1751)
);

CKINVDCx11_ASAP7_75t_R g1752 ( 
.A(n_1508),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_SL g1753 ( 
.A(n_1577),
.B(n_398),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1509),
.B(n_210),
.Y(n_1754)
);

BUFx6f_ASAP7_75t_L g1755 ( 
.A(n_1562),
.Y(n_1755)
);

AOI22xp33_ASAP7_75t_L g1756 ( 
.A1(n_1570),
.A2(n_210),
.B1(n_211),
.B2(n_213),
.Y(n_1756)
);

AOI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1620),
.A2(n_1619),
.B(n_1598),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1618),
.Y(n_1758)
);

AOI22xp33_ASAP7_75t_L g1759 ( 
.A1(n_1653),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_1759)
);

INVxp67_ASAP7_75t_SL g1760 ( 
.A(n_1541),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1594),
.B(n_214),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1575),
.Y(n_1762)
);

BUFx2_ASAP7_75t_L g1763 ( 
.A(n_1607),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1623),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1559),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1563),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1581),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1510),
.Y(n_1768)
);

A2O1A1Ixp33_ASAP7_75t_L g1769 ( 
.A1(n_1542),
.A2(n_216),
.B(n_218),
.C(n_219),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1599),
.B(n_216),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1639),
.B(n_218),
.Y(n_1771)
);

O2A1O1Ixp5_ASAP7_75t_L g1772 ( 
.A1(n_1646),
.A2(n_219),
.B(n_220),
.C(n_221),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1554),
.Y(n_1773)
);

INVxp67_ASAP7_75t_L g1774 ( 
.A(n_1493),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1530),
.B(n_220),
.Y(n_1775)
);

AOI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1634),
.A2(n_221),
.B(n_222),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_1544),
.Y(n_1777)
);

AND2x4_ASAP7_75t_L g1778 ( 
.A(n_1524),
.B(n_222),
.Y(n_1778)
);

BUFx6f_ASAP7_75t_L g1779 ( 
.A(n_1524),
.Y(n_1779)
);

BUFx2_ASAP7_75t_L g1780 ( 
.A(n_1525),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1566),
.B(n_223),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1498),
.B(n_223),
.Y(n_1782)
);

NAND3xp33_ASAP7_75t_L g1783 ( 
.A(n_1647),
.B(n_224),
.C(n_225),
.Y(n_1783)
);

OR2x6_ASAP7_75t_L g1784 ( 
.A(n_1650),
.B(n_1543),
.Y(n_1784)
);

AOI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1535),
.A2(n_1552),
.B1(n_1644),
.B2(n_1600),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1586),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1596),
.Y(n_1787)
);

AOI21xp5_ASAP7_75t_L g1788 ( 
.A1(n_1636),
.A2(n_224),
.B(n_225),
.Y(n_1788)
);

INVx5_ASAP7_75t_L g1789 ( 
.A(n_1569),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1574),
.B(n_226),
.Y(n_1790)
);

NOR2xp67_ASAP7_75t_SL g1791 ( 
.A(n_1638),
.B(n_226),
.Y(n_1791)
);

INVx3_ASAP7_75t_L g1792 ( 
.A(n_1554),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1654),
.B(n_227),
.Y(n_1793)
);

AND2x4_ASAP7_75t_L g1794 ( 
.A(n_1569),
.B(n_227),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1547),
.Y(n_1795)
);

HB1xp67_ASAP7_75t_L g1796 ( 
.A(n_1633),
.Y(n_1796)
);

INVxp67_ASAP7_75t_L g1797 ( 
.A(n_1511),
.Y(n_1797)
);

OAI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1647),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_1798)
);

BUFx6f_ASAP7_75t_L g1799 ( 
.A(n_1547),
.Y(n_1799)
);

AND2x4_ASAP7_75t_L g1800 ( 
.A(n_1543),
.B(n_228),
.Y(n_1800)
);

AOI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1615),
.A2(n_229),
.B(n_230),
.Y(n_1801)
);

OA21x2_ASAP7_75t_L g1802 ( 
.A1(n_1505),
.A2(n_400),
.B(n_399),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1502),
.B(n_231),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1556),
.Y(n_1804)
);

BUFx5_ASAP7_75t_L g1805 ( 
.A(n_1656),
.Y(n_1805)
);

O2A1O1Ixp33_ASAP7_75t_SL g1806 ( 
.A1(n_1587),
.A2(n_232),
.B(n_233),
.C(n_234),
.Y(n_1806)
);

AND2x4_ASAP7_75t_L g1807 ( 
.A(n_1643),
.B(n_1629),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1604),
.B(n_232),
.Y(n_1808)
);

INVx2_ASAP7_75t_SL g1809 ( 
.A(n_1602),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1539),
.Y(n_1810)
);

BUFx6f_ASAP7_75t_L g1811 ( 
.A(n_1611),
.Y(n_1811)
);

NOR2xp33_ASAP7_75t_L g1812 ( 
.A(n_1513),
.B(n_233),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1534),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1568),
.Y(n_1814)
);

BUFx3_ASAP7_75t_L g1815 ( 
.A(n_1610),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1582),
.B(n_234),
.Y(n_1816)
);

NAND2x1p5_ASAP7_75t_L g1817 ( 
.A(n_1506),
.B(n_401),
.Y(n_1817)
);

AND2x4_ASAP7_75t_L g1818 ( 
.A(n_1643),
.B(n_235),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1555),
.B(n_235),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1595),
.B(n_236),
.Y(n_1820)
);

AOI21xp5_ASAP7_75t_L g1821 ( 
.A1(n_1615),
.A2(n_236),
.B(n_237),
.Y(n_1821)
);

OAI21xp5_ASAP7_75t_L g1822 ( 
.A1(n_1576),
.A2(n_237),
.B(n_238),
.Y(n_1822)
);

INVx3_ASAP7_75t_L g1823 ( 
.A(n_1611),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1595),
.B(n_238),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1622),
.B(n_241),
.Y(n_1825)
);

OAI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1600),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_1826)
);

OAI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1593),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1658),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1520),
.Y(n_1829)
);

AOI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1707),
.A2(n_1605),
.B(n_1588),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1722),
.B(n_1578),
.Y(n_1831)
);

A2O1A1Ixp33_ASAP7_75t_L g1832 ( 
.A1(n_1785),
.A2(n_1593),
.B(n_1608),
.C(n_1624),
.Y(n_1832)
);

BUFx6f_ASAP7_75t_L g1833 ( 
.A(n_1779),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1780),
.B(n_1666),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1674),
.B(n_1669),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1734),
.B(n_1536),
.Y(n_1836)
);

A2O1A1Ixp33_ASAP7_75t_L g1837 ( 
.A1(n_1783),
.A2(n_1751),
.B(n_1769),
.C(n_1820),
.Y(n_1837)
);

BUFx2_ASAP7_75t_SL g1838 ( 
.A(n_1779),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1809),
.B(n_1567),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1672),
.Y(n_1840)
);

O2A1O1Ixp5_ASAP7_75t_L g1841 ( 
.A1(n_1798),
.A2(n_1621),
.B(n_1590),
.C(n_1645),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1797),
.B(n_1579),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1683),
.Y(n_1843)
);

INVx2_ASAP7_75t_SL g1844 ( 
.A(n_1740),
.Y(n_1844)
);

NAND2x1p5_ASAP7_75t_L g1845 ( 
.A(n_1739),
.B(n_1545),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1686),
.B(n_1626),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1815),
.B(n_1617),
.Y(n_1847)
);

AND2x4_ASAP7_75t_L g1848 ( 
.A(n_1694),
.B(n_1504),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1713),
.B(n_1631),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1709),
.B(n_1642),
.Y(n_1850)
);

AND2x4_ASAP7_75t_L g1851 ( 
.A(n_1724),
.B(n_1615),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1721),
.B(n_1621),
.Y(n_1852)
);

AND2x4_ASAP7_75t_L g1853 ( 
.A(n_1784),
.B(n_1637),
.Y(n_1853)
);

OA21x2_ASAP7_75t_L g1854 ( 
.A1(n_1746),
.A2(n_1652),
.B(n_1661),
.Y(n_1854)
);

AOI21xp5_ASAP7_75t_L g1855 ( 
.A1(n_1698),
.A2(n_1660),
.B(n_1663),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1762),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1754),
.B(n_1584),
.Y(n_1857)
);

AOI21xp5_ASAP7_75t_L g1858 ( 
.A1(n_1692),
.A2(n_1663),
.B(n_1655),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1699),
.B(n_1560),
.Y(n_1859)
);

NOR2xp33_ASAP7_75t_R g1860 ( 
.A(n_1687),
.B(n_1625),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1695),
.Y(n_1861)
);

O2A1O1Ixp5_ASAP7_75t_L g1862 ( 
.A1(n_1827),
.A2(n_1651),
.B(n_1657),
.C(n_1612),
.Y(n_1862)
);

BUFx6f_ASAP7_75t_L g1863 ( 
.A(n_1779),
.Y(n_1863)
);

INVx3_ASAP7_75t_L g1864 ( 
.A(n_1712),
.Y(n_1864)
);

CKINVDCx9p33_ASAP7_75t_R g1865 ( 
.A(n_1763),
.Y(n_1865)
);

O2A1O1Ixp33_ASAP7_75t_L g1866 ( 
.A1(n_1824),
.A2(n_1628),
.B(n_1662),
.C(n_1487),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1825),
.B(n_1804),
.Y(n_1867)
);

O2A1O1Ixp5_ASAP7_75t_L g1868 ( 
.A1(n_1826),
.A2(n_1527),
.B(n_1635),
.C(n_1668),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1766),
.B(n_1640),
.Y(n_1869)
);

INVx5_ASAP7_75t_L g1870 ( 
.A(n_1747),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1700),
.B(n_1496),
.Y(n_1871)
);

BUFx6f_ASAP7_75t_L g1872 ( 
.A(n_1799),
.Y(n_1872)
);

AND2x4_ASAP7_75t_L g1873 ( 
.A(n_1784),
.B(n_403),
.Y(n_1873)
);

BUFx2_ASAP7_75t_L g1874 ( 
.A(n_1697),
.Y(n_1874)
);

AND2x4_ASAP7_75t_L g1875 ( 
.A(n_1807),
.B(n_1799),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1758),
.B(n_1496),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1765),
.B(n_1533),
.Y(n_1877)
);

O2A1O1Ixp33_ASAP7_75t_L g1878 ( 
.A1(n_1719),
.A2(n_1655),
.B(n_1533),
.C(n_1571),
.Y(n_1878)
);

BUFx6f_ASAP7_75t_L g1879 ( 
.A(n_1799),
.Y(n_1879)
);

AOI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1684),
.A2(n_1571),
.B(n_245),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_1689),
.Y(n_1881)
);

AOI21xp5_ASAP7_75t_L g1882 ( 
.A1(n_1681),
.A2(n_246),
.B(n_247),
.Y(n_1882)
);

OR2x2_ASAP7_75t_L g1883 ( 
.A(n_1679),
.B(n_246),
.Y(n_1883)
);

OA21x2_ASAP7_75t_L g1884 ( 
.A1(n_1673),
.A2(n_247),
.B(n_248),
.Y(n_1884)
);

OAI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1720),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_1885)
);

A2O1A1Ixp33_ASAP7_75t_L g1886 ( 
.A1(n_1812),
.A2(n_249),
.B(n_251),
.C(n_252),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1767),
.B(n_253),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1742),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1764),
.B(n_254),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1743),
.Y(n_1890)
);

OR2x6_ASAP7_75t_L g1891 ( 
.A(n_1727),
.B(n_1749),
.Y(n_1891)
);

NOR2xp67_ASAP7_75t_L g1892 ( 
.A(n_1796),
.B(n_1768),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1786),
.B(n_254),
.Y(n_1893)
);

AND2x4_ASAP7_75t_L g1894 ( 
.A(n_1807),
.B(n_404),
.Y(n_1894)
);

A2O1A1Ixp33_ASAP7_75t_L g1895 ( 
.A1(n_1818),
.A2(n_255),
.B(n_256),
.C(n_257),
.Y(n_1895)
);

O2A1O1Ixp33_ASAP7_75t_L g1896 ( 
.A1(n_1737),
.A2(n_255),
.B(n_257),
.C(n_258),
.Y(n_1896)
);

NAND2x1p5_ASAP7_75t_L g1897 ( 
.A(n_1778),
.B(n_405),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1829),
.B(n_259),
.Y(n_1898)
);

BUFx3_ASAP7_75t_L g1899 ( 
.A(n_1675),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1774),
.B(n_260),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1800),
.B(n_260),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_SL g1902 ( 
.A(n_1777),
.B(n_406),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1703),
.Y(n_1903)
);

O2A1O1Ixp5_ASAP7_75t_L g1904 ( 
.A1(n_1690),
.A2(n_261),
.B(n_262),
.C(n_263),
.Y(n_1904)
);

BUFx4_ASAP7_75t_R g1905 ( 
.A(n_1795),
.Y(n_1905)
);

NOR2xp33_ASAP7_75t_L g1906 ( 
.A(n_1678),
.B(n_261),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1704),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1725),
.B(n_262),
.Y(n_1908)
);

HB1xp67_ASAP7_75t_L g1909 ( 
.A(n_1787),
.Y(n_1909)
);

O2A1O1Ixp33_ASAP7_75t_L g1910 ( 
.A1(n_1741),
.A2(n_407),
.B(n_408),
.C(n_410),
.Y(n_1910)
);

AOI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1676),
.A2(n_412),
.B(n_413),
.Y(n_1911)
);

OA21x2_ASAP7_75t_L g1912 ( 
.A1(n_1757),
.A2(n_416),
.B(n_418),
.Y(n_1912)
);

AOI21xp5_ASAP7_75t_L g1913 ( 
.A1(n_1706),
.A2(n_419),
.B(n_420),
.Y(n_1913)
);

A2O1A1Ixp33_ASAP7_75t_L g1914 ( 
.A1(n_1818),
.A2(n_421),
.B(n_422),
.C(n_423),
.Y(n_1914)
);

INVx1_ASAP7_75t_SL g1915 ( 
.A(n_1691),
.Y(n_1915)
);

NAND2x1p5_ASAP7_75t_L g1916 ( 
.A(n_1778),
.B(n_1789),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1800),
.B(n_424),
.Y(n_1917)
);

NOR2xp67_ASAP7_75t_L g1918 ( 
.A(n_1711),
.B(n_426),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1814),
.B(n_427),
.Y(n_1919)
);

NAND2x1p5_ASAP7_75t_L g1920 ( 
.A(n_1789),
.B(n_1792),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1705),
.Y(n_1921)
);

O2A1O1Ixp33_ASAP7_75t_L g1922 ( 
.A1(n_1806),
.A2(n_428),
.B(n_429),
.C(n_430),
.Y(n_1922)
);

INVx8_ASAP7_75t_L g1923 ( 
.A(n_1727),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1813),
.B(n_433),
.Y(n_1924)
);

BUFx3_ASAP7_75t_L g1925 ( 
.A(n_1738),
.Y(n_1925)
);

A2O1A1Ixp33_ASAP7_75t_L g1926 ( 
.A1(n_1748),
.A2(n_435),
.B(n_436),
.C(n_438),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1810),
.B(n_441),
.Y(n_1927)
);

AOI21xp5_ASAP7_75t_L g1928 ( 
.A1(n_1682),
.A2(n_442),
.B(n_444),
.Y(n_1928)
);

AOI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1744),
.A2(n_446),
.B(n_447),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1828),
.B(n_449),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1733),
.B(n_451),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1733),
.B(n_452),
.Y(n_1932)
);

BUFx3_ASAP7_75t_L g1933 ( 
.A(n_1899),
.Y(n_1933)
);

BUFx4f_ASAP7_75t_SL g1934 ( 
.A(n_1925),
.Y(n_1934)
);

AND2x4_ASAP7_75t_L g1935 ( 
.A(n_1870),
.B(n_1760),
.Y(n_1935)
);

OAI21xp33_ASAP7_75t_SL g1936 ( 
.A1(n_1891),
.A2(n_1793),
.B(n_1732),
.Y(n_1936)
);

BUFx3_ASAP7_75t_L g1937 ( 
.A(n_1844),
.Y(n_1937)
);

OAI22xp5_ASAP7_75t_L g1938 ( 
.A1(n_1832),
.A2(n_1756),
.B1(n_1759),
.B2(n_1822),
.Y(n_1938)
);

NOR2xp33_ASAP7_75t_L g1939 ( 
.A(n_1915),
.B(n_1752),
.Y(n_1939)
);

AOI22xp33_ASAP7_75t_SL g1940 ( 
.A1(n_1870),
.A2(n_1747),
.B1(n_1811),
.B2(n_1753),
.Y(n_1940)
);

OAI22xp5_ASAP7_75t_L g1941 ( 
.A1(n_1837),
.A2(n_1771),
.B1(n_1819),
.B2(n_1808),
.Y(n_1941)
);

AOI222xp33_ASAP7_75t_L g1942 ( 
.A1(n_1859),
.A2(n_1747),
.B1(n_1696),
.B2(n_1715),
.C1(n_1816),
.C2(n_1750),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1909),
.Y(n_1943)
);

INVx2_ASAP7_75t_SL g1944 ( 
.A(n_1874),
.Y(n_1944)
);

HB1xp67_ASAP7_75t_L g1945 ( 
.A(n_1892),
.Y(n_1945)
);

BUFx6f_ASAP7_75t_L g1946 ( 
.A(n_1872),
.Y(n_1946)
);

AOI22xp33_ASAP7_75t_L g1947 ( 
.A1(n_1850),
.A2(n_1791),
.B1(n_1773),
.B2(n_1811),
.Y(n_1947)
);

BUFx6f_ASAP7_75t_L g1948 ( 
.A(n_1872),
.Y(n_1948)
);

HB1xp67_ASAP7_75t_L g1949 ( 
.A(n_1834),
.Y(n_1949)
);

HB1xp67_ASAP7_75t_L g1950 ( 
.A(n_1846),
.Y(n_1950)
);

BUFx8_ASAP7_75t_L g1951 ( 
.A(n_1901),
.Y(n_1951)
);

INVx3_ASAP7_75t_L g1952 ( 
.A(n_1851),
.Y(n_1952)
);

AND2x4_ASAP7_75t_L g1953 ( 
.A(n_1870),
.B(n_1671),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1903),
.Y(n_1954)
);

HB1xp67_ASAP7_75t_L g1955 ( 
.A(n_1848),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1840),
.Y(n_1956)
);

OAI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1895),
.A2(n_1817),
.B1(n_1749),
.B2(n_1775),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1843),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1861),
.Y(n_1959)
);

BUFx4f_ASAP7_75t_SL g1960 ( 
.A(n_1842),
.Y(n_1960)
);

OAI22xp5_ASAP7_75t_L g1961 ( 
.A1(n_1891),
.A2(n_1781),
.B1(n_1770),
.B2(n_1782),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1836),
.B(n_1708),
.Y(n_1962)
);

BUFx4f_ASAP7_75t_SL g1963 ( 
.A(n_1867),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1835),
.B(n_1685),
.Y(n_1964)
);

AOI22xp33_ASAP7_75t_SL g1965 ( 
.A1(n_1923),
.A2(n_1811),
.B1(n_1823),
.B2(n_1805),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1888),
.B(n_1710),
.Y(n_1966)
);

AOI22xp33_ASAP7_75t_L g1967 ( 
.A1(n_1857),
.A2(n_1688),
.B1(n_1702),
.B2(n_1714),
.Y(n_1967)
);

BUFx6f_ASAP7_75t_L g1968 ( 
.A(n_1872),
.Y(n_1968)
);

AOI22xp33_ASAP7_75t_L g1969 ( 
.A1(n_1847),
.A2(n_1716),
.B1(n_1776),
.B2(n_1788),
.Y(n_1969)
);

AOI22xp33_ASAP7_75t_L g1970 ( 
.A1(n_1839),
.A2(n_1671),
.B1(n_1677),
.B2(n_1821),
.Y(n_1970)
);

CKINVDCx5p33_ASAP7_75t_R g1971 ( 
.A(n_1881),
.Y(n_1971)
);

OAI22xp5_ASAP7_75t_L g1972 ( 
.A1(n_1886),
.A2(n_1726),
.B1(n_1803),
.B2(n_1790),
.Y(n_1972)
);

OAI21xp33_ASAP7_75t_L g1973 ( 
.A1(n_1830),
.A2(n_1801),
.B(n_1723),
.Y(n_1973)
);

AOI22xp33_ASAP7_75t_L g1974 ( 
.A1(n_1831),
.A2(n_1677),
.B1(n_1693),
.B2(n_1731),
.Y(n_1974)
);

OAI22xp5_ASAP7_75t_L g1975 ( 
.A1(n_1852),
.A2(n_1794),
.B1(n_1735),
.B2(n_1745),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1907),
.Y(n_1976)
);

OAI21xp5_ASAP7_75t_SL g1977 ( 
.A1(n_1896),
.A2(n_1794),
.B(n_1717),
.Y(n_1977)
);

OAI21xp33_ASAP7_75t_L g1978 ( 
.A1(n_1882),
.A2(n_1761),
.B(n_1680),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1921),
.Y(n_1979)
);

AOI22xp33_ASAP7_75t_L g1980 ( 
.A1(n_1885),
.A2(n_1755),
.B1(n_1805),
.B2(n_1680),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1890),
.Y(n_1981)
);

BUFx2_ASAP7_75t_L g1982 ( 
.A(n_1865),
.Y(n_1982)
);

AOI22xp33_ASAP7_75t_L g1983 ( 
.A1(n_1923),
.A2(n_1755),
.B1(n_1805),
.B2(n_1789),
.Y(n_1983)
);

OAI22xp33_ASAP7_75t_L g1984 ( 
.A1(n_1902),
.A2(n_1728),
.B1(n_1712),
.B2(n_1755),
.Y(n_1984)
);

AOI22xp33_ASAP7_75t_L g1985 ( 
.A1(n_1876),
.A2(n_1805),
.B1(n_1701),
.B2(n_1728),
.Y(n_1985)
);

CKINVDCx5p33_ASAP7_75t_R g1986 ( 
.A(n_1860),
.Y(n_1986)
);

INVx3_ASAP7_75t_SL g1987 ( 
.A(n_1883),
.Y(n_1987)
);

BUFx6f_ASAP7_75t_L g1988 ( 
.A(n_1879),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1856),
.Y(n_1989)
);

OAI22xp5_ASAP7_75t_L g1990 ( 
.A1(n_1908),
.A2(n_1729),
.B1(n_1712),
.B2(n_1728),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1856),
.Y(n_1991)
);

OAI21xp5_ASAP7_75t_L g1992 ( 
.A1(n_1942),
.A2(n_1841),
.B(n_1868),
.Y(n_1992)
);

NOR2xp33_ASAP7_75t_SL g1993 ( 
.A(n_1986),
.B(n_1971),
.Y(n_1993)
);

OAI21x1_ASAP7_75t_SL g1994 ( 
.A1(n_1977),
.A2(n_1855),
.B(n_1878),
.Y(n_1994)
);

NOR2xp33_ASAP7_75t_L g1995 ( 
.A(n_1934),
.B(n_1906),
.Y(n_1995)
);

OAI21xp5_ASAP7_75t_L g1996 ( 
.A1(n_1942),
.A2(n_1922),
.B(n_1904),
.Y(n_1996)
);

BUFx3_ASAP7_75t_L g1997 ( 
.A(n_1933),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1949),
.B(n_1851),
.Y(n_1998)
);

AOI221x1_ASAP7_75t_L g1999 ( 
.A1(n_1973),
.A2(n_1880),
.B1(n_1893),
.B2(n_1898),
.C(n_1887),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1955),
.B(n_1848),
.Y(n_2000)
);

OAI21xp5_ASAP7_75t_L g2001 ( 
.A1(n_1941),
.A2(n_1914),
.B(n_1862),
.Y(n_2001)
);

OAI21xp5_ASAP7_75t_L g2002 ( 
.A1(n_1941),
.A2(n_1910),
.B(n_1866),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1952),
.B(n_1849),
.Y(n_2003)
);

O2A1O1Ixp33_ASAP7_75t_SL g2004 ( 
.A1(n_1944),
.A2(n_1926),
.B(n_1919),
.C(n_1869),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1952),
.B(n_1875),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1956),
.B(n_1875),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1958),
.B(n_1884),
.Y(n_2007)
);

NOR2x1_ASAP7_75t_L g2008 ( 
.A(n_1982),
.B(n_1864),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1959),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1976),
.B(n_1884),
.Y(n_2010)
);

AO32x2_ASAP7_75t_L g2011 ( 
.A1(n_1961),
.A2(n_1871),
.A3(n_1905),
.B1(n_1877),
.B2(n_1900),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1979),
.B(n_1854),
.Y(n_2012)
);

NOR2x1_ASAP7_75t_SL g2013 ( 
.A(n_1977),
.B(n_1838),
.Y(n_2013)
);

AOI211xp5_ASAP7_75t_L g2014 ( 
.A1(n_1938),
.A2(n_1889),
.B(n_1928),
.C(n_1917),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1981),
.B(n_1854),
.Y(n_2015)
);

A2O1A1Ixp33_ASAP7_75t_L g2016 ( 
.A1(n_1936),
.A2(n_1918),
.B(n_1873),
.C(n_1858),
.Y(n_2016)
);

OAI22xp5_ASAP7_75t_L g2017 ( 
.A1(n_1957),
.A2(n_1897),
.B1(n_1916),
.B2(n_1845),
.Y(n_2017)
);

INVx3_ASAP7_75t_L g2018 ( 
.A(n_1953),
.Y(n_2018)
);

AOI22xp33_ASAP7_75t_L g2019 ( 
.A1(n_1967),
.A2(n_1853),
.B1(n_1894),
.B2(n_1924),
.Y(n_2019)
);

OR2x2_ASAP7_75t_L g2020 ( 
.A(n_1950),
.B(n_1853),
.Y(n_2020)
);

NOR2xp33_ASAP7_75t_L g2021 ( 
.A(n_1960),
.B(n_1736),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1989),
.Y(n_2022)
);

OAI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_1961),
.A2(n_1730),
.B(n_1772),
.Y(n_2023)
);

AND2x4_ASAP7_75t_L g2024 ( 
.A(n_1953),
.B(n_1833),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1943),
.Y(n_2025)
);

AOI221xp5_ASAP7_75t_L g2026 ( 
.A1(n_1972),
.A2(n_1927),
.B1(n_1913),
.B2(n_1911),
.C(n_1718),
.Y(n_2026)
);

AOI221xp5_ASAP7_75t_L g2027 ( 
.A1(n_1975),
.A2(n_1932),
.B1(n_1931),
.B2(n_1929),
.C(n_1930),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_2007),
.Y(n_2028)
);

BUFx3_ASAP7_75t_L g2029 ( 
.A(n_1997),
.Y(n_2029)
);

HB1xp67_ASAP7_75t_L g2030 ( 
.A(n_2012),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_2012),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1998),
.B(n_2003),
.Y(n_2032)
);

BUFx2_ASAP7_75t_L g2033 ( 
.A(n_2008),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_2007),
.Y(n_2034)
);

AND2x4_ASAP7_75t_L g2035 ( 
.A(n_2018),
.B(n_2000),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2010),
.Y(n_2036)
);

OAI22xp5_ASAP7_75t_L g2037 ( 
.A1(n_1992),
.A2(n_1963),
.B1(n_1974),
.B2(n_1970),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1998),
.B(n_1937),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_2003),
.B(n_1964),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_2000),
.B(n_1945),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_2018),
.B(n_1987),
.Y(n_2041)
);

INVx2_ASAP7_75t_SL g2042 ( 
.A(n_2020),
.Y(n_2042)
);

INVx4_ASAP7_75t_L g2043 ( 
.A(n_1997),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_2015),
.B(n_1954),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_2010),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_2018),
.B(n_1939),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_2015),
.B(n_1962),
.Y(n_2047)
);

AND2x4_ASAP7_75t_SL g2048 ( 
.A(n_2024),
.B(n_1935),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_2022),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_2031),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_2031),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2049),
.Y(n_2052)
);

INVx3_ASAP7_75t_L g2053 ( 
.A(n_2035),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_2035),
.B(n_2013),
.Y(n_2054)
);

AO21x2_ASAP7_75t_L g2055 ( 
.A1(n_2028),
.A2(n_1994),
.B(n_2002),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_2031),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_2049),
.Y(n_2057)
);

OA21x2_ASAP7_75t_L g2058 ( 
.A1(n_2028),
.A2(n_1999),
.B(n_2001),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_2058),
.B(n_2030),
.Y(n_2059)
);

NAND2x1_ASAP7_75t_L g2060 ( 
.A(n_2054),
.B(n_2033),
.Y(n_2060)
);

HB1xp67_ASAP7_75t_L g2061 ( 
.A(n_2058),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_2054),
.B(n_2041),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_2053),
.B(n_2041),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_2058),
.B(n_2047),
.Y(n_2064)
);

AND2x2_ASAP7_75t_SL g2065 ( 
.A(n_2061),
.B(n_2058),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_2062),
.B(n_2063),
.Y(n_2066)
);

INVx1_ASAP7_75t_SL g2067 ( 
.A(n_2059),
.Y(n_2067)
);

HB1xp67_ASAP7_75t_L g2068 ( 
.A(n_2064),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2060),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2061),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2061),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_2062),
.B(n_2055),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_2062),
.B(n_2055),
.Y(n_2073)
);

AOI22xp33_ASAP7_75t_L g2074 ( 
.A1(n_2065),
.A2(n_2055),
.B1(n_1996),
.B2(n_1994),
.Y(n_2074)
);

A2O1A1Ixp33_ASAP7_75t_L g2075 ( 
.A1(n_2065),
.A2(n_2014),
.B(n_2037),
.C(n_2016),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2070),
.Y(n_2076)
);

AOI22xp5_ASAP7_75t_L g2077 ( 
.A1(n_2067),
.A2(n_2037),
.B1(n_2004),
.B2(n_2017),
.Y(n_2077)
);

OR2x2_ASAP7_75t_L g2078 ( 
.A(n_2068),
.B(n_2050),
.Y(n_2078)
);

HB1xp67_ASAP7_75t_L g2079 ( 
.A(n_2071),
.Y(n_2079)
);

INVx2_ASAP7_75t_SL g2080 ( 
.A(n_2066),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2066),
.Y(n_2081)
);

AOI22xp5_ASAP7_75t_L g2082 ( 
.A1(n_2072),
.A2(n_2027),
.B1(n_2026),
.B2(n_1990),
.Y(n_2082)
);

INVx2_ASAP7_75t_L g2083 ( 
.A(n_2072),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_2073),
.B(n_2052),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_2080),
.B(n_2073),
.Y(n_2085)
);

OR2x2_ASAP7_75t_L g2086 ( 
.A(n_2081),
.B(n_2069),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2079),
.Y(n_2087)
);

INVxp67_ASAP7_75t_SL g2088 ( 
.A(n_2074),
.Y(n_2088)
);

OR2x6_ASAP7_75t_L g2089 ( 
.A(n_2075),
.B(n_1995),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_2076),
.B(n_2069),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_2078),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_2083),
.B(n_2050),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2087),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2087),
.Y(n_2094)
);

NAND2x1p5_ASAP7_75t_L g2095 ( 
.A(n_2091),
.B(n_2043),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2086),
.Y(n_2096)
);

AND2x2_ASAP7_75t_SL g2097 ( 
.A(n_2096),
.B(n_2090),
.Y(n_2097)
);

INVxp67_ASAP7_75t_L g2098 ( 
.A(n_2093),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_2095),
.B(n_2085),
.Y(n_2099)
);

INVx1_ASAP7_75t_SL g2100 ( 
.A(n_2094),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_SL g2101 ( 
.A(n_2097),
.B(n_2077),
.Y(n_2101)
);

OAI211xp5_ASAP7_75t_L g2102 ( 
.A1(n_2100),
.A2(n_2088),
.B(n_2084),
.C(n_2082),
.Y(n_2102)
);

NAND3xp33_ASAP7_75t_L g2103 ( 
.A(n_2098),
.B(n_2089),
.C(n_2092),
.Y(n_2103)
);

NOR2xp33_ASAP7_75t_L g2104 ( 
.A(n_2099),
.B(n_2089),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2100),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2105),
.Y(n_2106)
);

A2O1A1Ixp33_ASAP7_75t_SL g2107 ( 
.A1(n_2104),
.A2(n_2102),
.B(n_2084),
.C(n_2101),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2103),
.Y(n_2108)
);

NAND4xp25_ASAP7_75t_SL g2109 ( 
.A(n_2102),
.B(n_2046),
.C(n_1993),
.D(n_1999),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2105),
.B(n_2050),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_2105),
.B(n_2051),
.Y(n_2111)
);

INVxp67_ASAP7_75t_L g2112 ( 
.A(n_2104),
.Y(n_2112)
);

NOR2xp33_ASAP7_75t_L g2113 ( 
.A(n_2104),
.B(n_2021),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_2105),
.B(n_2051),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_2105),
.B(n_2051),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2107),
.B(n_2029),
.Y(n_2116)
);

AOI221xp5_ASAP7_75t_L g2117 ( 
.A1(n_2109),
.A2(n_2023),
.B1(n_2057),
.B2(n_2052),
.C(n_2056),
.Y(n_2117)
);

NOR2xp33_ASAP7_75t_L g2118 ( 
.A(n_2112),
.B(n_1951),
.Y(n_2118)
);

OAI21xp5_ASAP7_75t_L g2119 ( 
.A1(n_2106),
.A2(n_2053),
.B(n_2046),
.Y(n_2119)
);

NAND3xp33_ASAP7_75t_L g2120 ( 
.A(n_2108),
.B(n_2043),
.C(n_2029),
.Y(n_2120)
);

AOI222xp33_ASAP7_75t_L g2121 ( 
.A1(n_2110),
.A2(n_2056),
.B1(n_1978),
.B2(n_2034),
.C1(n_2036),
.C2(n_2045),
.Y(n_2121)
);

AOI211xp5_ASAP7_75t_L g2122 ( 
.A1(n_2113),
.A2(n_2029),
.B(n_2033),
.C(n_1990),
.Y(n_2122)
);

NAND4xp25_ASAP7_75t_L g2123 ( 
.A(n_2111),
.B(n_2043),
.C(n_2053),
.D(n_1873),
.Y(n_2123)
);

AOI222xp33_ASAP7_75t_L g2124 ( 
.A1(n_2114),
.A2(n_2036),
.B1(n_2034),
.B2(n_2045),
.C1(n_2057),
.C2(n_1951),
.Y(n_2124)
);

AOI221x1_ASAP7_75t_L g2125 ( 
.A1(n_2115),
.A2(n_2043),
.B1(n_2053),
.B2(n_2025),
.C(n_2009),
.Y(n_2125)
);

O2A1O1Ixp33_ASAP7_75t_L g2126 ( 
.A1(n_2107),
.A2(n_2042),
.B(n_2040),
.C(n_1984),
.Y(n_2126)
);

BUFx12f_ASAP7_75t_L g2127 ( 
.A(n_2118),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_SL g2128 ( 
.A(n_2126),
.B(n_2116),
.Y(n_2128)
);

OR2x2_ASAP7_75t_L g2129 ( 
.A(n_2119),
.B(n_2042),
.Y(n_2129)
);

INVxp67_ASAP7_75t_L g2130 ( 
.A(n_2120),
.Y(n_2130)
);

BUFx2_ASAP7_75t_L g2131 ( 
.A(n_2123),
.Y(n_2131)
);

NOR2xp33_ASAP7_75t_L g2132 ( 
.A(n_2125),
.B(n_2038),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_2122),
.B(n_2040),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2117),
.Y(n_2134)
);

NAND2xp33_ASAP7_75t_L g2135 ( 
.A(n_2124),
.B(n_2038),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2121),
.B(n_2039),
.Y(n_2136)
);

NAND4xp75_ASAP7_75t_L g2137 ( 
.A(n_2128),
.B(n_1912),
.C(n_2039),
.D(n_2044),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2133),
.Y(n_2138)
);

NOR2xp67_ASAP7_75t_SL g2139 ( 
.A(n_2127),
.B(n_2020),
.Y(n_2139)
);

NOR2x1_ASAP7_75t_L g2140 ( 
.A(n_2134),
.B(n_2131),
.Y(n_2140)
);

NAND4xp75_ASAP7_75t_L g2141 ( 
.A(n_2132),
.B(n_1912),
.C(n_2044),
.D(n_1802),
.Y(n_2141)
);

NAND4xp75_ASAP7_75t_L g2142 ( 
.A(n_2136),
.B(n_1802),
.C(n_2032),
.D(n_2013),
.Y(n_2142)
);

NOR2xp33_ASAP7_75t_L g2143 ( 
.A(n_2129),
.B(n_1894),
.Y(n_2143)
);

OAI322xp33_ASAP7_75t_L g2144 ( 
.A1(n_2138),
.A2(n_2130),
.A3(n_2135),
.B1(n_1966),
.B2(n_2022),
.C1(n_2032),
.C2(n_1864),
.Y(n_2144)
);

OAI21xp33_ASAP7_75t_SL g2145 ( 
.A1(n_2142),
.A2(n_1947),
.B(n_1985),
.Y(n_2145)
);

NOR3xp33_ASAP7_75t_L g2146 ( 
.A(n_2140),
.B(n_2143),
.C(n_2137),
.Y(n_2146)
);

OR4x1_ASAP7_75t_L g2147 ( 
.A(n_2139),
.B(n_1991),
.C(n_2048),
.D(n_2035),
.Y(n_2147)
);

HB1xp67_ASAP7_75t_L g2148 ( 
.A(n_2141),
.Y(n_2148)
);

NOR3xp33_ASAP7_75t_L g2149 ( 
.A(n_2140),
.B(n_1940),
.C(n_1965),
.Y(n_2149)
);

HB1xp67_ASAP7_75t_L g2150 ( 
.A(n_2140),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2150),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2148),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2144),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2146),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2147),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_2151),
.B(n_2149),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2155),
.Y(n_2157)
);

NAND4xp75_ASAP7_75t_L g2158 ( 
.A(n_2152),
.B(n_2145),
.C(n_2006),
.D(n_2005),
.Y(n_2158)
);

OAI221xp5_ASAP7_75t_L g2159 ( 
.A1(n_2154),
.A2(n_1969),
.B1(n_2019),
.B2(n_1983),
.C(n_1980),
.Y(n_2159)
);

NAND3xp33_ASAP7_75t_SL g2160 ( 
.A(n_2156),
.B(n_2157),
.C(n_2153),
.Y(n_2160)
);

AOI21xp33_ASAP7_75t_L g2161 ( 
.A1(n_2158),
.A2(n_453),
.B(n_454),
.Y(n_2161)
);

NOR4xp25_ASAP7_75t_L g2162 ( 
.A(n_2159),
.B(n_2006),
.C(n_456),
.D(n_457),
.Y(n_2162)
);

OR5x1_ASAP7_75t_L g2163 ( 
.A(n_2157),
.B(n_2035),
.C(n_2048),
.D(n_2011),
.E(n_461),
.Y(n_2163)
);

NAND3xp33_ASAP7_75t_L g2164 ( 
.A(n_2157),
.B(n_1863),
.C(n_1833),
.Y(n_2164)
);

AOI221xp5_ASAP7_75t_L g2165 ( 
.A1(n_2160),
.A2(n_2048),
.B1(n_1946),
.B2(n_1948),
.C(n_1968),
.Y(n_2165)
);

OAI22xp5_ASAP7_75t_L g2166 ( 
.A1(n_2164),
.A2(n_1920),
.B1(n_1946),
.B2(n_1948),
.Y(n_2166)
);

OAI211xp5_ASAP7_75t_SL g2167 ( 
.A1(n_2161),
.A2(n_455),
.B(n_458),
.C(n_459),
.Y(n_2167)
);

AOI221xp5_ASAP7_75t_L g2168 ( 
.A1(n_2162),
.A2(n_1946),
.B1(n_1948),
.B2(n_1968),
.C(n_1988),
.Y(n_2168)
);

OAI21xp5_ASAP7_75t_L g2169 ( 
.A1(n_2167),
.A2(n_2163),
.B(n_1935),
.Y(n_2169)
);

AOI22xp5_ASAP7_75t_L g2170 ( 
.A1(n_2165),
.A2(n_1968),
.B1(n_1988),
.B2(n_2024),
.Y(n_2170)
);

INVxp67_ASAP7_75t_L g2171 ( 
.A(n_2168),
.Y(n_2171)
);

AOI22xp5_ASAP7_75t_L g2172 ( 
.A1(n_2171),
.A2(n_2166),
.B1(n_1988),
.B2(n_2024),
.Y(n_2172)
);

AOI21xp33_ASAP7_75t_L g2173 ( 
.A1(n_2169),
.A2(n_2170),
.B(n_464),
.Y(n_2173)
);

XNOR2xp5_ASAP7_75t_L g2174 ( 
.A(n_2171),
.B(n_462),
.Y(n_2174)
);

OR2x6_ASAP7_75t_L g2175 ( 
.A(n_2174),
.B(n_1838),
.Y(n_2175)
);

AOI22xp5_ASAP7_75t_L g2176 ( 
.A1(n_2172),
.A2(n_2173),
.B1(n_1833),
.B2(n_1863),
.Y(n_2176)
);

OR2x6_ASAP7_75t_L g2177 ( 
.A(n_2175),
.B(n_1863),
.Y(n_2177)
);

AO221x2_ASAP7_75t_SL g2178 ( 
.A1(n_2177),
.A2(n_2176),
.B1(n_467),
.B2(n_468),
.C(n_469),
.Y(n_2178)
);

OAI22xp5_ASAP7_75t_SL g2179 ( 
.A1(n_2178),
.A2(n_1879),
.B1(n_470),
.B2(n_471),
.Y(n_2179)
);

AOI211xp5_ASAP7_75t_L g2180 ( 
.A1(n_2179),
.A2(n_465),
.B(n_474),
.C(n_475),
.Y(n_2180)
);


endmodule