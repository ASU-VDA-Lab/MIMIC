module fake_netlist_5_1099_n_2016 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_2016);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_2016;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_326;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1406;
wire n_1279;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_783;
wire n_555;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1912;
wire n_1771;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1184;
wire n_1011;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1817;
wire n_1683;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g199 ( 
.A(n_86),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_147),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_46),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_41),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_41),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_100),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_8),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_154),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_158),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_38),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_57),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_11),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_153),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_181),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_115),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_172),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_43),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_119),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_139),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_167),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_91),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_174),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_59),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_39),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_79),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_103),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_166),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_117),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_31),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_113),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_173),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_58),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_64),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_192),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_99),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_145),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_58),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_159),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_89),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_24),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_143),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_62),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_15),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_157),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_34),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_163),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_175),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_3),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_125),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_136),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_168),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_26),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_11),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_161),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_111),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_83),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_170),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_142),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_82),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_6),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_69),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_150),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_24),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_185),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_182),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_48),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_189),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_164),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_9),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_48),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_13),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_171),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_169),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_47),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_92),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_70),
.Y(n_274)
);

INVxp67_ASAP7_75t_SL g275 ( 
.A(n_3),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_14),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_165),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_90),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_184),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_186),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_56),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_47),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_1),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_141),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_52),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_52),
.Y(n_286)
);

BUFx5_ASAP7_75t_L g287 ( 
.A(n_120),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_94),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_77),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_74),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_137),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_29),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_42),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_134),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_37),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_102),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_198),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_25),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_151),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_75),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_42),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_9),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_194),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_122),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_18),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_97),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_37),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_26),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_19),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_144),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_46),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_34),
.Y(n_312)
);

BUFx10_ASAP7_75t_L g313 ( 
.A(n_183),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_84),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_155),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_5),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_27),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_85),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_76),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_31),
.Y(n_320)
);

INVx4_ASAP7_75t_R g321 ( 
.A(n_160),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_188),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_39),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_45),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_118),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_44),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_98),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_114),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_128),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_20),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_10),
.Y(n_331)
);

BUFx10_ASAP7_75t_L g332 ( 
.A(n_55),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_5),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_131),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_180),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_53),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_43),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_60),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_44),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_4),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_30),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_21),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_135),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_53),
.Y(n_344)
);

BUFx10_ASAP7_75t_L g345 ( 
.A(n_66),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_73),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_126),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_110),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_176),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_45),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_55),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_80),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_132),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_71),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_21),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_17),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_93),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_178),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_127),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_33),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_121),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_146),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_133),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_62),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_105),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_4),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_67),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_19),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_104),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_162),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_107),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_96),
.Y(n_372)
);

BUFx10_ASAP7_75t_L g373 ( 
.A(n_30),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_18),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_108),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_61),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_138),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_65),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_156),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_8),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_40),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_179),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_72),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_1),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_63),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_197),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_40),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_64),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_123),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_140),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_38),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_0),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_15),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_60),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_2),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_191),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_212),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_220),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_378),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_271),
.B(n_0),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_245),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_223),
.Y(n_402)
);

NOR2xp67_ASAP7_75t_L g403 ( 
.A(n_309),
.B(n_2),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_240),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_367),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_240),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_240),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_247),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_249),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_252),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_240),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_253),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_257),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_274),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_240),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_260),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_288),
.B(n_6),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_309),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_323),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_263),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_211),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_236),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_211),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_265),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_323),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_248),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_256),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_270),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_381),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g430 ( 
.A(n_233),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_273),
.Y(n_431)
);

BUFx2_ASAP7_75t_SL g432 ( 
.A(n_271),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_289),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_381),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_246),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_246),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_317),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_290),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_317),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_338),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_R g441 ( 
.A(n_292),
.B(n_196),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_291),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_338),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_374),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_294),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_304),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_297),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_374),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_201),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_315),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_379),
.B(n_7),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_209),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_215),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_334),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_310),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_201),
.Y(n_456)
);

INVxp33_ASAP7_75t_SL g457 ( 
.A(n_202),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_222),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_314),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_202),
.Y(n_460)
);

NAND2xp33_ASAP7_75t_R g461 ( 
.A(n_200),
.B(n_7),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_227),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_238),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_318),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_322),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_327),
.Y(n_466)
);

INVxp67_ASAP7_75t_SL g467 ( 
.A(n_233),
.Y(n_467)
);

INVxp33_ASAP7_75t_L g468 ( 
.A(n_241),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_277),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_243),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_267),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_379),
.B(n_353),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_281),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_286),
.Y(n_474)
);

NOR2xp67_ASAP7_75t_L g475 ( 
.A(n_264),
.B(n_10),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_302),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_331),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_328),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_203),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_335),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_333),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_340),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_262),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_341),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_262),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_349),
.Y(n_486)
);

NOR2xp67_ASAP7_75t_L g487 ( 
.A(n_353),
.B(n_12),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_203),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_205),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_234),
.B(n_12),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_344),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_343),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_352),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_R g494 ( 
.A(n_346),
.B(n_195),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_356),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_386),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_279),
.B(n_13),
.Y(n_497)
);

INVxp67_ASAP7_75t_SL g498 ( 
.A(n_299),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_250),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_404),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_404),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_406),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_406),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_407),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_407),
.B(n_299),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_411),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_411),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_415),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_415),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_418),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_414),
.B(n_332),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_487),
.B(n_371),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_418),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_452),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_419),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_456),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_472),
.B(n_200),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_419),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_472),
.B(n_204),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_425),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_452),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_425),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_429),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_487),
.B(n_371),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_421),
.B(n_199),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_429),
.Y(n_526)
);

NAND2xp33_ASAP7_75t_L g527 ( 
.A(n_400),
.B(n_206),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_434),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_434),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_453),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_414),
.B(n_332),
.Y(n_531)
);

BUFx8_ASAP7_75t_L g532 ( 
.A(n_449),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_453),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_458),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_441),
.B(n_277),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_430),
.B(n_204),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_458),
.Y(n_537)
);

INVx5_ASAP7_75t_L g538 ( 
.A(n_423),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_467),
.B(n_213),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_423),
.Y(n_540)
);

AND3x2_ASAP7_75t_L g541 ( 
.A(n_417),
.B(n_275),
.C(n_364),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_462),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_462),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_423),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_463),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_463),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_496),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_470),
.Y(n_548)
);

INVx6_ASAP7_75t_L g549 ( 
.A(n_469),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_470),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_483),
.B(n_207),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_471),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_485),
.B(n_207),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_471),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_473),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_498),
.B(n_237),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_473),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_435),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_474),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_401),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_460),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_403),
.B(n_206),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_474),
.Y(n_563)
);

NAND2x1_ASAP7_75t_L g564 ( 
.A(n_400),
.B(n_321),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_476),
.Y(n_565)
);

BUFx8_ASAP7_75t_L g566 ( 
.A(n_449),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_476),
.Y(n_567)
);

INVx5_ASAP7_75t_L g568 ( 
.A(n_469),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_477),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_477),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_481),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_488),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_435),
.B(n_239),
.Y(n_573)
);

AND2x6_ASAP7_75t_L g574 ( 
.A(n_451),
.B(n_206),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_481),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_403),
.B(n_206),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_436),
.B(n_244),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_482),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_482),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_503),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_540),
.B(n_408),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_540),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_540),
.B(n_409),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_541),
.Y(n_584)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_538),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_568),
.B(n_410),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_574),
.A2(n_432),
.B1(n_399),
.B2(n_405),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_509),
.Y(n_588)
);

OAI22xp33_ASAP7_75t_SL g589 ( 
.A1(n_535),
.A2(n_457),
.B1(n_499),
.B2(n_497),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_574),
.A2(n_432),
.B1(n_489),
.B2(n_479),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_540),
.B(n_544),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_517),
.B(n_479),
.Y(n_592)
);

OAI22xp33_ASAP7_75t_L g593 ( 
.A1(n_511),
.A2(n_461),
.B1(n_295),
.B2(n_475),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_508),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_574),
.A2(n_489),
.B1(n_490),
.B2(n_475),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_509),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_561),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_503),
.Y(n_598)
);

NAND2xp33_ASAP7_75t_L g599 ( 
.A(n_574),
.B(n_494),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_568),
.B(n_412),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_509),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_509),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_500),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_500),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_508),
.Y(n_605)
);

NAND2x1p5_ASAP7_75t_L g606 ( 
.A(n_564),
.B(n_254),
.Y(n_606)
);

BUFx10_ASAP7_75t_L g607 ( 
.A(n_549),
.Y(n_607)
);

NAND2xp33_ASAP7_75t_L g608 ( 
.A(n_574),
.B(n_413),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_503),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_503),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_501),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_501),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_532),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_564),
.A2(n_420),
.B1(n_424),
.B2(n_416),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_502),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_568),
.B(n_428),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_502),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_532),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_538),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_504),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_504),
.Y(n_621)
);

INVx5_ASAP7_75t_L g622 ( 
.A(n_508),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_536),
.B(n_431),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_506),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_506),
.Y(n_625)
);

AND2x6_ASAP7_75t_L g626 ( 
.A(n_525),
.B(n_206),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_568),
.B(n_433),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_568),
.B(n_438),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_568),
.B(n_442),
.Y(n_629)
);

BUFx10_ASAP7_75t_L g630 ( 
.A(n_549),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_558),
.Y(n_631)
);

OR2x6_ASAP7_75t_L g632 ( 
.A(n_564),
.B(n_255),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_558),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_536),
.B(n_445),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_508),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_573),
.B(n_436),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_558),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_508),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_508),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_558),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_513),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_568),
.B(n_446),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_568),
.B(n_455),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_508),
.Y(n_644)
);

BUFx10_ASAP7_75t_L g645 ( 
.A(n_549),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_545),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_540),
.B(n_459),
.Y(n_647)
);

INVxp67_ASAP7_75t_SL g648 ( 
.A(n_544),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_579),
.Y(n_649)
);

INVx4_ASAP7_75t_SL g650 ( 
.A(n_574),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_579),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_551),
.B(n_464),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_513),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_544),
.B(n_465),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_579),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_568),
.B(n_466),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_508),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_579),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_579),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_513),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_545),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_511),
.A2(n_387),
.B1(n_324),
.B2(n_385),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_544),
.B(n_478),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_573),
.B(n_437),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_545),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_545),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_513),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_545),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_545),
.Y(n_669)
);

OR2x6_ASAP7_75t_L g670 ( 
.A(n_549),
.B(n_266),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_507),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_545),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_545),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_507),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_546),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_518),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_507),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_541),
.Y(n_678)
);

INVx6_ASAP7_75t_L g679 ( 
.A(n_538),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_518),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_547),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_507),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_544),
.B(n_480),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_546),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_546),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_517),
.B(n_437),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_551),
.B(n_486),
.Y(n_687)
);

NAND3xp33_ASAP7_75t_L g688 ( 
.A(n_519),
.B(n_493),
.C(n_440),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_546),
.Y(n_689)
);

INVx5_ASAP7_75t_L g690 ( 
.A(n_574),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_531),
.A2(n_342),
.B1(n_276),
.B2(n_376),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_518),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_518),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_553),
.B(n_468),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_535),
.B(n_277),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_522),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_574),
.A2(n_394),
.B1(n_366),
.B2(n_368),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_522),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_547),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_546),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_525),
.B(n_347),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_522),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_546),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_546),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_507),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_522),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_525),
.B(n_278),
.Y(n_707)
);

INVx4_ASAP7_75t_L g708 ( 
.A(n_538),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_523),
.Y(n_709)
);

NOR3xp33_ASAP7_75t_L g710 ( 
.A(n_516),
.B(n_384),
.C(n_380),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_531),
.A2(n_298),
.B1(n_235),
.B2(n_231),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_546),
.Y(n_712)
);

AND2x2_ASAP7_75t_SL g713 ( 
.A(n_527),
.B(n_232),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_552),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_523),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_552),
.Y(n_716)
);

AND2x4_ASAP7_75t_L g717 ( 
.A(n_505),
.B(n_280),
.Y(n_717)
);

BUFx2_ASAP7_75t_L g718 ( 
.A(n_532),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_505),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_539),
.B(n_284),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_552),
.Y(n_721)
);

INVx5_ASAP7_75t_L g722 ( 
.A(n_574),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_512),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_523),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_523),
.Y(n_725)
);

INVx5_ASAP7_75t_L g726 ( 
.A(n_574),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_561),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_526),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_516),
.A2(n_298),
.B1(n_235),
.B2(n_231),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_552),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_539),
.B(n_296),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_526),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_719),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_694),
.B(n_560),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_617),
.Y(n_735)
);

AO221x1_ASAP7_75t_L g736 ( 
.A1(n_593),
.A2(n_396),
.B1(n_232),
.B2(n_389),
.C(n_372),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_592),
.B(n_572),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_719),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_582),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_690),
.B(n_560),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_623),
.B(n_539),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_690),
.B(n_560),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_690),
.B(n_560),
.Y(n_743)
);

INVxp67_ASAP7_75t_SL g744 ( 
.A(n_582),
.Y(n_744)
);

OAI22xp33_ASAP7_75t_L g745 ( 
.A1(n_592),
.A2(n_686),
.B1(n_701),
.B2(n_711),
.Y(n_745)
);

NAND2xp33_ASAP7_75t_L g746 ( 
.A(n_626),
.B(n_574),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_634),
.B(n_560),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_636),
.B(n_572),
.Y(n_748)
);

INVxp33_ASAP7_75t_L g749 ( 
.A(n_727),
.Y(n_749)
);

O2A1O1Ixp33_ASAP7_75t_L g750 ( 
.A1(n_686),
.A2(n_527),
.B(n_519),
.C(n_556),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_588),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_652),
.B(n_556),
.Y(n_752)
);

INVx4_ASAP7_75t_L g753 ( 
.A(n_607),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_723),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_687),
.B(n_553),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_617),
.Y(n_756)
);

OAI22xp5_ASAP7_75t_L g757 ( 
.A1(n_595),
.A2(n_549),
.B1(n_397),
.B2(n_398),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_588),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_596),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_620),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_690),
.B(n_722),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_713),
.B(n_556),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_596),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_723),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_688),
.B(n_549),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_584),
.A2(n_402),
.B1(n_426),
.B2(n_427),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_636),
.B(n_573),
.Y(n_767)
);

NAND2xp33_ASAP7_75t_R g768 ( 
.A(n_613),
.B(n_422),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_601),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_601),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_591),
.A2(n_538),
.B(n_505),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_620),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_621),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_584),
.B(n_532),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_621),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_664),
.B(n_577),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_713),
.B(n_512),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_690),
.B(n_532),
.Y(n_778)
);

NOR3xp33_ASAP7_75t_SL g779 ( 
.A(n_695),
.B(n_208),
.C(n_205),
.Y(n_779)
);

HB1xp67_ASAP7_75t_L g780 ( 
.A(n_678),
.Y(n_780)
);

NAND3xp33_ASAP7_75t_L g781 ( 
.A(n_590),
.B(n_566),
.C(n_532),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_602),
.Y(n_782)
);

A2O1A1Ixp33_ASAP7_75t_L g783 ( 
.A1(n_707),
.A2(n_577),
.B(n_505),
.C(n_512),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_664),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_589),
.B(n_566),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_713),
.B(n_512),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_602),
.Y(n_787)
);

INVx8_ASAP7_75t_L g788 ( 
.A(n_670),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_717),
.B(n_577),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_678),
.A2(n_447),
.B1(n_454),
.B2(n_492),
.Y(n_790)
);

OAI22xp33_ASAP7_75t_L g791 ( 
.A1(n_711),
.A2(n_450),
.B1(n_375),
.B2(n_370),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_614),
.B(n_566),
.Y(n_792)
);

INVxp67_ASAP7_75t_L g793 ( 
.A(n_597),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_631),
.B(n_512),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_631),
.B(n_633),
.Y(n_795)
);

NOR2xp67_ASAP7_75t_L g796 ( 
.A(n_581),
.B(n_538),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_587),
.B(n_566),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_720),
.B(n_566),
.Y(n_798)
);

AND2x2_ASAP7_75t_SL g799 ( 
.A(n_613),
.B(n_232),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_633),
.B(n_512),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_599),
.A2(n_524),
.B1(n_505),
.B2(n_566),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_624),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_637),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_637),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_699),
.B(n_439),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_SL g806 ( 
.A(n_618),
.B(n_718),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_640),
.B(n_524),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_731),
.B(n_214),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_583),
.B(n_647),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_640),
.B(n_524),
.Y(n_810)
);

AOI221xp5_ASAP7_75t_L g811 ( 
.A1(n_729),
.A2(n_208),
.B1(n_210),
.B2(n_221),
.C(n_230),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_624),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_648),
.B(n_654),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_690),
.B(n_538),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_663),
.B(n_524),
.Y(n_815)
);

NOR2xp67_ASAP7_75t_L g816 ( 
.A(n_683),
.B(n_538),
.Y(n_816)
);

NOR2xp67_ASAP7_75t_L g817 ( 
.A(n_662),
.B(n_538),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_603),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_603),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_607),
.B(n_524),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_607),
.B(n_524),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_604),
.B(n_505),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_604),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_611),
.B(n_214),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_717),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_722),
.B(n_232),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_729),
.B(n_439),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_611),
.B(n_562),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_630),
.B(n_216),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_717),
.B(n_514),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_612),
.B(n_562),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_612),
.B(n_562),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_615),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_615),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_722),
.B(n_232),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_630),
.B(n_216),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_625),
.B(n_717),
.Y(n_837)
);

INVx1_ASAP7_75t_SL g838 ( 
.A(n_681),
.Y(n_838)
);

BUFx2_ASAP7_75t_L g839 ( 
.A(n_662),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_697),
.A2(n_393),
.B1(n_562),
.B2(n_576),
.Y(n_840)
);

NAND3xp33_ASAP7_75t_L g841 ( 
.A(n_710),
.B(n_691),
.C(n_608),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_625),
.B(n_562),
.Y(n_842)
);

BUFx6f_ASAP7_75t_SL g843 ( 
.A(n_632),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_691),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_630),
.B(n_217),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_722),
.B(n_372),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_649),
.B(n_217),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_649),
.B(n_562),
.Y(n_848)
);

A2O1A1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_651),
.A2(n_362),
.B(n_306),
.C(n_348),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_651),
.B(n_218),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_632),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_655),
.B(n_576),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_626),
.A2(n_576),
.B1(n_396),
.B2(n_389),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_655),
.B(n_576),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_670),
.B(n_514),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_658),
.B(n_218),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_L g857 ( 
.A1(n_670),
.A2(n_303),
.B1(n_319),
.B2(n_325),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_641),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_632),
.A2(n_576),
.B1(n_369),
.B2(n_377),
.Y(n_859)
);

NOR2x1p5_ASAP7_75t_L g860 ( 
.A(n_618),
.B(n_210),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_658),
.B(n_576),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_722),
.B(n_372),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_659),
.A2(n_329),
.B(n_520),
.C(n_578),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_722),
.B(n_372),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_718),
.B(n_440),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_645),
.B(n_219),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_670),
.B(n_443),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_659),
.B(n_552),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_645),
.B(n_219),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_670),
.A2(n_224),
.B1(n_377),
.B2(n_382),
.Y(n_870)
);

AND2x6_ASAP7_75t_L g871 ( 
.A(n_650),
.B(n_372),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_726),
.B(n_389),
.Y(n_872)
);

O2A1O1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_606),
.A2(n_578),
.B(n_537),
.C(n_570),
.Y(n_873)
);

BUFx6f_ASAP7_75t_SL g874 ( 
.A(n_632),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_632),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_626),
.A2(n_226),
.B1(n_225),
.B2(n_390),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_671),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_726),
.B(n_389),
.Y(n_878)
);

INVx1_ASAP7_75t_SL g879 ( 
.A(n_606),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_671),
.B(n_674),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_671),
.Y(n_881)
);

OR2x2_ASAP7_75t_L g882 ( 
.A(n_606),
.B(n_443),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_732),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_646),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_674),
.B(n_552),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_586),
.A2(n_300),
.B1(n_224),
.B2(n_225),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_674),
.B(n_552),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_650),
.B(n_521),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_677),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_677),
.B(n_552),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_732),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_641),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_677),
.B(n_571),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_682),
.B(n_571),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_682),
.B(n_705),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_653),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_645),
.B(n_226),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_653),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_726),
.B(n_389),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_682),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_705),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_705),
.B(n_571),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_SL g903 ( 
.A1(n_626),
.A2(n_313),
.B1(n_345),
.B2(n_332),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_626),
.B(n_571),
.Y(n_904)
);

O2A1O1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_762),
.A2(n_616),
.B(n_627),
.C(n_600),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_818),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_809),
.B(n_726),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_818),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_SL g909 ( 
.A(n_838),
.B(n_313),
.Y(n_909)
);

BUFx2_ASAP7_75t_SL g910 ( 
.A(n_748),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_888),
.Y(n_911)
);

INVxp67_ASAP7_75t_L g912 ( 
.A(n_805),
.Y(n_912)
);

NAND3xp33_ASAP7_75t_L g913 ( 
.A(n_755),
.B(n_258),
.C(n_251),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_737),
.B(n_444),
.Y(n_914)
);

INVx3_ASAP7_75t_L g915 ( 
.A(n_888),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_820),
.A2(n_726),
.B(n_629),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_821),
.A2(n_726),
.B(n_642),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_755),
.B(n_626),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_815),
.A2(n_643),
.B(n_628),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_738),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_819),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_813),
.A2(n_656),
.B(n_619),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_741),
.B(n_661),
.Y(n_923)
);

INVxp67_ASAP7_75t_L g924 ( 
.A(n_780),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_809),
.B(n_650),
.Y(n_925)
);

INVxp67_ASAP7_75t_L g926 ( 
.A(n_793),
.Y(n_926)
);

O2A1O1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_745),
.A2(n_752),
.B(n_750),
.C(n_784),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_819),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_808),
.B(n_626),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_823),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_776),
.B(n_444),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_794),
.A2(n_619),
.B(n_585),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_734),
.B(n_661),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_800),
.A2(n_619),
.B(n_585),
.Y(n_934)
);

NOR2x1_ASAP7_75t_L g935 ( 
.A(n_747),
.B(n_665),
.Y(n_935)
);

BUFx12f_ASAP7_75t_L g936 ( 
.A(n_844),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_777),
.A2(n_668),
.B(n_665),
.Y(n_937)
);

OAI21xp33_ASAP7_75t_L g938 ( 
.A1(n_811),
.A2(n_230),
.B(n_221),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_807),
.A2(n_708),
.B(n_585),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_791),
.B(n_668),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_810),
.A2(n_708),
.B(n_666),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_767),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_761),
.A2(n_783),
.B(n_786),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_837),
.A2(n_895),
.B(n_880),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_761),
.A2(n_708),
.B(n_666),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_754),
.B(n_650),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_754),
.B(n_721),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_841),
.A2(n_521),
.B(n_567),
.C(n_563),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_738),
.B(n_537),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_822),
.A2(n_672),
.B(n_669),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_848),
.A2(n_672),
.B(n_669),
.Y(n_951)
);

INVxp67_ASAP7_75t_L g952 ( 
.A(n_827),
.Y(n_952)
);

AO21x1_ASAP7_75t_L g953 ( 
.A1(n_797),
.A2(n_675),
.B(n_673),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_823),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_754),
.A2(n_666),
.B(n_646),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_767),
.Y(n_956)
);

INVx2_ASAP7_75t_SL g957 ( 
.A(n_865),
.Y(n_957)
);

AOI21x1_ASAP7_75t_L g958 ( 
.A1(n_828),
.A2(n_675),
.B(n_673),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_834),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_SL g960 ( 
.A(n_792),
.B(n_313),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_754),
.A2(n_666),
.B(n_646),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_764),
.A2(n_666),
.B(n_646),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_808),
.B(n_721),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_749),
.B(n_448),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_833),
.B(n_721),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_764),
.B(n_646),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_764),
.A2(n_730),
.B(n_685),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_764),
.A2(n_730),
.B(n_685),
.Y(n_968)
);

OAI21xp33_ASAP7_75t_L g969 ( 
.A1(n_824),
.A2(n_355),
.B(n_354),
.Y(n_969)
);

BUFx4f_ASAP7_75t_L g970 ( 
.A(n_855),
.Y(n_970)
);

OAI21xp33_ASAP7_75t_L g971 ( 
.A1(n_824),
.A2(n_355),
.B(n_354),
.Y(n_971)
);

NOR3xp33_ASAP7_75t_L g972 ( 
.A(n_757),
.B(n_839),
.C(n_785),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_831),
.A2(n_842),
.B(n_832),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_789),
.B(n_684),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_SL g975 ( 
.A(n_792),
.B(n_774),
.Y(n_975)
);

HB1xp67_ASAP7_75t_L g976 ( 
.A(n_789),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_852),
.A2(n_689),
.B(n_684),
.Y(n_977)
);

BUFx3_ASAP7_75t_L g978 ( 
.A(n_855),
.Y(n_978)
);

AOI22xp33_ASAP7_75t_L g979 ( 
.A1(n_736),
.A2(n_781),
.B1(n_799),
.B2(n_853),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_735),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_735),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_733),
.B(n_689),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_798),
.A2(n_703),
.B1(n_700),
.B2(n_704),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_774),
.B(n_700),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_733),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_798),
.A2(n_712),
.B1(n_703),
.B2(n_704),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_854),
.A2(n_861),
.B(n_795),
.Y(n_987)
);

O2A1O1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_751),
.A2(n_555),
.B(n_542),
.C(n_548),
.Y(n_988)
);

NOR2xp67_ASAP7_75t_L g989 ( 
.A(n_766),
.B(n_448),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_830),
.B(n_712),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_756),
.Y(n_991)
);

OAI21xp5_ASAP7_75t_L g992 ( 
.A1(n_885),
.A2(n_716),
.B(n_714),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_760),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_830),
.B(n_714),
.Y(n_994)
);

AOI21x1_ASAP7_75t_L g995 ( 
.A1(n_771),
.A2(n_716),
.B(n_598),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_847),
.B(n_594),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_884),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_879),
.B(n_594),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_847),
.B(n_594),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_739),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_739),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_753),
.A2(n_635),
.B(n_605),
.Y(n_1002)
);

AOI21xp33_ASAP7_75t_L g1003 ( 
.A1(n_882),
.A2(n_261),
.B(n_259),
.Y(n_1003)
);

AOI21x1_ASAP7_75t_L g1004 ( 
.A1(n_904),
.A2(n_598),
.B(n_580),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_765),
.A2(n_563),
.B(n_570),
.C(n_567),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_867),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_850),
.B(n_605),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_850),
.B(n_605),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_760),
.Y(n_1009)
);

BUFx4f_ASAP7_75t_L g1010 ( 
.A(n_788),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_753),
.A2(n_638),
.B(n_635),
.Y(n_1011)
);

OR2x2_ASAP7_75t_L g1012 ( 
.A(n_790),
.B(n_542),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_758),
.A2(n_559),
.B(n_557),
.C(n_555),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_856),
.B(n_635),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_744),
.A2(n_639),
.B(n_638),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_765),
.B(n_268),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_875),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_825),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_817),
.B(n_638),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_772),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_856),
.B(n_639),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_759),
.B(n_639),
.Y(n_1022)
);

NOR2x1_ASAP7_75t_L g1023 ( 
.A(n_860),
.B(n_644),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_887),
.A2(n_893),
.B(n_890),
.Y(n_1024)
);

NOR2xp67_ASAP7_75t_L g1025 ( 
.A(n_870),
.B(n_548),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_763),
.B(n_644),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_799),
.B(n_644),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_801),
.A2(n_228),
.B1(n_229),
.B2(n_242),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_772),
.Y(n_1029)
);

AOI21x1_ASAP7_75t_L g1030 ( 
.A1(n_868),
.A2(n_609),
.B(n_580),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_884),
.A2(n_657),
.B(n_622),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_884),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_769),
.B(n_657),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_884),
.A2(n_902),
.B(n_894),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_788),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_851),
.A2(n_877),
.B1(n_889),
.B2(n_881),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_770),
.B(n_269),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_746),
.A2(n_657),
.B(n_622),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_900),
.B(n_660),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_740),
.A2(n_622),
.B(n_660),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_773),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_779),
.B(n_903),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_773),
.Y(n_1043)
);

NAND3xp33_ASAP7_75t_L g1044 ( 
.A(n_886),
.B(n_282),
.C(n_272),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_806),
.B(n_550),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_775),
.Y(n_1046)
);

AOI21xp33_ASAP7_75t_L g1047 ( 
.A1(n_768),
.A2(n_285),
.B(n_283),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_853),
.A2(n_559),
.B(n_554),
.C(n_550),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_901),
.B(n_667),
.Y(n_1049)
);

INVx4_ASAP7_75t_L g1050 ( 
.A(n_788),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_740),
.A2(n_743),
.B(n_742),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_782),
.A2(n_728),
.B(n_725),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_742),
.A2(n_743),
.B(n_796),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_787),
.B(n_667),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_816),
.A2(n_622),
.B(n_725),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_803),
.B(n_554),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_804),
.B(n_676),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_859),
.A2(n_228),
.B1(n_229),
.B2(n_242),
.Y(n_1058)
);

OR2x2_ASAP7_75t_L g1059 ( 
.A(n_802),
.B(n_557),
.Y(n_1059)
);

INVxp67_ASAP7_75t_L g1060 ( 
.A(n_768),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_802),
.B(n_345),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_812),
.B(n_676),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_858),
.B(n_883),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_858),
.B(n_680),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_873),
.B(n_680),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_840),
.A2(n_520),
.B(n_495),
.C(n_491),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_883),
.B(n_692),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_891),
.B(n_692),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_814),
.A2(n_622),
.B(n_724),
.Y(n_1069)
);

INVx4_ASAP7_75t_L g1070 ( 
.A(n_843),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_891),
.B(n_693),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_892),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_829),
.B(n_293),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_840),
.B(n_345),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_814),
.A2(n_622),
.B(n_724),
.Y(n_1075)
);

AO21x1_ASAP7_75t_L g1076 ( 
.A1(n_778),
.A2(n_728),
.B(n_715),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_892),
.B(n_693),
.Y(n_1077)
);

AOI21xp33_ASAP7_75t_L g1078 ( 
.A1(n_836),
.A2(n_308),
.B(n_301),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_863),
.A2(n_715),
.B(n_709),
.C(n_706),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_778),
.A2(n_383),
.B1(n_357),
.B2(n_358),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_826),
.A2(n_709),
.B(n_706),
.Y(n_1081)
);

A2O1A1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_896),
.A2(n_898),
.B(n_876),
.C(n_849),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_898),
.B(n_696),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_826),
.A2(n_702),
.B(n_698),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_899),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_871),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_899),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_R g1088 ( 
.A(n_843),
.B(n_300),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_897),
.B(n_305),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_835),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_845),
.B(n_307),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_835),
.A2(n_702),
.B(n_698),
.Y(n_1092)
);

AOI21x1_ASAP7_75t_L g1093 ( 
.A1(n_846),
.A2(n_610),
.B(n_609),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_979),
.A2(n_874),
.B1(n_857),
.B2(n_360),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_911),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_979),
.A2(n_874),
.B1(n_360),
.B2(n_388),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_911),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_923),
.B(n_696),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_1016),
.A2(n_869),
.B(n_866),
.C(n_878),
.Y(n_1099)
);

AO22x1_ASAP7_75t_L g1100 ( 
.A1(n_1074),
.A2(n_388),
.B1(n_391),
.B2(n_392),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1016),
.B(n_530),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_975),
.A2(n_361),
.B1(n_363),
.B2(n_365),
.Y(n_1102)
);

O2A1O1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_960),
.A2(n_878),
.B(n_872),
.C(n_864),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_978),
.B(n_484),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_978),
.B(n_484),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_970),
.B(n_357),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_SL g1107 ( 
.A1(n_910),
.A2(n_373),
.B1(n_392),
.B2(n_391),
.Y(n_1107)
);

CKINVDCx8_ASAP7_75t_R g1108 ( 
.A(n_1035),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_923),
.B(n_520),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_908),
.B(n_520),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_927),
.B(n_520),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_952),
.B(n_610),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_906),
.Y(n_1113)
);

AOI21x1_ASAP7_75t_L g1114 ( 
.A1(n_907),
.A2(n_872),
.B(n_864),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_972),
.A2(n_846),
.B(n_862),
.C(n_383),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_921),
.Y(n_1116)
);

INVxp67_ASAP7_75t_L g1117 ( 
.A(n_964),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_919),
.A2(n_862),
.B(n_871),
.Y(n_1118)
);

INVx4_ASAP7_75t_L g1119 ( 
.A(n_1035),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_912),
.B(n_373),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_915),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_SL g1122 ( 
.A1(n_936),
.A2(n_1060),
.B1(n_1089),
.B2(n_1073),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_943),
.A2(n_973),
.B(n_1005),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_970),
.B(n_358),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_1006),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_940),
.A2(n_382),
.B(n_359),
.C(n_361),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_987),
.A2(n_871),
.B(n_679),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_931),
.B(n_871),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_928),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_957),
.B(n_914),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_1006),
.A2(n_871),
.B1(n_287),
.B2(n_396),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1051),
.A2(n_922),
.B(n_1019),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1061),
.B(n_373),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_SL g1134 ( 
.A(n_1070),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1019),
.A2(n_679),
.B(n_575),
.Y(n_1135)
);

NAND2xp33_ASAP7_75t_SL g1136 ( 
.A(n_1035),
.B(n_1050),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_944),
.A2(n_679),
.B(n_575),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_942),
.B(n_491),
.Y(n_1138)
);

INVxp67_ASAP7_75t_L g1139 ( 
.A(n_926),
.Y(n_1139)
);

AOI21xp33_ASAP7_75t_L g1140 ( 
.A1(n_940),
.A2(n_495),
.B(n_395),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1041),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_991),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_920),
.B(n_359),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_1035),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_R g1145 ( 
.A(n_1010),
.B(n_363),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_920),
.B(n_365),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_924),
.B(n_311),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_930),
.B(n_571),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1053),
.A2(n_679),
.B(n_575),
.Y(n_1149)
);

CKINVDCx6p67_ASAP7_75t_R g1150 ( 
.A(n_1070),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_942),
.B(n_312),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_954),
.B(n_571),
.Y(n_1152)
);

O2A1O1Ixp5_ASAP7_75t_L g1153 ( 
.A1(n_983),
.A2(n_953),
.B(n_1076),
.C(n_929),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_959),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_956),
.B(n_316),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_950),
.A2(n_575),
.B(n_530),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1059),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_980),
.Y(n_1158)
);

BUFx12f_ASAP7_75t_L g1159 ( 
.A(n_920),
.Y(n_1159)
);

O2A1O1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_1003),
.A2(n_569),
.B(n_565),
.C(n_543),
.Y(n_1160)
);

A2O1A1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_1073),
.A2(n_369),
.B(n_390),
.C(n_336),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_1050),
.B(n_530),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_948),
.B(n_918),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_905),
.A2(n_530),
.B(n_569),
.Y(n_1164)
);

A2O1A1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1089),
.A2(n_320),
.B(n_337),
.C(n_339),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_907),
.A2(n_569),
.B(n_565),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_991),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_993),
.Y(n_1168)
);

AO22x1_ASAP7_75t_L g1169 ( 
.A1(n_1091),
.A2(n_395),
.B1(n_330),
.B2(n_350),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_948),
.A2(n_533),
.B(n_565),
.C(n_543),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1029),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_920),
.B(n_571),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1017),
.B(n_533),
.Y(n_1173)
);

OAI22x1_ASAP7_75t_L g1174 ( 
.A1(n_1042),
.A2(n_326),
.B1(n_351),
.B2(n_17),
.Y(n_1174)
);

NOR2xp67_ASAP7_75t_L g1175 ( 
.A(n_913),
.B(n_87),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_993),
.B(n_1043),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_976),
.B(n_571),
.Y(n_1177)
);

NOR3xp33_ASAP7_75t_SL g1178 ( 
.A(n_938),
.B(n_14),
.C(n_16),
.Y(n_1178)
);

BUFx2_ASAP7_75t_SL g1179 ( 
.A(n_1017),
.Y(n_1179)
);

BUFx8_ASAP7_75t_L g1180 ( 
.A(n_1045),
.Y(n_1180)
);

NOR2xp67_ASAP7_75t_SL g1181 ( 
.A(n_1086),
.B(n_396),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_992),
.A2(n_569),
.B(n_565),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_951),
.A2(n_543),
.B(n_534),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_963),
.A2(n_543),
.B(n_534),
.Y(n_1184)
);

O2A1O1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1047),
.A2(n_534),
.B(n_533),
.C(n_529),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_996),
.A2(n_534),
.B(n_533),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_997),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_956),
.B(n_16),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_976),
.B(n_528),
.Y(n_1189)
);

BUFx8_ASAP7_75t_SL g1190 ( 
.A(n_1010),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1043),
.B(n_529),
.Y(n_1191)
);

NOR3xp33_ASAP7_75t_L g1192 ( 
.A(n_1091),
.B(n_529),
.C(n_528),
.Y(n_1192)
);

INVxp67_ASAP7_75t_SL g1193 ( 
.A(n_997),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_949),
.B(n_529),
.Y(n_1194)
);

NAND2x1p5_ASAP7_75t_L g1195 ( 
.A(n_915),
.B(n_396),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_1012),
.B(n_528),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_969),
.B(n_20),
.Y(n_1197)
);

O2A1O1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_971),
.A2(n_528),
.B(n_526),
.C(n_25),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1046),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_999),
.A2(n_526),
.B(n_515),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1037),
.B(n_22),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_949),
.B(n_515),
.Y(n_1202)
);

BUFx4f_ASAP7_75t_L g1203 ( 
.A(n_1086),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1007),
.A2(n_510),
.B(n_515),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_997),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_997),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1008),
.A2(n_1021),
.B(n_1014),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1046),
.B(n_515),
.Y(n_1208)
);

BUFx3_ASAP7_75t_L g1209 ( 
.A(n_1056),
.Y(n_1209)
);

AOI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1037),
.A2(n_287),
.B1(n_515),
.B2(n_510),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1025),
.A2(n_515),
.B(n_510),
.C(n_287),
.Y(n_1211)
);

AOI222xp33_ASAP7_75t_L g1212 ( 
.A1(n_1058),
.A2(n_515),
.B1(n_510),
.B2(n_27),
.C1(n_28),
.C2(n_29),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1048),
.A2(n_510),
.B1(n_515),
.B2(n_28),
.Y(n_1213)
);

O2A1O1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1005),
.A2(n_1078),
.B(n_1080),
.C(n_1028),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_SL g1215 ( 
.A1(n_984),
.A2(n_287),
.B(n_129),
.C(n_193),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1056),
.B(n_510),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_981),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1023),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_1088),
.Y(n_1219)
);

NAND3xp33_ASAP7_75t_SL g1220 ( 
.A(n_909),
.B(n_1088),
.C(n_1044),
.Y(n_1220)
);

A2O1A1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_937),
.A2(n_510),
.B(n_287),
.C(n_32),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_916),
.A2(n_510),
.B(n_124),
.Y(n_1222)
);

NOR3xp33_ASAP7_75t_L g1223 ( 
.A(n_989),
.B(n_287),
.C(n_23),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1048),
.A2(n_22),
.B1(n_23),
.B2(n_32),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1072),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1018),
.B(n_287),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1032),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_984),
.A2(n_287),
.B(n_35),
.C(n_36),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_1032),
.Y(n_1229)
);

INVx2_ASAP7_75t_SL g1230 ( 
.A(n_974),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_917),
.A2(n_190),
.B(n_187),
.Y(n_1231)
);

NAND3xp33_ASAP7_75t_SL g1232 ( 
.A(n_988),
.B(n_33),
.C(n_35),
.Y(n_1232)
);

OR2x6_ASAP7_75t_SL g1233 ( 
.A(n_1036),
.B(n_36),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_985),
.B(n_177),
.Y(n_1234)
);

NAND2x1p5_ASAP7_75t_L g1235 ( 
.A(n_1032),
.B(n_152),
.Y(n_1235)
);

INVxp67_ASAP7_75t_L g1236 ( 
.A(n_990),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1009),
.Y(n_1237)
);

AOI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_994),
.A2(n_149),
.B1(n_148),
.B2(n_130),
.Y(n_1238)
);

NOR3xp33_ASAP7_75t_SL g1239 ( 
.A(n_1013),
.B(n_49),
.C(n_50),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1020),
.B(n_49),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_985),
.Y(n_1241)
);

OAI21xp33_ASAP7_75t_SL g1242 ( 
.A1(n_1027),
.A2(n_925),
.B(n_986),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1066),
.A2(n_1027),
.B1(n_1000),
.B2(n_1001),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1000),
.B(n_1001),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1063),
.Y(n_1245)
);

O2A1O1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1082),
.A2(n_50),
.B(n_51),
.C(n_54),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_925),
.B(n_51),
.Y(n_1247)
);

NAND2x1p5_ASAP7_75t_L g1248 ( 
.A(n_1032),
.B(n_116),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1034),
.A2(n_112),
.B(n_109),
.Y(n_1249)
);

AOI221xp5_ASAP7_75t_L g1250 ( 
.A1(n_1066),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.C(n_59),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1087),
.Y(n_1251)
);

OR2x2_ASAP7_75t_L g1252 ( 
.A(n_1117),
.B(n_1085),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1139),
.Y(n_1253)
);

INVx3_ASAP7_75t_L g1254 ( 
.A(n_1108),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1207),
.A2(n_933),
.B(n_1024),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1167),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1236),
.B(n_998),
.Y(n_1257)
);

OAI22x1_ASAP7_75t_L g1258 ( 
.A1(n_1201),
.A2(n_998),
.B1(n_933),
.B2(n_1090),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1132),
.A2(n_1065),
.B(n_941),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1164),
.A2(n_1030),
.B(n_1004),
.Y(n_1260)
);

OA21x2_ASAP7_75t_L g1261 ( 
.A1(n_1123),
.A2(n_1065),
.B(n_1052),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1166),
.A2(n_995),
.B(n_1093),
.Y(n_1262)
);

AO31x2_ASAP7_75t_L g1263 ( 
.A1(n_1221),
.A2(n_1082),
.A3(n_977),
.B(n_967),
.Y(n_1263)
);

A2O1A1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1214),
.A2(n_935),
.B(n_1079),
.C(n_968),
.Y(n_1264)
);

INVx3_ASAP7_75t_L g1265 ( 
.A(n_1144),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_1159),
.Y(n_1266)
);

NAND3x1_ASAP7_75t_L g1267 ( 
.A(n_1197),
.B(n_965),
.C(n_63),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1123),
.A2(n_966),
.B(n_955),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1133),
.B(n_1039),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1101),
.A2(n_966),
.B(n_962),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1163),
.A2(n_961),
.B(n_982),
.Y(n_1271)
);

AO32x2_ASAP7_75t_L g1272 ( 
.A1(n_1224),
.A2(n_958),
.A3(n_1067),
.B1(n_1068),
.B2(n_1071),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1158),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1184),
.A2(n_1092),
.B(n_1084),
.Y(n_1274)
);

BUFx2_ASAP7_75t_SL g1275 ( 
.A(n_1134),
.Y(n_1275)
);

BUFx2_ASAP7_75t_R g1276 ( 
.A(n_1190),
.Y(n_1276)
);

AOI221x1_ASAP7_75t_L g1277 ( 
.A1(n_1140),
.A2(n_1015),
.B1(n_1040),
.B2(n_1055),
.C(n_1011),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1186),
.A2(n_1081),
.B(n_1002),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_1130),
.B(n_1086),
.Y(n_1279)
);

AO31x2_ASAP7_75t_L g1280 ( 
.A1(n_1111),
.A2(n_1033),
.A3(n_1026),
.B(n_1022),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1204),
.A2(n_1038),
.B(n_1039),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1163),
.A2(n_1127),
.B(n_1118),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1157),
.B(n_1057),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1098),
.A2(n_939),
.B(n_934),
.Y(n_1284)
);

INVx3_ASAP7_75t_SL g1285 ( 
.A(n_1150),
.Y(n_1285)
);

BUFx10_ASAP7_75t_L g1286 ( 
.A(n_1134),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1230),
.B(n_1054),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1138),
.B(n_1049),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1122),
.A2(n_947),
.B1(n_946),
.B2(n_1049),
.Y(n_1289)
);

AOI221x1_ASAP7_75t_L g1290 ( 
.A1(n_1140),
.A2(n_1062),
.B1(n_1075),
.B2(n_1069),
.C(n_1083),
.Y(n_1290)
);

OAI22x1_ASAP7_75t_L g1291 ( 
.A1(n_1247),
.A2(n_1188),
.B1(n_1251),
.B2(n_1102),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1171),
.Y(n_1292)
);

AOI21xp33_ASAP7_75t_SL g1293 ( 
.A1(n_1174),
.A2(n_61),
.B(n_65),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1098),
.A2(n_932),
.B(n_947),
.Y(n_1294)
);

AOI221x1_ASAP7_75t_L g1295 ( 
.A1(n_1228),
.A2(n_1064),
.B1(n_1031),
.B2(n_945),
.C(n_1086),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1180),
.Y(n_1296)
);

BUFx2_ASAP7_75t_L g1297 ( 
.A(n_1180),
.Y(n_1297)
);

A2O1A1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1099),
.A2(n_946),
.B(n_1071),
.C(n_1068),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1125),
.B(n_1077),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1200),
.A2(n_1077),
.B(n_1067),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1168),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_L g1302 ( 
.A(n_1209),
.Y(n_1302)
);

AO221x2_ASAP7_75t_L g1303 ( 
.A1(n_1224),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.C(n_69),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1149),
.A2(n_81),
.B(n_101),
.Y(n_1304)
);

AO31x2_ASAP7_75t_L g1305 ( 
.A1(n_1111),
.A2(n_68),
.A3(n_70),
.B(n_71),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1196),
.A2(n_78),
.B1(n_88),
.B2(n_95),
.Y(n_1306)
);

BUFx10_ASAP7_75t_L g1307 ( 
.A(n_1151),
.Y(n_1307)
);

AND2x4_ASAP7_75t_L g1308 ( 
.A(n_1173),
.B(n_106),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1245),
.B(n_1244),
.Y(n_1309)
);

AOI221xp5_ASAP7_75t_L g1310 ( 
.A1(n_1169),
.A2(n_1100),
.B1(n_1096),
.B2(n_1165),
.C(n_1220),
.Y(n_1310)
);

NAND2x1_ASAP7_75t_L g1311 ( 
.A(n_1119),
.B(n_1095),
.Y(n_1311)
);

AOI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1156),
.A2(n_1183),
.B(n_1182),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1109),
.A2(n_1137),
.B(n_1242),
.Y(n_1313)
);

OAI22x1_ASAP7_75t_L g1314 ( 
.A1(n_1212),
.A2(n_1218),
.B1(n_1233),
.B2(n_1146),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_1173),
.B(n_1104),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1213),
.A2(n_1178),
.B1(n_1113),
.B2(n_1116),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1109),
.A2(n_1153),
.B(n_1243),
.Y(n_1317)
);

OAI21xp33_ASAP7_75t_L g1318 ( 
.A1(n_1155),
.A2(n_1212),
.B(n_1147),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1199),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1243),
.A2(n_1249),
.B(n_1103),
.Y(n_1320)
);

AO21x1_ASAP7_75t_L g1321 ( 
.A1(n_1213),
.A2(n_1246),
.B(n_1198),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1128),
.A2(n_1222),
.B(n_1176),
.Y(n_1322)
);

OR2x2_ASAP7_75t_L g1323 ( 
.A(n_1112),
.B(n_1120),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1211),
.A2(n_1160),
.B(n_1170),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1128),
.A2(n_1216),
.B(n_1191),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1217),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_SL g1327 ( 
.A1(n_1107),
.A2(n_1096),
.B1(n_1094),
.B2(n_1219),
.Y(n_1327)
);

NOR4xp25_ASAP7_75t_L g1328 ( 
.A(n_1232),
.B(n_1250),
.C(n_1126),
.D(n_1094),
.Y(n_1328)
);

AO21x2_ASAP7_75t_L g1329 ( 
.A1(n_1215),
.A2(n_1192),
.B(n_1210),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1237),
.Y(n_1330)
);

A2O1A1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1161),
.A2(n_1175),
.B(n_1115),
.C(n_1223),
.Y(n_1331)
);

INVxp67_ASAP7_75t_SL g1332 ( 
.A(n_1187),
.Y(n_1332)
);

NAND2x1p5_ASAP7_75t_L g1333 ( 
.A(n_1119),
.B(n_1144),
.Y(n_1333)
);

A2O1A1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1239),
.A2(n_1112),
.B(n_1238),
.C(n_1231),
.Y(n_1334)
);

CKINVDCx11_ASAP7_75t_R g1335 ( 
.A(n_1144),
.Y(n_1335)
);

BUFx8_ASAP7_75t_L g1336 ( 
.A(n_1229),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1191),
.A2(n_1148),
.B(n_1152),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1114),
.A2(n_1208),
.B(n_1152),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1194),
.B(n_1105),
.Y(n_1339)
);

OA21x2_ASAP7_75t_L g1340 ( 
.A1(n_1148),
.A2(n_1208),
.B(n_1110),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1129),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1154),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_1104),
.Y(n_1343)
);

AOI211x1_ASAP7_75t_L g1344 ( 
.A1(n_1240),
.A2(n_1143),
.B(n_1106),
.C(n_1124),
.Y(n_1344)
);

NOR2xp67_ASAP7_75t_L g1345 ( 
.A(n_1241),
.B(n_1105),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1135),
.A2(n_1177),
.B(n_1172),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1225),
.Y(n_1347)
);

AOI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1234),
.A2(n_1179),
.B1(n_1189),
.B2(n_1202),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1189),
.Y(n_1349)
);

AOI221x1_ASAP7_75t_L g1350 ( 
.A1(n_1226),
.A2(n_1136),
.B1(n_1110),
.B2(n_1234),
.C(n_1205),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_1145),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_SL g1352 ( 
.A(n_1095),
.B(n_1097),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1162),
.B(n_1097),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1195),
.A2(n_1185),
.B(n_1235),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1131),
.A2(n_1141),
.B(n_1195),
.Y(n_1355)
);

CKINVDCx11_ASAP7_75t_R g1356 ( 
.A(n_1187),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1121),
.B(n_1162),
.Y(n_1357)
);

INVx2_ASAP7_75t_SL g1358 ( 
.A(n_1203),
.Y(n_1358)
);

OAI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1248),
.A2(n_1121),
.B(n_1193),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_SL g1360 ( 
.A1(n_1203),
.A2(n_1181),
.B(n_1187),
.Y(n_1360)
);

A2O1A1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1206),
.A2(n_755),
.B(n_1201),
.C(n_1214),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1206),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1206),
.Y(n_1363)
);

A2O1A1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1227),
.A2(n_755),
.B(n_1201),
.C(n_1214),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1227),
.B(n_755),
.Y(n_1365)
);

AOI211xp5_ASAP7_75t_L g1366 ( 
.A1(n_1140),
.A2(n_1201),
.B(n_791),
.C(n_745),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1245),
.B(n_755),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1125),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1207),
.A2(n_821),
.B(n_820),
.Y(n_1369)
);

BUFx6f_ASAP7_75t_L g1370 ( 
.A(n_1159),
.Y(n_1370)
);

INVx1_ASAP7_75t_SL g1371 ( 
.A(n_1125),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1245),
.B(n_755),
.Y(n_1372)
);

OAI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1153),
.A2(n_1163),
.B(n_1123),
.Y(n_1373)
);

NOR2xp67_ASAP7_75t_SL g1374 ( 
.A(n_1108),
.B(n_613),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_SL g1375 ( 
.A1(n_1099),
.A2(n_753),
.B(n_778),
.Y(n_1375)
);

AO32x2_ASAP7_75t_L g1376 ( 
.A1(n_1224),
.A2(n_1213),
.A3(n_1094),
.B1(n_1243),
.B2(n_1096),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1132),
.A2(n_1030),
.B(n_1164),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1245),
.B(n_755),
.Y(n_1378)
);

O2A1O1Ixp33_ASAP7_75t_L g1379 ( 
.A1(n_1201),
.A2(n_1140),
.B(n_755),
.C(n_960),
.Y(n_1379)
);

OAI221xp5_ASAP7_75t_L g1380 ( 
.A1(n_1201),
.A2(n_691),
.B1(n_662),
.B2(n_511),
.C(n_531),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1207),
.A2(n_821),
.B(n_820),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1219),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_1180),
.Y(n_1383)
);

AO21x2_ASAP7_75t_L g1384 ( 
.A1(n_1123),
.A2(n_1207),
.B(n_1132),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1133),
.B(n_910),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1117),
.B(n_838),
.Y(n_1386)
);

BUFx2_ASAP7_75t_SL g1387 ( 
.A(n_1108),
.Y(n_1387)
);

O2A1O1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1201),
.A2(n_1140),
.B(n_755),
.C(n_960),
.Y(n_1388)
);

AOI221x1_ASAP7_75t_L g1389 ( 
.A1(n_1201),
.A2(n_1140),
.B1(n_972),
.B2(n_1228),
.C(n_1224),
.Y(n_1389)
);

NAND2xp33_ASAP7_75t_R g1390 ( 
.A(n_1219),
.B(n_547),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1245),
.B(n_755),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1158),
.Y(n_1392)
);

BUFx10_ASAP7_75t_L g1393 ( 
.A(n_1134),
.Y(n_1393)
);

AOI221x1_ASAP7_75t_L g1394 ( 
.A1(n_1201),
.A2(n_1140),
.B1(n_972),
.B2(n_1228),
.C(n_1224),
.Y(n_1394)
);

OA21x2_ASAP7_75t_L g1395 ( 
.A1(n_1123),
.A2(n_1153),
.B(n_1207),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1158),
.Y(n_1396)
);

O2A1O1Ixp33_ASAP7_75t_SL g1397 ( 
.A1(n_1099),
.A2(n_1221),
.B(n_1228),
.C(n_797),
.Y(n_1397)
);

OAI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1153),
.A2(n_1163),
.B(n_1123),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1132),
.A2(n_1030),
.B(n_1164),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1142),
.Y(n_1400)
);

OAI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1153),
.A2(n_1163),
.B(n_1123),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1139),
.B(n_496),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1153),
.A2(n_1163),
.B(n_1123),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1245),
.B(n_755),
.Y(n_1404)
);

BUFx10_ASAP7_75t_L g1405 ( 
.A(n_1134),
.Y(n_1405)
);

AO32x2_ASAP7_75t_L g1406 ( 
.A1(n_1224),
.A2(n_1213),
.A3(n_1094),
.B1(n_1243),
.B2(n_1096),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1207),
.A2(n_821),
.B(n_820),
.Y(n_1407)
);

BUFx6f_ASAP7_75t_L g1408 ( 
.A(n_1159),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1207),
.A2(n_821),
.B(n_820),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1245),
.B(n_755),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1133),
.B(n_910),
.Y(n_1411)
);

INVx3_ASAP7_75t_SL g1412 ( 
.A(n_1382),
.Y(n_1412)
);

INVx6_ASAP7_75t_L g1413 ( 
.A(n_1336),
.Y(n_1413)
);

BUFx8_ASAP7_75t_L g1414 ( 
.A(n_1266),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1366),
.A2(n_1318),
.B1(n_1380),
.B2(n_1388),
.Y(n_1415)
);

INVx6_ASAP7_75t_L g1416 ( 
.A(n_1336),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1303),
.A2(n_1327),
.B1(n_1310),
.B2(n_1321),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_SL g1418 ( 
.A1(n_1303),
.A2(n_1327),
.B1(n_1398),
.B2(n_1401),
.Y(n_1418)
);

BUFx8_ASAP7_75t_SL g1419 ( 
.A(n_1297),
.Y(n_1419)
);

BUFx4f_ASAP7_75t_SL g1420 ( 
.A(n_1266),
.Y(n_1420)
);

INVx4_ASAP7_75t_L g1421 ( 
.A(n_1266),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_SL g1422 ( 
.A1(n_1373),
.A2(n_1401),
.B1(n_1403),
.B2(n_1398),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1370),
.Y(n_1423)
);

BUFx2_ASAP7_75t_SL g1424 ( 
.A(n_1370),
.Y(n_1424)
);

CKINVDCx11_ASAP7_75t_R g1425 ( 
.A(n_1286),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1314),
.A2(n_1291),
.B1(n_1403),
.B2(n_1373),
.Y(n_1426)
);

CKINVDCx6p67_ASAP7_75t_R g1427 ( 
.A(n_1285),
.Y(n_1427)
);

INVx6_ASAP7_75t_L g1428 ( 
.A(n_1408),
.Y(n_1428)
);

AO22x1_ASAP7_75t_L g1429 ( 
.A1(n_1385),
.A2(n_1411),
.B1(n_1351),
.B2(n_1402),
.Y(n_1429)
);

INVx4_ASAP7_75t_L g1430 ( 
.A(n_1408),
.Y(n_1430)
);

BUFx6f_ASAP7_75t_L g1431 ( 
.A(n_1356),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1367),
.A2(n_1410),
.B1(n_1378),
.B2(n_1404),
.Y(n_1432)
);

INVx4_ASAP7_75t_L g1433 ( 
.A(n_1408),
.Y(n_1433)
);

AOI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1366),
.A2(n_1390),
.B1(n_1269),
.B2(n_1307),
.Y(n_1434)
);

INVx2_ASAP7_75t_SL g1435 ( 
.A(n_1286),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1256),
.Y(n_1436)
);

BUFx10_ASAP7_75t_L g1437 ( 
.A(n_1296),
.Y(n_1437)
);

CKINVDCx11_ASAP7_75t_R g1438 ( 
.A(n_1393),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1367),
.A2(n_1410),
.B1(n_1404),
.B2(n_1391),
.Y(n_1439)
);

OAI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1379),
.A2(n_1364),
.B(n_1361),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1301),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1400),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1276),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1372),
.A2(n_1378),
.B1(n_1391),
.B2(n_1316),
.Y(n_1444)
);

INVx6_ASAP7_75t_L g1445 ( 
.A(n_1393),
.Y(n_1445)
);

BUFx2_ASAP7_75t_L g1446 ( 
.A(n_1253),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1292),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1368),
.Y(n_1448)
);

BUFx6f_ASAP7_75t_L g1449 ( 
.A(n_1335),
.Y(n_1449)
);

CKINVDCx20_ASAP7_75t_R g1450 ( 
.A(n_1307),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1372),
.A2(n_1316),
.B1(n_1323),
.B2(n_1288),
.Y(n_1451)
);

INVx1_ASAP7_75t_SL g1452 ( 
.A(n_1371),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1257),
.A2(n_1255),
.B1(n_1306),
.B2(n_1258),
.Y(n_1453)
);

INVx6_ASAP7_75t_L g1454 ( 
.A(n_1405),
.Y(n_1454)
);

CKINVDCx20_ASAP7_75t_R g1455 ( 
.A(n_1302),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1315),
.A2(n_1339),
.B1(n_1348),
.B2(n_1267),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1306),
.A2(n_1320),
.B1(n_1317),
.B2(n_1326),
.Y(n_1457)
);

OAI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1389),
.A2(n_1394),
.B1(n_1293),
.B2(n_1365),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_SL g1459 ( 
.A1(n_1376),
.A2(n_1406),
.B1(n_1387),
.B2(n_1395),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1330),
.A2(n_1342),
.B1(n_1341),
.B2(n_1283),
.Y(n_1460)
);

OAI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1365),
.A2(n_1287),
.B1(n_1371),
.B2(n_1350),
.Y(n_1461)
);

CKINVDCx16_ASAP7_75t_R g1462 ( 
.A(n_1405),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1289),
.A2(n_1344),
.B1(n_1386),
.B2(n_1345),
.Y(n_1463)
);

OAI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1309),
.A2(n_1252),
.B1(n_1392),
.B2(n_1396),
.Y(n_1464)
);

BUFx2_ASAP7_75t_SL g1465 ( 
.A(n_1254),
.Y(n_1465)
);

CKINVDCx11_ASAP7_75t_R g1466 ( 
.A(n_1343),
.Y(n_1466)
);

CKINVDCx6p67_ASAP7_75t_R g1467 ( 
.A(n_1275),
.Y(n_1467)
);

INVx6_ASAP7_75t_L g1468 ( 
.A(n_1353),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1349),
.B(n_1299),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1319),
.Y(n_1470)
);

BUFx4_ASAP7_75t_R g1471 ( 
.A(n_1374),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1309),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1334),
.A2(n_1331),
.B1(n_1254),
.B2(n_1358),
.Y(n_1473)
);

CKINVDCx6p67_ASAP7_75t_R g1474 ( 
.A(n_1308),
.Y(n_1474)
);

OAI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1359),
.A2(n_1357),
.B1(n_1279),
.B2(n_1353),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1362),
.B(n_1363),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1384),
.Y(n_1477)
);

BUFx8_ASAP7_75t_L g1478 ( 
.A(n_1383),
.Y(n_1478)
);

INVx2_ASAP7_75t_SL g1479 ( 
.A(n_1265),
.Y(n_1479)
);

AOI21xp5_ASAP7_75t_SL g1480 ( 
.A1(n_1359),
.A2(n_1264),
.B(n_1298),
.Y(n_1480)
);

BUFx3_ASAP7_75t_L g1481 ( 
.A(n_1333),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1395),
.A2(n_1384),
.B1(n_1406),
.B2(n_1376),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1328),
.B(n_1352),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1305),
.Y(n_1484)
);

BUFx6f_ASAP7_75t_L g1485 ( 
.A(n_1311),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1355),
.A2(n_1375),
.B1(n_1313),
.B2(n_1409),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_SL g1487 ( 
.A1(n_1376),
.A2(n_1406),
.B1(n_1328),
.B2(n_1261),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_SL g1488 ( 
.A1(n_1332),
.A2(n_1355),
.B1(n_1261),
.B2(n_1324),
.Y(n_1488)
);

INVx6_ASAP7_75t_L g1489 ( 
.A(n_1360),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1272),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_SL g1491 ( 
.A1(n_1324),
.A2(n_1397),
.B1(n_1282),
.B2(n_1329),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1329),
.A2(n_1325),
.B1(n_1271),
.B2(n_1340),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1340),
.A2(n_1337),
.B1(n_1322),
.B2(n_1369),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1381),
.A2(n_1407),
.B1(n_1268),
.B2(n_1294),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_SL g1495 ( 
.A1(n_1354),
.A2(n_1304),
.B1(n_1259),
.B2(n_1305),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1346),
.A2(n_1270),
.B1(n_1284),
.B2(n_1300),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1312),
.A2(n_1295),
.B1(n_1272),
.B2(n_1277),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1272),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1280),
.B(n_1263),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1338),
.A2(n_1399),
.B1(n_1377),
.B2(n_1260),
.Y(n_1500)
);

AOI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1281),
.A2(n_1278),
.B1(n_1262),
.B2(n_1274),
.Y(n_1501)
);

INVxp33_ASAP7_75t_L g1502 ( 
.A(n_1290),
.Y(n_1502)
);

AOI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1280),
.A2(n_1255),
.B(n_1369),
.Y(n_1503)
);

CKINVDCx20_ASAP7_75t_R g1504 ( 
.A(n_1280),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_SL g1505 ( 
.A1(n_1303),
.A2(n_960),
.B1(n_1380),
.B2(n_1327),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_1382),
.Y(n_1506)
);

BUFx4f_ASAP7_75t_SL g1507 ( 
.A(n_1336),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1347),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1347),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1273),
.Y(n_1510)
);

OAI21xp5_ASAP7_75t_SL g1511 ( 
.A1(n_1318),
.A2(n_691),
.B(n_662),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_1382),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1318),
.A2(n_1201),
.B1(n_1303),
.B2(n_1140),
.Y(n_1513)
);

CKINVDCx11_ASAP7_75t_R g1514 ( 
.A(n_1286),
.Y(n_1514)
);

INVx4_ASAP7_75t_L g1515 ( 
.A(n_1266),
.Y(n_1515)
);

BUFx2_ASAP7_75t_SL g1516 ( 
.A(n_1266),
.Y(n_1516)
);

BUFx12f_ASAP7_75t_L g1517 ( 
.A(n_1335),
.Y(n_1517)
);

CKINVDCx11_ASAP7_75t_R g1518 ( 
.A(n_1286),
.Y(n_1518)
);

BUFx10_ASAP7_75t_L g1519 ( 
.A(n_1382),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1366),
.A2(n_1318),
.B1(n_1380),
.B2(n_755),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1318),
.A2(n_1201),
.B1(n_1303),
.B2(n_1140),
.Y(n_1521)
);

CKINVDCx6p67_ASAP7_75t_R g1522 ( 
.A(n_1285),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1347),
.Y(n_1523)
);

BUFx6f_ASAP7_75t_L g1524 ( 
.A(n_1356),
.Y(n_1524)
);

CKINVDCx11_ASAP7_75t_R g1525 ( 
.A(n_1286),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1318),
.A2(n_1201),
.B1(n_1303),
.B2(n_1140),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1273),
.Y(n_1527)
);

BUFx6f_ASAP7_75t_SL g1528 ( 
.A(n_1266),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_SL g1529 ( 
.A1(n_1303),
.A2(n_960),
.B1(n_1380),
.B2(n_1327),
.Y(n_1529)
);

BUFx12f_ASAP7_75t_L g1530 ( 
.A(n_1335),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_1266),
.Y(n_1531)
);

OAI21xp5_ASAP7_75t_SL g1532 ( 
.A1(n_1318),
.A2(n_691),
.B(n_662),
.Y(n_1532)
);

OAI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1380),
.A2(n_960),
.B1(n_975),
.B2(n_1389),
.Y(n_1533)
);

CKINVDCx20_ASAP7_75t_R g1534 ( 
.A(n_1382),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1318),
.A2(n_1201),
.B1(n_1303),
.B2(n_1140),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1339),
.B(n_910),
.Y(n_1536)
);

INVx2_ASAP7_75t_SL g1537 ( 
.A(n_1286),
.Y(n_1537)
);

BUFx2_ASAP7_75t_L g1538 ( 
.A(n_1253),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1318),
.A2(n_1201),
.B1(n_1303),
.B2(n_1140),
.Y(n_1539)
);

BUFx12f_ASAP7_75t_L g1540 ( 
.A(n_1335),
.Y(n_1540)
);

CKINVDCx20_ASAP7_75t_R g1541 ( 
.A(n_1382),
.Y(n_1541)
);

INVx6_ASAP7_75t_L g1542 ( 
.A(n_1336),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1318),
.A2(n_1201),
.B1(n_1303),
.B2(n_1140),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1367),
.B(n_755),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1366),
.A2(n_1318),
.B1(n_1380),
.B2(n_755),
.Y(n_1545)
);

CKINVDCx6p67_ASAP7_75t_R g1546 ( 
.A(n_1285),
.Y(n_1546)
);

CKINVDCx20_ASAP7_75t_R g1547 ( 
.A(n_1382),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1382),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1318),
.A2(n_1201),
.B1(n_1303),
.B2(n_1140),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1266),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1253),
.Y(n_1551)
);

BUFx3_ASAP7_75t_L g1552 ( 
.A(n_1266),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1484),
.Y(n_1553)
);

AOI21xp33_ASAP7_75t_SL g1554 ( 
.A1(n_1520),
.A2(n_1545),
.B(n_1415),
.Y(n_1554)
);

OAI21xp33_ASAP7_75t_SL g1555 ( 
.A1(n_1480),
.A2(n_1417),
.B(n_1440),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1483),
.B(n_1499),
.Y(n_1556)
);

INVx1_ASAP7_75t_SL g1557 ( 
.A(n_1446),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1418),
.B(n_1487),
.Y(n_1558)
);

OR2x6_ASAP7_75t_L g1559 ( 
.A(n_1503),
.B(n_1486),
.Y(n_1559)
);

INVx2_ASAP7_75t_SL g1560 ( 
.A(n_1445),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1477),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1477),
.Y(n_1562)
);

OAI21x1_ASAP7_75t_L g1563 ( 
.A1(n_1500),
.A2(n_1493),
.B(n_1496),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1544),
.B(n_1432),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1490),
.Y(n_1565)
);

INVx4_ASAP7_75t_L g1566 ( 
.A(n_1489),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1447),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1498),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1418),
.B(n_1487),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1504),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1432),
.B(n_1439),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1482),
.B(n_1426),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1459),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1459),
.B(n_1422),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1422),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1482),
.B(n_1426),
.Y(n_1576)
);

INVxp67_ASAP7_75t_L g1577 ( 
.A(n_1448),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1502),
.B(n_1469),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_L g1579 ( 
.A(n_1434),
.B(n_1536),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1510),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1417),
.B(n_1451),
.Y(n_1581)
);

AO21x2_ASAP7_75t_L g1582 ( 
.A1(n_1501),
.A2(n_1497),
.B(n_1533),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1452),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1527),
.Y(n_1584)
);

INVx6_ASAP7_75t_L g1585 ( 
.A(n_1414),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1451),
.B(n_1472),
.Y(n_1586)
);

AO21x2_ASAP7_75t_L g1587 ( 
.A1(n_1533),
.A2(n_1461),
.B(n_1458),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1470),
.Y(n_1588)
);

OAI21x1_ASAP7_75t_L g1589 ( 
.A1(n_1500),
.A2(n_1493),
.B(n_1496),
.Y(n_1589)
);

BUFx3_ASAP7_75t_L g1590 ( 
.A(n_1445),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1444),
.B(n_1453),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1488),
.Y(n_1592)
);

AOI21x1_ASAP7_75t_L g1593 ( 
.A1(n_1463),
.A2(n_1473),
.B(n_1475),
.Y(n_1593)
);

NOR2x1_ASAP7_75t_R g1594 ( 
.A(n_1517),
.B(n_1530),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_1443),
.Y(n_1595)
);

BUFx4f_ASAP7_75t_SL g1596 ( 
.A(n_1540),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1444),
.B(n_1453),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1505),
.B(n_1529),
.Y(n_1598)
);

OAI21x1_ASAP7_75t_L g1599 ( 
.A1(n_1494),
.A2(n_1492),
.B(n_1457),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1538),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1464),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1464),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1551),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1436),
.Y(n_1604)
);

OAI21x1_ASAP7_75t_L g1605 ( 
.A1(n_1494),
.A2(n_1492),
.B(n_1457),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1476),
.Y(n_1606)
);

OAI21xp33_ASAP7_75t_L g1607 ( 
.A1(n_1513),
.A2(n_1521),
.B(n_1535),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1513),
.A2(n_1539),
.B1(n_1543),
.B2(n_1521),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1441),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1439),
.B(n_1461),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1442),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1491),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1491),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_L g1614 ( 
.A(n_1455),
.B(n_1412),
.Y(n_1614)
);

OA21x2_ASAP7_75t_L g1615 ( 
.A1(n_1526),
.A2(n_1539),
.B(n_1535),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1495),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1495),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1508),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1509),
.Y(n_1619)
);

AO21x2_ASAP7_75t_L g1620 ( 
.A1(n_1458),
.A2(n_1456),
.B(n_1511),
.Y(n_1620)
);

NAND2xp33_ASAP7_75t_L g1621 ( 
.A(n_1526),
.B(n_1543),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1523),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_1506),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1549),
.B(n_1532),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1460),
.Y(n_1625)
);

BUFx3_ASAP7_75t_L g1626 ( 
.A(n_1445),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1460),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1481),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1505),
.B(n_1529),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1489),
.Y(n_1630)
);

BUFx4f_ASAP7_75t_SL g1631 ( 
.A(n_1534),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1479),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1489),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1412),
.B(n_1548),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1485),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1549),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1429),
.B(n_1474),
.Y(n_1637)
);

AND2x4_ASAP7_75t_L g1638 ( 
.A(n_1435),
.B(n_1537),
.Y(n_1638)
);

AO21x2_ASAP7_75t_L g1639 ( 
.A1(n_1471),
.A2(n_1465),
.B(n_1468),
.Y(n_1639)
);

BUFx12f_ASAP7_75t_L g1640 ( 
.A(n_1431),
.Y(n_1640)
);

NAND2x1p5_ASAP7_75t_L g1641 ( 
.A(n_1421),
.B(n_1430),
.Y(n_1641)
);

INVx3_ASAP7_75t_L g1642 ( 
.A(n_1454),
.Y(n_1642)
);

OAI21x1_ASAP7_75t_L g1643 ( 
.A1(n_1454),
.A2(n_1471),
.B(n_1467),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1431),
.B(n_1449),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1454),
.Y(n_1645)
);

OAI21x1_ASAP7_75t_L g1646 ( 
.A1(n_1528),
.A2(n_1413),
.B(n_1542),
.Y(n_1646)
);

INVx2_ASAP7_75t_SL g1647 ( 
.A(n_1428),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1423),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1528),
.Y(n_1649)
);

BUFx3_ASAP7_75t_L g1650 ( 
.A(n_1450),
.Y(n_1650)
);

AO21x1_ASAP7_75t_L g1651 ( 
.A1(n_1421),
.A2(n_1515),
.B(n_1433),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1466),
.A2(n_1413),
.B1(n_1542),
.B2(n_1416),
.Y(n_1652)
);

INVx2_ASAP7_75t_SL g1653 ( 
.A(n_1416),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1512),
.B(n_1541),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1430),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1552),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1424),
.Y(n_1657)
);

INVx2_ASAP7_75t_SL g1658 ( 
.A(n_1437),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1516),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1462),
.B(n_1524),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1507),
.A2(n_1420),
.B1(n_1427),
.B2(n_1522),
.Y(n_1661)
);

A2O1A1Ixp33_ASAP7_75t_L g1662 ( 
.A1(n_1555),
.A2(n_1524),
.B(n_1431),
.C(n_1449),
.Y(n_1662)
);

OAI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1554),
.A2(n_1547),
.B(n_1531),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1570),
.B(n_1578),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1570),
.B(n_1449),
.Y(n_1665)
);

AO32x2_ASAP7_75t_L g1666 ( 
.A1(n_1608),
.A2(n_1556),
.A3(n_1566),
.B1(n_1560),
.B2(n_1573),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1578),
.B(n_1449),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1646),
.B(n_1550),
.Y(n_1668)
);

NAND2x1p5_ASAP7_75t_L g1669 ( 
.A(n_1566),
.B(n_1524),
.Y(n_1669)
);

BUFx12f_ASAP7_75t_L g1670 ( 
.A(n_1640),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1579),
.B(n_1524),
.Y(n_1671)
);

AOI221xp5_ASAP7_75t_L g1672 ( 
.A1(n_1554),
.A2(n_1431),
.B1(n_1437),
.B2(n_1518),
.C(n_1425),
.Y(n_1672)
);

OAI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1555),
.A2(n_1519),
.B(n_1525),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1606),
.B(n_1519),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1586),
.B(n_1546),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1559),
.A2(n_1420),
.B(n_1507),
.Y(n_1676)
);

OA21x2_ASAP7_75t_L g1677 ( 
.A1(n_1563),
.A2(n_1438),
.B(n_1514),
.Y(n_1677)
);

OAI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1621),
.A2(n_1414),
.B(n_1419),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1607),
.B(n_1478),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1624),
.B(n_1478),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1586),
.B(n_1575),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1564),
.B(n_1583),
.Y(n_1682)
);

INVx1_ASAP7_75t_SL g1683 ( 
.A(n_1557),
.Y(n_1683)
);

AO21x2_ASAP7_75t_L g1684 ( 
.A1(n_1563),
.A2(n_1589),
.B(n_1587),
.Y(n_1684)
);

OR2x6_ASAP7_75t_L g1685 ( 
.A(n_1559),
.B(n_1643),
.Y(n_1685)
);

AND2x4_ASAP7_75t_L g1686 ( 
.A(n_1646),
.B(n_1580),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1559),
.A2(n_1605),
.B(n_1599),
.Y(n_1687)
);

AOI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1607),
.A2(n_1620),
.B1(n_1598),
.B2(n_1629),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_SL g1689 ( 
.A(n_1595),
.B(n_1623),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1575),
.B(n_1592),
.Y(n_1690)
);

OAI21x1_ASAP7_75t_L g1691 ( 
.A1(n_1589),
.A2(n_1605),
.B(n_1599),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1600),
.B(n_1603),
.Y(n_1692)
);

O2A1O1Ixp33_ASAP7_75t_SL g1693 ( 
.A1(n_1636),
.A2(n_1637),
.B(n_1592),
.C(n_1630),
.Y(n_1693)
);

INVx2_ASAP7_75t_SL g1694 ( 
.A(n_1567),
.Y(n_1694)
);

AO32x1_ASAP7_75t_L g1695 ( 
.A1(n_1598),
.A2(n_1629),
.A3(n_1569),
.B1(n_1558),
.B2(n_1574),
.Y(n_1695)
);

AOI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1559),
.A2(n_1587),
.B(n_1620),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1577),
.B(n_1571),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1580),
.B(n_1584),
.Y(n_1698)
);

AO32x2_ASAP7_75t_L g1699 ( 
.A1(n_1566),
.A2(n_1560),
.A3(n_1573),
.B1(n_1587),
.B2(n_1574),
.Y(n_1699)
);

AOI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1559),
.A2(n_1620),
.B(n_1639),
.Y(n_1700)
);

OAI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1615),
.A2(n_1636),
.B1(n_1610),
.B2(n_1581),
.Y(n_1701)
);

OR2x6_ASAP7_75t_L g1702 ( 
.A(n_1643),
.B(n_1593),
.Y(n_1702)
);

AOI221x1_ASAP7_75t_SL g1703 ( 
.A1(n_1612),
.A2(n_1613),
.B1(n_1601),
.B2(n_1602),
.C(n_1617),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1610),
.B(n_1572),
.Y(n_1704)
);

O2A1O1Ixp33_ASAP7_75t_L g1705 ( 
.A1(n_1591),
.A2(n_1597),
.B(n_1581),
.C(n_1615),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1639),
.B(n_1644),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1553),
.Y(n_1707)
);

OA21x2_ASAP7_75t_L g1708 ( 
.A1(n_1616),
.A2(n_1617),
.B(n_1612),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1639),
.B(n_1644),
.Y(n_1709)
);

OR2x2_ASAP7_75t_L g1710 ( 
.A(n_1572),
.B(n_1576),
.Y(n_1710)
);

OA21x2_ASAP7_75t_L g1711 ( 
.A1(n_1616),
.A2(n_1613),
.B(n_1602),
.Y(n_1711)
);

AOI221xp5_ASAP7_75t_L g1712 ( 
.A1(n_1591),
.A2(n_1597),
.B1(n_1569),
.B2(n_1558),
.C(n_1627),
.Y(n_1712)
);

AO21x2_ASAP7_75t_L g1713 ( 
.A1(n_1582),
.A2(n_1593),
.B(n_1561),
.Y(n_1713)
);

AO21x1_ASAP7_75t_L g1714 ( 
.A1(n_1566),
.A2(n_1630),
.B(n_1633),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1615),
.A2(n_1576),
.B1(n_1627),
.B2(n_1625),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1625),
.B(n_1562),
.Y(n_1716)
);

CKINVDCx20_ASAP7_75t_R g1717 ( 
.A(n_1631),
.Y(n_1717)
);

OA21x2_ASAP7_75t_L g1718 ( 
.A1(n_1562),
.A2(n_1565),
.B(n_1568),
.Y(n_1718)
);

OAI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1615),
.A2(n_1652),
.B1(n_1585),
.B2(n_1649),
.Y(n_1719)
);

OAI221xp5_ASAP7_75t_L g1720 ( 
.A1(n_1653),
.A2(n_1614),
.B1(n_1660),
.B2(n_1649),
.C(n_1650),
.Y(n_1720)
);

AOI221xp5_ASAP7_75t_L g1721 ( 
.A1(n_1582),
.A2(n_1638),
.B1(n_1632),
.B2(n_1611),
.C(n_1622),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1585),
.A2(n_1653),
.B1(n_1657),
.B2(n_1659),
.Y(n_1722)
);

INVxp67_ASAP7_75t_L g1723 ( 
.A(n_1711),
.Y(n_1723)
);

INVx3_ASAP7_75t_L g1724 ( 
.A(n_1686),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1707),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1706),
.B(n_1709),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1711),
.B(n_1582),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1707),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1684),
.B(n_1568),
.Y(n_1729)
);

INVx2_ASAP7_75t_SL g1730 ( 
.A(n_1686),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1708),
.B(n_1588),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1681),
.B(n_1635),
.Y(n_1732)
);

INVx2_ASAP7_75t_SL g1733 ( 
.A(n_1686),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1718),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1718),
.Y(n_1735)
);

HB1xp67_ASAP7_75t_L g1736 ( 
.A(n_1718),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1684),
.B(n_1609),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_SL g1738 ( 
.A1(n_1696),
.A2(n_1585),
.B1(n_1640),
.B2(n_1650),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1699),
.B(n_1604),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1699),
.B(n_1638),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1708),
.B(n_1618),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1699),
.B(n_1638),
.Y(n_1742)
);

OAI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1688),
.A2(n_1585),
.B1(n_1660),
.B2(n_1650),
.Y(n_1743)
);

CKINVDCx14_ASAP7_75t_R g1744 ( 
.A(n_1717),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1698),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1699),
.B(n_1664),
.Y(n_1746)
);

HB1xp67_ASAP7_75t_L g1747 ( 
.A(n_1694),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1710),
.B(n_1628),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1691),
.B(n_1687),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1691),
.B(n_1619),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1685),
.B(n_1619),
.Y(n_1751)
);

NOR2x1p5_ASAP7_75t_L g1752 ( 
.A(n_1670),
.B(n_1626),
.Y(n_1752)
);

INVxp67_ASAP7_75t_SL g1753 ( 
.A(n_1716),
.Y(n_1753)
);

NOR2x1_ASAP7_75t_L g1754 ( 
.A(n_1741),
.B(n_1713),
.Y(n_1754)
);

INVx4_ASAP7_75t_L g1755 ( 
.A(n_1748),
.Y(n_1755)
);

OAI21xp33_ASAP7_75t_SL g1756 ( 
.A1(n_1740),
.A2(n_1721),
.B(n_1695),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1740),
.B(n_1700),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1725),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1725),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1753),
.B(n_1715),
.Y(n_1760)
);

OAI21xp33_ASAP7_75t_L g1761 ( 
.A1(n_1743),
.A2(n_1712),
.B(n_1679),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1728),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1742),
.B(n_1685),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1727),
.B(n_1677),
.Y(n_1764)
);

NAND2x1p5_ASAP7_75t_SL g1765 ( 
.A(n_1749),
.B(n_1679),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1742),
.B(n_1739),
.Y(n_1766)
);

OAI211xp5_ASAP7_75t_SL g1767 ( 
.A1(n_1738),
.A2(n_1672),
.B(n_1697),
.C(n_1678),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1746),
.B(n_1715),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1735),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1728),
.Y(n_1770)
);

HB1xp67_ASAP7_75t_L g1771 ( 
.A(n_1723),
.Y(n_1771)
);

OAI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1743),
.A2(n_1662),
.B1(n_1695),
.B2(n_1705),
.Y(n_1772)
);

NAND3xp33_ASAP7_75t_SL g1773 ( 
.A(n_1738),
.B(n_1662),
.C(n_1673),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1739),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1746),
.B(n_1685),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1737),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1726),
.B(n_1666),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1748),
.A2(n_1701),
.B1(n_1704),
.B2(n_1690),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1744),
.B(n_1720),
.Y(n_1779)
);

AND2x4_ASAP7_75t_SL g1780 ( 
.A(n_1747),
.B(n_1702),
.Y(n_1780)
);

INVx1_ASAP7_75t_SL g1781 ( 
.A(n_1747),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1724),
.B(n_1666),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1723),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1730),
.B(n_1666),
.Y(n_1784)
);

INVx4_ASAP7_75t_L g1785 ( 
.A(n_1751),
.Y(n_1785)
);

NAND2x1p5_ASAP7_75t_L g1786 ( 
.A(n_1737),
.B(n_1677),
.Y(n_1786)
);

BUFx3_ASAP7_75t_L g1787 ( 
.A(n_1751),
.Y(n_1787)
);

OAI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1727),
.A2(n_1695),
.B1(n_1705),
.B2(n_1701),
.Y(n_1788)
);

HB1xp67_ASAP7_75t_L g1789 ( 
.A(n_1734),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1758),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1758),
.Y(n_1791)
);

AND2x4_ASAP7_75t_L g1792 ( 
.A(n_1785),
.B(n_1730),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1768),
.B(n_1729),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1774),
.B(n_1731),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1759),
.Y(n_1795)
);

NOR2xp67_ASAP7_75t_L g1796 ( 
.A(n_1785),
.B(n_1734),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1766),
.B(n_1733),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1766),
.B(n_1733),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1766),
.B(n_1733),
.Y(n_1799)
);

AND2x4_ASAP7_75t_SL g1800 ( 
.A(n_1755),
.B(n_1668),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1769),
.Y(n_1801)
);

INVx3_ASAP7_75t_L g1802 ( 
.A(n_1785),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1759),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1776),
.B(n_1731),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1776),
.B(n_1736),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1782),
.B(n_1784),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1769),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1768),
.B(n_1729),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1762),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1784),
.B(n_1745),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1762),
.Y(n_1811)
);

INVx4_ASAP7_75t_L g1812 ( 
.A(n_1755),
.Y(n_1812)
);

NAND2x1p5_ASAP7_75t_L g1813 ( 
.A(n_1754),
.B(n_1677),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1776),
.B(n_1736),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1760),
.B(n_1729),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_1779),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1784),
.B(n_1751),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_SL g1818 ( 
.A(n_1772),
.B(n_1714),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1775),
.B(n_1732),
.Y(n_1819)
);

INVx3_ASAP7_75t_SL g1820 ( 
.A(n_1780),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1775),
.B(n_1732),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1770),
.Y(n_1822)
);

AND2x4_ASAP7_75t_L g1823 ( 
.A(n_1785),
.B(n_1750),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1820),
.B(n_1800),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1820),
.B(n_1775),
.Y(n_1825)
);

INVx2_ASAP7_75t_SL g1826 ( 
.A(n_1800),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1820),
.B(n_1757),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1818),
.B(n_1755),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1820),
.B(n_1757),
.Y(n_1829)
);

INVxp67_ASAP7_75t_SL g1830 ( 
.A(n_1818),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1800),
.B(n_1757),
.Y(n_1831)
);

OAI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1813),
.A2(n_1756),
.B(n_1788),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1793),
.B(n_1760),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1793),
.B(n_1755),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1806),
.B(n_1792),
.Y(n_1835)
);

OAI32xp33_ASAP7_75t_L g1836 ( 
.A1(n_1813),
.A2(n_1756),
.A3(n_1772),
.B1(n_1788),
.B2(n_1761),
.Y(n_1836)
);

AND2x4_ASAP7_75t_L g1837 ( 
.A(n_1812),
.B(n_1796),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1808),
.B(n_1815),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1806),
.B(n_1763),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1808),
.B(n_1764),
.Y(n_1840)
);

NOR2x1p5_ASAP7_75t_L g1841 ( 
.A(n_1816),
.B(n_1773),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1790),
.Y(n_1842)
);

HB1xp67_ASAP7_75t_L g1843 ( 
.A(n_1790),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1791),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1815),
.B(n_1764),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1791),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1806),
.B(n_1763),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1795),
.Y(n_1848)
);

A2O1A1Ixp33_ASAP7_75t_L g1849 ( 
.A1(n_1796),
.A2(n_1761),
.B(n_1767),
.C(n_1773),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1801),
.Y(n_1850)
);

OAI21xp33_ASAP7_75t_SL g1851 ( 
.A1(n_1812),
.A2(n_1755),
.B(n_1785),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1795),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1819),
.B(n_1777),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1803),
.Y(n_1854)
);

INVx2_ASAP7_75t_SL g1855 ( 
.A(n_1802),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1803),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1809),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1792),
.B(n_1763),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1794),
.B(n_1764),
.Y(n_1859)
);

INVx2_ASAP7_75t_SL g1860 ( 
.A(n_1802),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1809),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1811),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1811),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1822),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1792),
.B(n_1777),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1822),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1810),
.Y(n_1867)
);

AND2x4_ASAP7_75t_L g1868 ( 
.A(n_1812),
.B(n_1780),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1801),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1830),
.B(n_1819),
.Y(n_1870)
);

AND3x2_ASAP7_75t_L g1871 ( 
.A(n_1824),
.B(n_1689),
.C(n_1837),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1839),
.B(n_1847),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1843),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1842),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1835),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1849),
.B(n_1819),
.Y(n_1876)
);

INVx1_ASAP7_75t_SL g1877 ( 
.A(n_1824),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1842),
.Y(n_1878)
);

OAI31xp33_ASAP7_75t_L g1879 ( 
.A1(n_1841),
.A2(n_1767),
.A3(n_1813),
.B(n_1802),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1853),
.B(n_1794),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1839),
.B(n_1802),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1847),
.B(n_1802),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1844),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_L g1884 ( 
.A(n_1836),
.B(n_1596),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1825),
.B(n_1817),
.Y(n_1885)
);

AND2x4_ASAP7_75t_L g1886 ( 
.A(n_1835),
.B(n_1812),
.Y(n_1886)
);

NAND4xp25_ASAP7_75t_L g1887 ( 
.A(n_1836),
.B(n_1663),
.C(n_1778),
.D(n_1703),
.Y(n_1887)
);

NOR2xp67_ASAP7_75t_SL g1888 ( 
.A(n_1828),
.B(n_1670),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1833),
.B(n_1821),
.Y(n_1889)
);

AOI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1832),
.A2(n_1719),
.B1(n_1778),
.B2(n_1812),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1825),
.B(n_1827),
.Y(n_1891)
);

INVxp67_ASAP7_75t_L g1892 ( 
.A(n_1827),
.Y(n_1892)
);

AND2x2_ASAP7_75t_SL g1893 ( 
.A(n_1868),
.B(n_1671),
.Y(n_1893)
);

CKINVDCx16_ASAP7_75t_R g1894 ( 
.A(n_1829),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1833),
.B(n_1821),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1829),
.B(n_1817),
.Y(n_1896)
);

INVx1_ASAP7_75t_SL g1897 ( 
.A(n_1868),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1838),
.B(n_1794),
.Y(n_1898)
);

AOI21xp33_ASAP7_75t_SL g1899 ( 
.A1(n_1826),
.A2(n_1661),
.B(n_1765),
.Y(n_1899)
);

NOR2xp67_ASAP7_75t_SL g1900 ( 
.A(n_1826),
.B(n_1623),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1858),
.B(n_1831),
.Y(n_1901)
);

AND2x4_ASAP7_75t_L g1902 ( 
.A(n_1868),
.B(n_1792),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1858),
.B(n_1817),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1838),
.B(n_1821),
.Y(n_1904)
);

AOI22xp33_ASAP7_75t_L g1905 ( 
.A1(n_1831),
.A2(n_1834),
.B1(n_1837),
.B2(n_1702),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1844),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1846),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1874),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1874),
.Y(n_1909)
);

OAI22xp33_ASAP7_75t_L g1910 ( 
.A1(n_1887),
.A2(n_1890),
.B1(n_1876),
.B2(n_1894),
.Y(n_1910)
);

NOR3xp33_ASAP7_75t_L g1911 ( 
.A(n_1884),
.B(n_1851),
.C(n_1594),
.Y(n_1911)
);

OAI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1879),
.A2(n_1813),
.B(n_1680),
.Y(n_1912)
);

OR2x2_ASAP7_75t_L g1913 ( 
.A(n_1870),
.B(n_1840),
.Y(n_1913)
);

OAI22xp5_ASAP7_75t_L g1914 ( 
.A1(n_1877),
.A2(n_1893),
.B1(n_1897),
.B2(n_1899),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1892),
.B(n_1865),
.Y(n_1915)
);

NAND3xp33_ASAP7_75t_L g1916 ( 
.A(n_1888),
.B(n_1840),
.C(n_1845),
.Y(n_1916)
);

OAI22xp33_ASAP7_75t_L g1917 ( 
.A1(n_1875),
.A2(n_1845),
.B1(n_1867),
.B2(n_1786),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1878),
.Y(n_1918)
);

OAI22xp33_ASAP7_75t_L g1919 ( 
.A1(n_1875),
.A2(n_1786),
.B1(n_1787),
.B2(n_1859),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1878),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1891),
.B(n_1872),
.Y(n_1921)
);

OAI21xp33_ASAP7_75t_L g1922 ( 
.A1(n_1891),
.A2(n_1859),
.B(n_1865),
.Y(n_1922)
);

AOI221x1_ASAP7_75t_L g1923 ( 
.A1(n_1873),
.A2(n_1837),
.B1(n_1866),
.B2(n_1848),
.C(n_1846),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1883),
.Y(n_1924)
);

INVxp67_ASAP7_75t_L g1925 ( 
.A(n_1900),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1883),
.Y(n_1926)
);

INVxp67_ASAP7_75t_L g1927 ( 
.A(n_1900),
.Y(n_1927)
);

AOI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1893),
.A2(n_1792),
.B1(n_1823),
.B2(n_1668),
.Y(n_1928)
);

OAI22xp5_ASAP7_75t_L g1929 ( 
.A1(n_1905),
.A2(n_1895),
.B1(n_1889),
.B2(n_1902),
.Y(n_1929)
);

O2A1O1Ixp33_ASAP7_75t_L g1930 ( 
.A1(n_1873),
.A2(n_1860),
.B(n_1855),
.C(n_1665),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1906),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1901),
.B(n_1810),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1872),
.B(n_1852),
.Y(n_1933)
);

XNOR2x1_ASAP7_75t_L g1934 ( 
.A(n_1871),
.B(n_1752),
.Y(n_1934)
);

OAI21xp33_ASAP7_75t_L g1935 ( 
.A1(n_1910),
.A2(n_1901),
.B(n_1904),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_L g1936 ( 
.A(n_1925),
.B(n_1888),
.Y(n_1936)
);

OAI22xp33_ASAP7_75t_L g1937 ( 
.A1(n_1923),
.A2(n_1898),
.B1(n_1880),
.B2(n_1786),
.Y(n_1937)
);

AOI222xp33_ASAP7_75t_L g1938 ( 
.A1(n_1914),
.A2(n_1885),
.B1(n_1896),
.B2(n_1903),
.C1(n_1886),
.C2(n_1882),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1932),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1927),
.B(n_1885),
.Y(n_1940)
);

OAI22xp5_ASAP7_75t_L g1941 ( 
.A1(n_1916),
.A2(n_1902),
.B1(n_1886),
.B2(n_1903),
.Y(n_1941)
);

AOI222xp33_ASAP7_75t_L g1942 ( 
.A1(n_1914),
.A2(n_1896),
.B1(n_1886),
.B2(n_1881),
.C1(n_1882),
.C2(n_1907),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1908),
.Y(n_1943)
);

AOI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1911),
.A2(n_1934),
.B1(n_1929),
.B2(n_1912),
.Y(n_1944)
);

NAND4xp25_ASAP7_75t_SL g1945 ( 
.A(n_1912),
.B(n_1881),
.C(n_1880),
.D(n_1898),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1909),
.Y(n_1946)
);

NOR2xp33_ASAP7_75t_L g1947 ( 
.A(n_1921),
.B(n_1594),
.Y(n_1947)
);

OAI332xp33_ASAP7_75t_L g1948 ( 
.A1(n_1915),
.A2(n_1907),
.A3(n_1906),
.B1(n_1860),
.B2(n_1855),
.B3(n_1683),
.C1(n_1848),
.C2(n_1862),
.Y(n_1948)
);

AOI321xp33_ASAP7_75t_L g1949 ( 
.A1(n_1922),
.A2(n_1902),
.A3(n_1680),
.B1(n_1754),
.B2(n_1675),
.C(n_1692),
.Y(n_1949)
);

AOI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1928),
.A2(n_1854),
.B1(n_1856),
.B2(n_1864),
.Y(n_1950)
);

AND2x4_ASAP7_75t_L g1951 ( 
.A(n_1918),
.B(n_1857),
.Y(n_1951)
);

OAI22xp5_ASAP7_75t_L g1952 ( 
.A1(n_1913),
.A2(n_1786),
.B1(n_1752),
.B2(n_1823),
.Y(n_1952)
);

NOR2x1_ASAP7_75t_L g1953 ( 
.A(n_1920),
.B(n_1717),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1933),
.B(n_1810),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1924),
.Y(n_1955)
);

AOI22xp5_ASAP7_75t_L g1956 ( 
.A1(n_1945),
.A2(n_1917),
.B1(n_1919),
.B2(n_1931),
.Y(n_1956)
);

O2A1O1Ixp33_ASAP7_75t_L g1957 ( 
.A1(n_1937),
.A2(n_1926),
.B(n_1930),
.C(n_1771),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1935),
.B(n_1861),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1951),
.Y(n_1959)
);

AOI21xp33_ASAP7_75t_SL g1960 ( 
.A1(n_1941),
.A2(n_1595),
.B(n_1634),
.Y(n_1960)
);

AOI21xp5_ASAP7_75t_SL g1961 ( 
.A1(n_1936),
.A2(n_1654),
.B(n_1658),
.Y(n_1961)
);

AND2x4_ASAP7_75t_L g1962 ( 
.A(n_1953),
.B(n_1863),
.Y(n_1962)
);

O2A1O1Ixp33_ASAP7_75t_L g1963 ( 
.A1(n_1942),
.A2(n_1783),
.B(n_1771),
.C(n_1658),
.Y(n_1963)
);

NAND4xp75_ASAP7_75t_SL g1964 ( 
.A(n_1947),
.B(n_1799),
.C(n_1798),
.D(n_1797),
.Y(n_1964)
);

NOR2xp33_ASAP7_75t_L g1965 ( 
.A(n_1940),
.B(n_1674),
.Y(n_1965)
);

AOI21xp5_ASAP7_75t_L g1966 ( 
.A1(n_1948),
.A2(n_1866),
.B(n_1862),
.Y(n_1966)
);

NAND3xp33_ASAP7_75t_L g1967 ( 
.A(n_1938),
.B(n_1869),
.C(n_1850),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1951),
.Y(n_1968)
);

NAND2xp33_ASAP7_75t_SL g1969 ( 
.A(n_1962),
.B(n_1939),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_SL g1970 ( 
.A(n_1962),
.B(n_1949),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1959),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1968),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1958),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1967),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1965),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1960),
.B(n_1944),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1966),
.Y(n_1977)
);

NOR2xp33_ASAP7_75t_L g1978 ( 
.A(n_1961),
.B(n_1943),
.Y(n_1978)
);

AOI21xp5_ASAP7_75t_L g1979 ( 
.A1(n_1957),
.A2(n_1955),
.B(n_1946),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_L g1980 ( 
.A(n_1956),
.B(n_1950),
.Y(n_1980)
);

O2A1O1Ixp33_ASAP7_75t_L g1981 ( 
.A1(n_1977),
.A2(n_1963),
.B(n_1952),
.C(n_1949),
.Y(n_1981)
);

AOI221xp5_ASAP7_75t_L g1982 ( 
.A1(n_1980),
.A2(n_1954),
.B1(n_1964),
.B2(n_1869),
.C(n_1850),
.Y(n_1982)
);

INVxp67_ASAP7_75t_L g1983 ( 
.A(n_1969),
.Y(n_1983)
);

O2A1O1Ixp33_ASAP7_75t_L g1984 ( 
.A1(n_1974),
.A2(n_1783),
.B(n_1693),
.C(n_1789),
.Y(n_1984)
);

NAND4xp75_ASAP7_75t_L g1985 ( 
.A(n_1970),
.B(n_1651),
.C(n_1676),
.D(n_1657),
.Y(n_1985)
);

O2A1O1Ixp33_ASAP7_75t_L g1986 ( 
.A1(n_1980),
.A2(n_1693),
.B(n_1789),
.C(n_1645),
.Y(n_1986)
);

CKINVDCx5p33_ASAP7_75t_R g1987 ( 
.A(n_1983),
.Y(n_1987)
);

AOI221xp5_ASAP7_75t_L g1988 ( 
.A1(n_1981),
.A2(n_1979),
.B1(n_1978),
.B2(n_1973),
.C(n_1976),
.Y(n_1988)
);

OAI22xp33_ASAP7_75t_R g1989 ( 
.A1(n_1985),
.A2(n_1972),
.B1(n_1971),
.B2(n_1975),
.Y(n_1989)
);

OAI22xp33_ASAP7_75t_L g1990 ( 
.A1(n_1982),
.A2(n_1978),
.B1(n_1805),
.B2(n_1814),
.Y(n_1990)
);

NAND3xp33_ASAP7_75t_SL g1991 ( 
.A(n_1984),
.B(n_1651),
.C(n_1669),
.Y(n_1991)
);

NAND3xp33_ASAP7_75t_SL g1992 ( 
.A(n_1986),
.B(n_1669),
.C(n_1641),
.Y(n_1992)
);

OAI211xp5_ASAP7_75t_L g1993 ( 
.A1(n_1983),
.A2(n_1590),
.B(n_1626),
.C(n_1648),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1987),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1988),
.B(n_1823),
.Y(n_1995)
);

CKINVDCx14_ASAP7_75t_R g1996 ( 
.A(n_1991),
.Y(n_1996)
);

OAI211xp5_ASAP7_75t_L g1997 ( 
.A1(n_1993),
.A2(n_1626),
.B(n_1590),
.C(n_1642),
.Y(n_1997)
);

AOI21xp5_ASAP7_75t_L g1998 ( 
.A1(n_1990),
.A2(n_1642),
.B(n_1682),
.Y(n_1998)
);

NAND4xp75_ASAP7_75t_L g1999 ( 
.A(n_1989),
.B(n_1659),
.C(n_1647),
.D(n_1667),
.Y(n_1999)
);

NOR2x1p5_ASAP7_75t_L g2000 ( 
.A(n_1999),
.B(n_1992),
.Y(n_2000)
);

NAND4xp25_ASAP7_75t_L g2001 ( 
.A(n_1995),
.B(n_1590),
.C(n_1642),
.D(n_1722),
.Y(n_2001)
);

AOI22xp5_ASAP7_75t_L g2002 ( 
.A1(n_1994),
.A2(n_1823),
.B1(n_1668),
.B2(n_1656),
.Y(n_2002)
);

INVx1_ASAP7_75t_SL g2003 ( 
.A(n_1998),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_2000),
.Y(n_2004)
);

AOI22xp5_ASAP7_75t_L g2005 ( 
.A1(n_2004),
.A2(n_1996),
.B1(n_2001),
.B2(n_2003),
.Y(n_2005)
);

XNOR2x1_ASAP7_75t_L g2006 ( 
.A(n_2005),
.B(n_2002),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_2005),
.B(n_1997),
.Y(n_2007)
);

OAI22xp5_ASAP7_75t_L g2008 ( 
.A1(n_2007),
.A2(n_1814),
.B1(n_1805),
.B2(n_1804),
.Y(n_2008)
);

OAI31xp33_ASAP7_75t_L g2009 ( 
.A1(n_2006),
.A2(n_1641),
.A3(n_1823),
.B(n_1781),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_2008),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_2009),
.Y(n_2011)
);

AOI221xp5_ASAP7_75t_L g2012 ( 
.A1(n_2010),
.A2(n_1807),
.B1(n_1801),
.B2(n_1765),
.C(n_1781),
.Y(n_2012)
);

XNOR2xp5_ASAP7_75t_L g2013 ( 
.A(n_2012),
.B(n_2011),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_2013),
.Y(n_2014)
);

OAI221xp5_ASAP7_75t_R g2015 ( 
.A1(n_2014),
.A2(n_1765),
.B1(n_1814),
.B2(n_1805),
.C(n_1807),
.Y(n_2015)
);

AOI211xp5_ASAP7_75t_L g2016 ( 
.A1(n_2015),
.A2(n_1647),
.B(n_1655),
.C(n_1656),
.Y(n_2016)
);


endmodule