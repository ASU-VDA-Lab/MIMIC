module fake_jpeg_17753_n_86 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_86);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_86;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx6_ASAP7_75t_SL g14 ( 
.A(n_7),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx4_ASAP7_75t_SL g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_15),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_19),
.B1(n_20),
.B2(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_2),
.Y(n_27)
);

AO21x1_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_31),
.B(n_32),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_22),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_3),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_19),
.Y(n_44)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_12),
.B(n_3),
.Y(n_31)
);

HAxp5_ASAP7_75t_SL g32 ( 
.A(n_20),
.B(n_4),
.CON(n_32),
.SN(n_32)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_33),
.A2(n_43),
.B1(n_5),
.B2(n_9),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_28),
.A2(n_19),
.B1(n_16),
.B2(n_17),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_34),
.A2(n_47),
.B1(n_45),
.B2(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_16),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_44),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_17),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_42),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_21),
.C(n_18),
.Y(n_42)
);

AND2x6_ASAP7_75t_L g43 ( 
.A(n_23),
.B(n_4),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_16),
.Y(n_45)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_45),
.B(n_46),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_17),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_21),
.C(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_50),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_26),
.B(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_27),
.B(n_14),
.Y(n_50)
);

AO32x1_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_14),
.A3(n_21),
.B1(n_8),
.B2(n_9),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_56),
.B1(n_57),
.B2(n_63),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_10),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_39),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_55),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_66),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_40),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_52),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_44),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_44),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_70),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_36),
.C(n_49),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_43),
.C(n_35),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_SL g72 ( 
.A(n_54),
.B(n_10),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_76),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_52),
.B1(n_57),
.B2(n_58),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_62),
.B(n_11),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_75),
.C(n_61),
.Y(n_82)
);

NOR2x1_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_72),
.Y(n_79)
);

OAI31xp33_ASAP7_75t_L g84 ( 
.A1(n_79),
.A2(n_81),
.A3(n_78),
.B(n_69),
.Y(n_84)
);

NOR2x1_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_67),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_75),
.C(n_79),
.Y(n_83)
);

O2A1O1Ixp33_ASAP7_75t_SL g85 ( 
.A1(n_84),
.A2(n_81),
.B(n_78),
.C(n_80),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_83),
.C(n_80),
.Y(n_86)
);


endmodule