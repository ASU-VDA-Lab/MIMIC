module fake_netlist_6_1724_n_1881 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1881);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1881;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1821;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_7),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_168),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_61),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_92),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_130),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_138),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_59),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_3),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_159),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_90),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_153),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_17),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_13),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_43),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_68),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_78),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_88),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g193 ( 
.A(n_58),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_147),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_49),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_56),
.Y(n_197)
);

INVxp33_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_107),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_117),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_165),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_172),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_76),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_40),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_102),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_60),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_47),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_41),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_108),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_152),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_134),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_17),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_1),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_158),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_32),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_35),
.Y(n_216)
);

BUFx2_ASAP7_75t_SL g217 ( 
.A(n_64),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_40),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_66),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_58),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_91),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_25),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_63),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_101),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_120),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_109),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_57),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_7),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_49),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_82),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_62),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_113),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_129),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_29),
.Y(n_234)
);

INVxp33_ASAP7_75t_L g235 ( 
.A(n_116),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_16),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_16),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_166),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_83),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_119),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_139),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_111),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_56),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_41),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_20),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_160),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_94),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_44),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_26),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_65),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_95),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_155),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_106),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_14),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_24),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_47),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_32),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_63),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_87),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_118),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_64),
.Y(n_261)
);

BUFx10_ASAP7_75t_L g262 ( 
.A(n_60),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_2),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_25),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_128),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_142),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_74),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_148),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_93),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_3),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_14),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_37),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_156),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_105),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_137),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_45),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_33),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_70),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_141),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_132),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_44),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_26),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_59),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_135),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_133),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_170),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_86),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_103),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_21),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_37),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_157),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_171),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_4),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_110),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_50),
.Y(n_295)
);

BUFx5_ASAP7_75t_L g296 ( 
.A(n_97),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_174),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_115),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_104),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_89),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_85),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_66),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_84),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_126),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_143),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_50),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_53),
.Y(n_307)
);

BUFx10_ASAP7_75t_L g308 ( 
.A(n_124),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_10),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_151),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_169),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_114),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_77),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_51),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_39),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_52),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_30),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_61),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_80),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_0),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_34),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_127),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_4),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_20),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_73),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_150),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_36),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_33),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_1),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_28),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_167),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_149),
.Y(n_332)
);

BUFx5_ASAP7_75t_L g333 ( 
.A(n_13),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_154),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_98),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_2),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_6),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_55),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_46),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_38),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_72),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_27),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_65),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_54),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_21),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_55),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_161),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_6),
.Y(n_348)
);

NOR2xp67_ASAP7_75t_L g349 ( 
.A(n_181),
.B(n_0),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_193),
.Y(n_350)
);

INVxp33_ASAP7_75t_SL g351 ( 
.A(n_261),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_176),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_193),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_210),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_193),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_211),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_313),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_193),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_193),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_265),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_334),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_302),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_247),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_193),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_193),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_177),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_306),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_214),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_193),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_257),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_333),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_198),
.B(n_5),
.Y(n_372)
);

NOR2xp67_ASAP7_75t_L g373 ( 
.A(n_181),
.B(n_5),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_333),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_221),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_224),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_235),
.B(n_8),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_333),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_312),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_333),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_226),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_232),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_238),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_333),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_333),
.Y(n_385)
);

INVxp33_ASAP7_75t_SL g386 ( 
.A(n_175),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_239),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_240),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_242),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_333),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_246),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_333),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_216),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_251),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_252),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_216),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_257),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_267),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_273),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_185),
.B(n_8),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_279),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_280),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_288),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_294),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_216),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_216),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_185),
.B(n_9),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_201),
.B(n_9),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_R g409 ( 
.A(n_298),
.B(n_122),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_201),
.B(n_10),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_300),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_308),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_301),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_212),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_192),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_216),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_228),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_215),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_218),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_228),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_228),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_228),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_219),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_228),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_179),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_307),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_179),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_220),
.Y(n_428)
);

BUFx10_ASAP7_75t_L g429 ( 
.A(n_259),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_175),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_188),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_259),
.B(n_11),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_182),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_180),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_307),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_222),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_359),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_360),
.B(n_192),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_393),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_360),
.B(n_241),
.Y(n_440)
);

NOR2x1_ASAP7_75t_L g441 ( 
.A(n_360),
.B(n_241),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_372),
.B(n_307),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_393),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_431),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_396),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_377),
.B(n_400),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_396),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_405),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_359),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_415),
.B(n_274),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_392),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_405),
.B(n_274),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_406),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_360),
.B(n_326),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_392),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_406),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_416),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_350),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_350),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_414),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_430),
.Y(n_461)
);

OA21x2_ASAP7_75t_L g462 ( 
.A1(n_353),
.A2(n_213),
.B(n_197),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_416),
.B(n_326),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_353),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_355),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_417),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_417),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_355),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_358),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_358),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_420),
.B(n_307),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_433),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_420),
.B(n_307),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_364),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_364),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_421),
.Y(n_476)
);

AND2x6_ASAP7_75t_L g477 ( 
.A(n_365),
.B(n_265),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_379),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_365),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_412),
.B(n_308),
.Y(n_480)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_429),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_421),
.Y(n_482)
);

AND2x6_ASAP7_75t_L g483 ( 
.A(n_369),
.B(n_265),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_422),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_422),
.B(n_209),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_424),
.B(n_329),
.Y(n_486)
);

AND2x6_ASAP7_75t_L g487 ( 
.A(n_369),
.B(n_265),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_407),
.B(n_329),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_371),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_410),
.B(n_329),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_412),
.B(n_308),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_432),
.B(n_329),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_424),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_371),
.Y(n_494)
);

AND2x6_ASAP7_75t_L g495 ( 
.A(n_374),
.B(n_265),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_426),
.B(n_209),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_354),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_426),
.B(n_284),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_435),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_435),
.B(n_374),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_378),
.B(n_329),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_378),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_380),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_380),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_384),
.Y(n_505)
);

CKINVDCx6p67_ASAP7_75t_R g506 ( 
.A(n_363),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_384),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_385),
.B(n_180),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_385),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_390),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_390),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_429),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_349),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_351),
.A2(n_276),
.B1(n_345),
.B2(n_196),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_446),
.B(n_356),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_437),
.Y(n_516)
);

BUFx10_ASAP7_75t_L g517 ( 
.A(n_497),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_450),
.B(n_418),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_455),
.Y(n_519)
);

NAND2xp33_ASAP7_75t_L g520 ( 
.A(n_488),
.B(n_266),
.Y(n_520)
);

CKINVDCx16_ASAP7_75t_R g521 ( 
.A(n_444),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_450),
.B(n_419),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_512),
.B(n_368),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_512),
.B(n_375),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_462),
.Y(n_525)
);

OR2x6_ASAP7_75t_L g526 ( 
.A(n_460),
.B(n_217),
.Y(n_526)
);

INVx1_ASAP7_75t_SL g527 ( 
.A(n_444),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_446),
.A2(n_408),
.B1(n_367),
.B2(n_362),
.Y(n_528)
);

BUFx6f_ASAP7_75t_SL g529 ( 
.A(n_481),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_462),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_450),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_437),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_438),
.B(n_349),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_462),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_470),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_461),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_437),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_455),
.Y(n_538)
);

CKINVDCx6p67_ASAP7_75t_R g539 ( 
.A(n_506),
.Y(n_539)
);

AND2x6_ASAP7_75t_L g540 ( 
.A(n_512),
.B(n_284),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_478),
.A2(n_382),
.B1(n_388),
.B2(n_381),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_462),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_437),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_462),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_478),
.B(n_376),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_512),
.B(n_383),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_481),
.B(n_387),
.Y(n_547)
);

AND2x6_ASAP7_75t_L g548 ( 
.A(n_512),
.B(n_291),
.Y(n_548)
);

OAI21xp33_ASAP7_75t_L g549 ( 
.A1(n_442),
.A2(n_386),
.B(n_423),
.Y(n_549)
);

BUFx4f_ASAP7_75t_L g550 ( 
.A(n_462),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_481),
.B(n_389),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_455),
.Y(n_552)
);

AND2x2_ASAP7_75t_SL g553 ( 
.A(n_442),
.B(n_291),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_481),
.B(n_391),
.Y(n_554)
);

CKINVDCx6p67_ASAP7_75t_R g555 ( 
.A(n_506),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_481),
.B(n_394),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_455),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_480),
.A2(n_401),
.B1(n_411),
.B2(n_395),
.Y(n_558)
);

OAI221xp5_ASAP7_75t_L g559 ( 
.A1(n_488),
.A2(n_373),
.B1(n_213),
.B2(n_264),
.C(n_263),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_460),
.B(n_398),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_471),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_437),
.Y(n_562)
);

OR2x6_ASAP7_75t_L g563 ( 
.A(n_460),
.B(n_231),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_471),
.Y(n_564)
);

BUFx10_ASAP7_75t_L g565 ( 
.A(n_461),
.Y(n_565)
);

NOR3xp33_ASAP7_75t_L g566 ( 
.A(n_514),
.B(n_366),
.C(n_370),
.Y(n_566)
);

CKINVDCx16_ASAP7_75t_R g567 ( 
.A(n_472),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_472),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_471),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_459),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_506),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_513),
.B(n_428),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_473),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_473),
.Y(n_574)
);

INVx5_ASAP7_75t_L g575 ( 
.A(n_477),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_508),
.B(n_399),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_459),
.Y(n_577)
);

OR2x2_ASAP7_75t_L g578 ( 
.A(n_508),
.B(n_366),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_480),
.B(n_402),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_490),
.B(n_403),
.Y(n_580)
);

AND2x6_ASAP7_75t_L g581 ( 
.A(n_438),
.B(n_331),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_473),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_486),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_486),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_459),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_490),
.B(n_436),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_486),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_492),
.B(n_503),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_503),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_491),
.B(n_404),
.Y(n_590)
);

BUFx4f_ASAP7_75t_L g591 ( 
.A(n_470),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_504),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_459),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_504),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_492),
.B(n_429),
.Y(n_595)
);

BUFx10_ASAP7_75t_L g596 ( 
.A(n_463),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_500),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_491),
.B(n_413),
.Y(n_598)
);

BUFx8_ASAP7_75t_SL g599 ( 
.A(n_514),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_500),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_513),
.B(n_429),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_438),
.B(n_178),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_464),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_464),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_452),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_500),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_464),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_500),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_464),
.Y(n_609)
);

OR2x6_ASAP7_75t_L g610 ( 
.A(n_463),
.B(n_231),
.Y(n_610)
);

INVx4_ASAP7_75t_L g611 ( 
.A(n_470),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_468),
.Y(n_612)
);

NAND3xp33_ASAP7_75t_L g613 ( 
.A(n_452),
.B(n_397),
.C(n_229),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_465),
.B(n_425),
.Y(n_614)
);

NAND3xp33_ASAP7_75t_L g615 ( 
.A(n_452),
.B(n_234),
.C(n_227),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_438),
.B(n_299),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_500),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_438),
.B(n_440),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_440),
.B(n_331),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_463),
.A2(n_373),
.B1(n_248),
.B2(n_278),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_463),
.A2(n_434),
.B1(n_427),
.B2(n_244),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_458),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_470),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_458),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_463),
.B(n_409),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_437),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_468),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_468),
.Y(n_628)
);

NAND2xp33_ASAP7_75t_L g629 ( 
.A(n_477),
.B(n_266),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_437),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_437),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_440),
.B(n_183),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_440),
.B(n_184),
.Y(n_633)
);

NAND3xp33_ASAP7_75t_SL g634 ( 
.A(n_501),
.B(n_324),
.C(n_207),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_468),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_SL g636 ( 
.A(n_441),
.B(n_352),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_440),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_470),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_458),
.Y(n_639)
);

INVx4_ASAP7_75t_L g640 ( 
.A(n_470),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_465),
.B(n_361),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_489),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_465),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_454),
.B(n_485),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_489),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_469),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_454),
.B(n_190),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_489),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_489),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_454),
.B(n_183),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_469),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_454),
.B(n_465),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_469),
.Y(n_653)
);

BUFx4f_ASAP7_75t_L g654 ( 
.A(n_470),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_465),
.Y(n_655)
);

AND2x6_ASAP7_75t_L g656 ( 
.A(n_454),
.B(n_266),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_470),
.Y(n_657)
);

NOR2x1p5_ASAP7_75t_L g658 ( 
.A(n_501),
.B(n_182),
.Y(n_658)
);

NAND2xp33_ASAP7_75t_L g659 ( 
.A(n_477),
.B(n_266),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_474),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_449),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_474),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_449),
.Y(n_663)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_494),
.B(n_337),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_494),
.B(n_357),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_441),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_474),
.Y(n_667)
);

NOR2xp67_ASAP7_75t_SL g668 ( 
.A(n_575),
.B(n_266),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_515),
.B(n_494),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_586),
.B(n_494),
.Y(n_670)
);

CKINVDCx11_ASAP7_75t_R g671 ( 
.A(n_517),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_553),
.B(n_494),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_553),
.B(n_474),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_531),
.B(n_191),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_531),
.B(n_191),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_580),
.B(n_194),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_550),
.B(n_474),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_550),
.B(n_474),
.Y(n_678)
);

BUFx8_ASAP7_75t_L g679 ( 
.A(n_536),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_605),
.B(n_474),
.Y(n_680)
);

NOR2xp67_ASAP7_75t_L g681 ( 
.A(n_541),
.B(n_439),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_550),
.B(n_600),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_595),
.B(n_474),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_644),
.Y(n_684)
);

CKINVDCx20_ASAP7_75t_R g685 ( 
.A(n_521),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_525),
.A2(n_289),
.B1(n_283),
.B2(n_272),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_588),
.B(n_475),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_661),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_576),
.B(n_475),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_644),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_589),
.B(n_475),
.Y(n_691)
);

NOR3xp33_ASAP7_75t_L g692 ( 
.A(n_621),
.B(n_249),
.C(n_236),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_578),
.B(n_194),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_600),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_569),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_606),
.Y(n_696)
);

HB1xp67_ASAP7_75t_L g697 ( 
.A(n_527),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_578),
.B(n_199),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_606),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_589),
.B(n_475),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_592),
.B(n_594),
.Y(n_701)
);

AO21x2_ASAP7_75t_L g702 ( 
.A1(n_525),
.A2(n_200),
.B(n_195),
.Y(n_702)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_536),
.B(n_187),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_592),
.B(n_475),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_530),
.A2(n_254),
.B1(n_208),
.B2(n_206),
.Y(n_705)
);

BUFx5_ASAP7_75t_L g706 ( 
.A(n_530),
.Y(n_706)
);

NOR2xp67_ASAP7_75t_L g707 ( 
.A(n_579),
.B(n_439),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_569),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_608),
.B(n_475),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_549),
.B(n_199),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_596),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_608),
.B(n_617),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_617),
.B(n_475),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_594),
.B(n_573),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_597),
.B(n_475),
.Y(n_715)
);

INVx8_ASAP7_75t_L g716 ( 
.A(n_526),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_663),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_637),
.B(n_505),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_573),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_545),
.B(n_203),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_518),
.A2(n_322),
.B1(n_325),
.B2(n_332),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_637),
.B(n_505),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_574),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_518),
.B(n_257),
.Y(n_724)
);

INVxp67_ASAP7_75t_L g725 ( 
.A(n_568),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_596),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_522),
.B(n_203),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_519),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_582),
.Y(n_729)
);

A2O1A1Ixp33_ASAP7_75t_SL g730 ( 
.A1(n_534),
.A2(n_275),
.B(n_319),
.C(n_297),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_522),
.B(n_572),
.Y(n_731)
);

BUFx12f_ASAP7_75t_L g732 ( 
.A(n_517),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_582),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_572),
.B(n_268),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_583),
.Y(n_735)
);

NAND2x1_ASAP7_75t_L g736 ( 
.A(n_534),
.B(n_477),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_618),
.B(n_583),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_584),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_584),
.B(n_505),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_587),
.B(n_505),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_587),
.B(n_505),
.Y(n_741)
);

INVxp67_ASAP7_75t_SL g742 ( 
.A(n_542),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_542),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_664),
.B(n_268),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_666),
.B(n_505),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_596),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_666),
.B(n_505),
.Y(n_747)
);

OR2x2_ASAP7_75t_L g748 ( 
.A(n_568),
.B(n_567),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_519),
.Y(n_749)
);

BUFx10_ASAP7_75t_L g750 ( 
.A(n_658),
.Y(n_750)
);

OR2x2_ASAP7_75t_L g751 ( 
.A(n_664),
.B(n_187),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_601),
.B(n_262),
.Y(n_752)
);

NAND3xp33_ASAP7_75t_L g753 ( 
.A(n_528),
.B(n_255),
.C(n_250),
.Y(n_753)
);

OAI21xp33_ASAP7_75t_L g754 ( 
.A1(n_601),
.A2(n_204),
.B(n_186),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_523),
.A2(n_335),
.B1(n_292),
.B2(n_287),
.Y(n_755)
);

AND2x6_ASAP7_75t_L g756 ( 
.A(n_544),
.B(n_205),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_614),
.B(n_303),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_561),
.B(n_505),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_564),
.B(n_507),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_547),
.B(n_507),
.Y(n_760)
);

OAI22xp33_ASAP7_75t_L g761 ( 
.A1(n_559),
.A2(n_321),
.B1(n_245),
.B2(n_243),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_634),
.B(n_303),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_554),
.B(n_507),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_524),
.B(n_546),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_652),
.B(n_507),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_619),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_544),
.B(n_507),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_565),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_633),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_L g770 ( 
.A1(n_551),
.A2(n_285),
.B1(n_286),
.B2(n_269),
.Y(n_770)
);

O2A1O1Ixp5_ASAP7_75t_L g771 ( 
.A1(n_647),
.A2(n_485),
.B(n_496),
.C(n_498),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_643),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_533),
.B(n_507),
.Y(n_773)
);

OR2x6_ASAP7_75t_L g774 ( 
.A(n_526),
.B(n_223),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_538),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_655),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_538),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_533),
.B(n_507),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_533),
.B(n_507),
.Y(n_779)
);

INVx1_ASAP7_75t_SL g780 ( 
.A(n_565),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_556),
.B(n_510),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_602),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_616),
.B(n_510),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_516),
.B(n_510),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_610),
.B(n_225),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_552),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_622),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_613),
.B(n_304),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_615),
.B(n_304),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_516),
.B(n_510),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_516),
.B(n_510),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_532),
.B(n_510),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_581),
.A2(n_346),
.B1(n_323),
.B2(n_330),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_L g794 ( 
.A1(n_641),
.A2(n_260),
.B1(n_253),
.B2(n_233),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_532),
.B(n_510),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_532),
.B(n_510),
.Y(n_796)
);

BUFx6f_ASAP7_75t_SL g797 ( 
.A(n_517),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_543),
.B(n_511),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_581),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_552),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_557),
.Y(n_801)
);

NAND2xp33_ASAP7_75t_L g802 ( 
.A(n_581),
.B(n_202),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_665),
.B(n_511),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_565),
.B(n_262),
.Y(n_804)
);

NAND3xp33_ASAP7_75t_L g805 ( 
.A(n_620),
.B(n_271),
.C(n_295),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_543),
.B(n_511),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_563),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_563),
.B(n_262),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_543),
.B(n_511),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_563),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_563),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_562),
.B(n_511),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_562),
.B(n_626),
.Y(n_813)
);

BUFx6f_ASAP7_75t_SL g814 ( 
.A(n_526),
.Y(n_814)
);

NOR3xp33_ASAP7_75t_L g815 ( 
.A(n_590),
.B(n_277),
.C(n_256),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_636),
.B(n_511),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_632),
.A2(n_310),
.B1(n_341),
.B2(n_332),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_557),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_570),
.Y(n_819)
);

NOR3xp33_ASAP7_75t_L g820 ( 
.A(n_598),
.B(n_270),
.C(n_281),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_562),
.B(n_511),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_570),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_626),
.B(n_511),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_575),
.B(n_479),
.Y(n_824)
);

INVxp33_ASAP7_75t_L g825 ( 
.A(n_566),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_624),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_577),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_581),
.Y(n_828)
);

OR2x6_ASAP7_75t_L g829 ( 
.A(n_526),
.B(n_237),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_626),
.B(n_509),
.Y(n_830)
);

BUFx5_ASAP7_75t_L g831 ( 
.A(n_581),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_631),
.B(n_509),
.Y(n_832)
);

OR2x2_ASAP7_75t_L g833 ( 
.A(n_560),
.B(n_189),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_631),
.B(n_509),
.Y(n_834)
);

NOR3xp33_ASAP7_75t_L g835 ( 
.A(n_731),
.B(n_558),
.C(n_650),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_731),
.A2(n_625),
.B1(n_581),
.B2(n_610),
.Y(n_836)
);

O2A1O1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_737),
.A2(n_672),
.B(n_712),
.C(n_794),
.Y(n_837)
);

A2O1A1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_720),
.A2(n_520),
.B(n_230),
.C(n_631),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_720),
.B(n_610),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_677),
.A2(n_654),
.B(n_591),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_764),
.A2(n_610),
.B1(n_540),
.B2(n_548),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_673),
.A2(n_529),
.B1(n_591),
.B2(n_654),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_782),
.A2(n_548),
.B1(n_540),
.B2(n_529),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_SL g844 ( 
.A(n_732),
.B(n_797),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_676),
.B(n_540),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_677),
.A2(n_654),
.B(n_591),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_SL g847 ( 
.A(n_797),
.B(n_571),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_678),
.A2(n_611),
.B(n_535),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_697),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_676),
.B(n_540),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_695),
.B(n_540),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_708),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_711),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_695),
.Y(n_854)
);

BUFx12f_ASAP7_75t_L g855 ( 
.A(n_671),
.Y(n_855)
);

CKINVDCx20_ASAP7_75t_R g856 ( 
.A(n_685),
.Y(n_856)
);

BUFx2_ASAP7_75t_L g857 ( 
.A(n_748),
.Y(n_857)
);

INVxp67_ASAP7_75t_SL g858 ( 
.A(n_743),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_707),
.B(n_575),
.Y(n_859)
);

BUFx8_ASAP7_75t_L g860 ( 
.A(n_814),
.Y(n_860)
);

NOR3xp33_ASAP7_75t_L g861 ( 
.A(n_757),
.B(n_310),
.C(n_305),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_725),
.B(n_539),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_678),
.A2(n_611),
.B(n_535),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_684),
.B(n_336),
.Y(n_864)
);

OAI21xp33_ASAP7_75t_L g865 ( 
.A1(n_757),
.A2(n_258),
.B(n_189),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_742),
.B(n_540),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_711),
.B(n_575),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_690),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_773),
.A2(n_611),
.B(n_535),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_727),
.B(n_539),
.Y(n_870)
);

O2A1O1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_737),
.A2(n_520),
.B(n_639),
.C(n_653),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_711),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_669),
.A2(n_529),
.B1(n_651),
.B2(n_646),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_727),
.B(n_693),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_778),
.A2(n_640),
.B(n_623),
.Y(n_875)
);

O2A1O1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_712),
.A2(n_639),
.B(n_646),
.C(n_651),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_711),
.B(n_575),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_769),
.B(n_548),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_719),
.B(n_548),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_679),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_723),
.B(n_548),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_734),
.B(n_305),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_779),
.A2(n_640),
.B(n_623),
.Y(n_883)
);

O2A1O1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_714),
.A2(n_733),
.B(n_735),
.C(n_729),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_779),
.A2(n_640),
.B(n_623),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_SL g886 ( 
.A(n_780),
.B(n_555),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_783),
.A2(n_630),
.B(n_537),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_689),
.A2(n_630),
.B(n_537),
.Y(n_888)
);

A2O1A1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_710),
.A2(n_653),
.B(n_660),
.C(n_638),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_734),
.B(n_311),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_814),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_706),
.B(n_537),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_687),
.A2(n_630),
.B(n_537),
.Y(n_893)
);

OAI22xp5_ASAP7_75t_L g894 ( 
.A1(n_743),
.A2(n_667),
.B1(n_660),
.B2(n_657),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_745),
.A2(n_630),
.B(n_537),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_738),
.B(n_548),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_706),
.B(n_638),
.Y(n_897)
);

O2A1O1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_682),
.A2(n_701),
.B(n_816),
.C(n_694),
.Y(n_898)
);

INVx5_ASAP7_75t_L g899 ( 
.A(n_799),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_747),
.A2(n_630),
.B(n_662),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_724),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_744),
.B(n_311),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_781),
.A2(n_662),
.B(n_667),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_781),
.A2(n_662),
.B(n_667),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_760),
.A2(n_662),
.B(n_660),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_693),
.B(n_555),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_799),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_744),
.B(n_322),
.Y(n_908)
);

AOI21x1_ASAP7_75t_L g909 ( 
.A1(n_767),
.A2(n_593),
.B(n_604),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_816),
.A2(n_656),
.B1(n_657),
.B2(n_638),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_696),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_699),
.A2(n_657),
.B1(n_325),
.B2(n_341),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_736),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_706),
.B(n_577),
.Y(n_914)
);

O2A1O1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_682),
.A2(n_629),
.B(n_659),
.C(n_593),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_763),
.A2(n_662),
.B(n_612),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_767),
.A2(n_604),
.B(n_585),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_680),
.A2(n_612),
.B(n_585),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_765),
.A2(n_627),
.B(n_603),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_698),
.B(n_603),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_787),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_765),
.A2(n_627),
.B(n_607),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_710),
.A2(n_670),
.B(n_789),
.C(n_788),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_706),
.B(n_607),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_718),
.A2(n_628),
.B(n_609),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_819),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_706),
.B(n_609),
.Y(n_927)
);

OAI21xp33_ASAP7_75t_L g928 ( 
.A1(n_698),
.A2(n_258),
.B(n_309),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_752),
.B(n_309),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_679),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_766),
.B(n_628),
.Y(n_931)
);

O2A1O1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_770),
.A2(n_659),
.B(n_629),
.C(n_649),
.Y(n_932)
);

AOI21x1_ASAP7_75t_L g933 ( 
.A1(n_718),
.A2(n_649),
.B(n_648),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_825),
.B(n_635),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_722),
.A2(n_648),
.B(n_645),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_751),
.B(n_635),
.Y(n_936)
);

NOR2xp67_ASAP7_75t_L g937 ( 
.A(n_768),
.B(n_347),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_804),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_771),
.A2(n_642),
.B(n_479),
.Y(n_939)
);

A2O1A1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_670),
.A2(n_496),
.B(n_485),
.C(n_498),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_683),
.A2(n_502),
.B(n_479),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_803),
.A2(n_502),
.B(n_451),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_803),
.A2(n_502),
.B(n_451),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_810),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_807),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_813),
.A2(n_451),
.B(n_449),
.Y(n_946)
);

O2A1O1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_755),
.A2(n_754),
.B(n_740),
.C(n_761),
.Y(n_947)
);

AO21x1_ASAP7_75t_L g948 ( 
.A1(n_762),
.A2(n_498),
.B(n_496),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_739),
.A2(n_451),
.B(n_449),
.Y(n_949)
);

O2A1O1Ixp33_ASAP7_75t_SL g950 ( 
.A1(n_730),
.A2(n_348),
.B(n_342),
.C(n_338),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_703),
.B(n_314),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_789),
.B(n_347),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_674),
.B(n_656),
.Y(n_953)
);

O2A1O1Ixp33_ASAP7_75t_SL g954 ( 
.A1(n_730),
.A2(n_339),
.B(n_499),
.C(n_457),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_674),
.B(n_656),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_826),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_L g957 ( 
.A1(n_686),
.A2(n_485),
.B1(n_496),
.B2(n_498),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_741),
.A2(n_451),
.B(n_449),
.Y(n_958)
);

INVx5_ASAP7_75t_L g959 ( 
.A(n_799),
.Y(n_959)
);

AOI22xp5_ASAP7_75t_L g960 ( 
.A1(n_788),
.A2(n_656),
.B1(n_485),
.B2(n_496),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_758),
.A2(n_498),
.B(n_499),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_750),
.Y(n_962)
);

NAND3xp33_ASAP7_75t_L g963 ( 
.A(n_762),
.B(n_293),
.C(n_290),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_822),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_726),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_772),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_675),
.B(n_202),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_759),
.A2(n_445),
.B(n_443),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_833),
.B(n_282),
.Y(n_969)
);

AOI22xp5_ASAP7_75t_L g970 ( 
.A1(n_681),
.A2(n_656),
.B1(n_448),
.B2(n_447),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_753),
.B(n_314),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_686),
.B(n_656),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_705),
.B(n_445),
.Y(n_973)
);

NOR3xp33_ASAP7_75t_L g974 ( 
.A(n_692),
.B(n_315),
.C(n_316),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_822),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_831),
.B(n_202),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_721),
.B(n_315),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_784),
.A2(n_453),
.B(n_447),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_790),
.A2(n_456),
.B(n_448),
.Y(n_979)
);

AND2x2_ASAP7_75t_SL g980 ( 
.A(n_705),
.B(n_599),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_791),
.A2(n_456),
.B(n_453),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_R g982 ( 
.A(n_811),
.B(n_316),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_726),
.B(n_457),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_792),
.A2(n_466),
.B(n_467),
.Y(n_984)
);

INVxp67_ASAP7_75t_L g985 ( 
.A(n_808),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_795),
.A2(n_467),
.B(n_476),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_750),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_709),
.A2(n_477),
.B(n_495),
.Y(n_988)
);

AOI33xp33_ASAP7_75t_L g989 ( 
.A1(n_761),
.A2(n_599),
.A3(n_343),
.B1(n_340),
.B2(n_318),
.B3(n_320),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_688),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_799),
.Y(n_991)
);

OAI21xp5_ASAP7_75t_L g992 ( 
.A1(n_709),
.A2(n_495),
.B(n_477),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_796),
.A2(n_476),
.B(n_493),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_SL g994 ( 
.A1(n_824),
.A2(n_482),
.B(n_484),
.C(n_202),
.Y(n_994)
);

BUFx12f_ASAP7_75t_L g995 ( 
.A(n_774),
.Y(n_995)
);

A2O1A1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_776),
.A2(n_482),
.B(n_484),
.C(n_317),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_828),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_746),
.B(n_495),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_774),
.B(n_829),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_746),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_798),
.A2(n_495),
.B(n_487),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_785),
.B(n_202),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_828),
.A2(n_328),
.B1(n_317),
.B2(n_318),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_774),
.Y(n_1004)
);

NOR2x1_ASAP7_75t_L g1005 ( 
.A(n_829),
.B(n_320),
.Y(n_1005)
);

AOI21x1_ASAP7_75t_L g1006 ( 
.A1(n_713),
.A2(n_495),
.B(n_487),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_691),
.A2(n_343),
.B(n_327),
.C(n_328),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_700),
.B(n_495),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_704),
.B(n_495),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_702),
.B(n_827),
.Y(n_1010)
);

INVx5_ASAP7_75t_L g1011 ( 
.A(n_828),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_702),
.B(n_495),
.Y(n_1012)
);

AOI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_756),
.A2(n_793),
.B1(n_828),
.B2(n_713),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_728),
.B(n_495),
.Y(n_1014)
);

AOI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_785),
.A2(n_495),
.B1(n_487),
.B2(n_483),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_749),
.B(n_775),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_806),
.A2(n_487),
.B(n_483),
.Y(n_1017)
);

BUFx12f_ASAP7_75t_L g1018 ( 
.A(n_860),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_923),
.A2(n_802),
.B(n_832),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_874),
.A2(n_820),
.B(n_815),
.C(n_817),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_852),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_853),
.Y(n_1022)
);

NAND3xp33_ASAP7_75t_SL g1023 ( 
.A(n_874),
.B(n_793),
.C(n_327),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_858),
.A2(n_834),
.B(n_830),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_856),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_936),
.B(n_756),
.Y(n_1026)
);

O2A1O1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_996),
.A2(n_715),
.B(n_777),
.C(n_786),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_SL g1028 ( 
.A1(n_878),
.A2(n_809),
.B(n_823),
.C(n_821),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_858),
.A2(n_812),
.B(n_717),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_845),
.A2(n_800),
.B(n_818),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_980),
.B(n_831),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_L g1032 ( 
.A1(n_909),
.A2(n_801),
.B(n_824),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_868),
.Y(n_1033)
);

INVx4_ASAP7_75t_L g1034 ( 
.A(n_853),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_850),
.A2(n_831),
.B(n_716),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_853),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_929),
.B(n_829),
.Y(n_1037)
);

OAI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_898),
.A2(n_756),
.B(n_805),
.Y(n_1038)
);

O2A1O1Ixp5_ASAP7_75t_L g1039 ( 
.A1(n_967),
.A2(n_668),
.B(n_756),
.C(n_831),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_888),
.A2(n_831),
.B(n_716),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_853),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_839),
.A2(n_756),
.B1(n_340),
.B2(n_344),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_866),
.A2(n_487),
.B(n_483),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_936),
.B(n_344),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_884),
.A2(n_296),
.B(n_202),
.C(n_15),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_840),
.A2(n_487),
.B(n_483),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_839),
.A2(n_296),
.B(n_202),
.C(n_15),
.Y(n_1047)
);

NOR3xp33_ASAP7_75t_L g1048 ( 
.A(n_974),
.B(n_870),
.C(n_969),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_980),
.B(n_296),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_846),
.A2(n_487),
.B(n_483),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_872),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_835),
.A2(n_296),
.B(n_12),
.C(n_18),
.Y(n_1052)
);

INVx2_ASAP7_75t_SL g1053 ( 
.A(n_849),
.Y(n_1053)
);

BUFx3_ASAP7_75t_L g1054 ( 
.A(n_857),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_951),
.B(n_296),
.Y(n_1055)
);

INVx1_ASAP7_75t_SL g1056 ( 
.A(n_849),
.Y(n_1056)
);

OAI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_901),
.A2(n_11),
.B1(n_12),
.B2(n_18),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_872),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_944),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_870),
.B(n_19),
.Y(n_1060)
);

O2A1O1Ixp33_ASAP7_75t_SL g1061 ( 
.A1(n_976),
.A2(n_296),
.B(n_164),
.C(n_163),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_872),
.Y(n_1062)
);

XOR2xp5_ASAP7_75t_L g1063 ( 
.A(n_891),
.B(n_146),
.Y(n_1063)
);

O2A1O1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_835),
.A2(n_296),
.B(n_22),
.C(n_23),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_868),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_934),
.B(n_487),
.Y(n_1066)
);

BUFx2_ASAP7_75t_L g1067 ( 
.A(n_944),
.Y(n_1067)
);

OA21x2_ASAP7_75t_L g1068 ( 
.A1(n_1010),
.A2(n_487),
.B(n_483),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_893),
.A2(n_940),
.B(n_887),
.Y(n_1069)
);

O2A1O1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_947),
.A2(n_296),
.B(n_22),
.C(n_23),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_1004),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_854),
.B(n_934),
.Y(n_1072)
);

O2A1O1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_1007),
.A2(n_19),
.B(n_24),
.C(n_27),
.Y(n_1073)
);

INVx4_ASAP7_75t_L g1074 ( 
.A(n_872),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_854),
.B(n_487),
.Y(n_1075)
);

NAND3xp33_ASAP7_75t_SL g1076 ( 
.A(n_861),
.B(n_28),
.C(n_29),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_1004),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_911),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_921),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_836),
.A2(n_121),
.B1(n_75),
.B2(n_145),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_889),
.A2(n_483),
.B(n_477),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_926),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_956),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_920),
.B(n_30),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_966),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_1013),
.A2(n_144),
.B1(n_140),
.B2(n_136),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_964),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_975),
.Y(n_1088)
);

BUFx8_ASAP7_75t_L g1089 ( 
.A(n_880),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_1013),
.A2(n_131),
.B1(n_123),
.B2(n_112),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_920),
.B(n_31),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_969),
.B(n_906),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_906),
.B(n_882),
.Y(n_1093)
);

INVx5_ASAP7_75t_L g1094 ( 
.A(n_907),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_977),
.B(n_31),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_905),
.A2(n_100),
.B(n_99),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_892),
.A2(n_955),
.B(n_953),
.Y(n_1097)
);

INVx3_ASAP7_75t_SL g1098 ( 
.A(n_930),
.Y(n_1098)
);

CKINVDCx8_ASAP7_75t_R g1099 ( 
.A(n_864),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_945),
.B(n_96),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_938),
.B(n_81),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_861),
.B(n_79),
.Y(n_1102)
);

HB1xp67_ASAP7_75t_L g1103 ( 
.A(n_945),
.Y(n_1103)
);

BUFx3_ASAP7_75t_L g1104 ( 
.A(n_987),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_990),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_974),
.A2(n_971),
.B1(n_977),
.B2(n_952),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_862),
.B(n_34),
.Y(n_1107)
);

AOI22xp33_ASAP7_75t_L g1108 ( 
.A1(n_971),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_890),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_1109)
);

AND2x4_ASAP7_75t_L g1110 ( 
.A(n_985),
.B(n_71),
.Y(n_1110)
);

NAND2xp33_ASAP7_75t_SL g1111 ( 
.A(n_907),
.B(n_42),
.Y(n_1111)
);

INVx2_ASAP7_75t_SL g1112 ( 
.A(n_864),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_865),
.B(n_928),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_999),
.B(n_45),
.Y(n_1114)
);

CKINVDCx20_ASAP7_75t_R g1115 ( 
.A(n_860),
.Y(n_1115)
);

O2A1O1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_973),
.A2(n_46),
.B(n_48),
.C(n_51),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_841),
.A2(n_48),
.B(n_52),
.C(n_53),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_892),
.A2(n_54),
.B(n_57),
.Y(n_1118)
);

NAND3xp33_ASAP7_75t_L g1119 ( 
.A(n_902),
.B(n_62),
.C(n_67),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_907),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_907),
.Y(n_1121)
);

INVx1_ASAP7_75t_SL g1122 ( 
.A(n_982),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_908),
.B(n_67),
.Y(n_1123)
);

INVx11_ASAP7_75t_L g1124 ( 
.A(n_995),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_931),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_899),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_1126)
);

BUFx4f_ASAP7_75t_L g1127 ( 
.A(n_855),
.Y(n_1127)
);

OR2x2_ASAP7_75t_L g1128 ( 
.A(n_1003),
.B(n_69),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_965),
.B(n_1000),
.Y(n_1129)
);

AOI22xp5_ASAP7_75t_SL g1130 ( 
.A1(n_962),
.A2(n_989),
.B1(n_1000),
.B2(n_965),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_963),
.B(n_899),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_915),
.A2(n_896),
.B(n_879),
.C(n_881),
.Y(n_1132)
);

NOR3xp33_ASAP7_75t_SL g1133 ( 
.A(n_1002),
.B(n_912),
.C(n_976),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_R g1134 ( 
.A(n_847),
.B(n_886),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_983),
.B(n_914),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_899),
.A2(n_959),
.B1(n_1011),
.B2(n_851),
.Y(n_1136)
);

BUFx8_ASAP7_75t_L g1137 ( 
.A(n_991),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1005),
.B(n_937),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_991),
.Y(n_1139)
);

O2A1O1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_838),
.A2(n_994),
.B(n_950),
.C(n_871),
.Y(n_1140)
);

OR2x6_ASAP7_75t_L g1141 ( 
.A(n_991),
.B(n_997),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_899),
.A2(n_1011),
.B1(n_959),
.B2(n_991),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_972),
.A2(n_960),
.B(n_876),
.C(n_843),
.Y(n_1143)
);

NOR2xp67_ASAP7_75t_L g1144 ( 
.A(n_1015),
.B(n_970),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_SL g1145 ( 
.A(n_844),
.B(n_959),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_959),
.B(n_1011),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1011),
.A2(n_997),
.B1(n_913),
.B2(n_842),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_R g1148 ( 
.A(n_997),
.B(n_913),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_982),
.B(n_1016),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_916),
.A2(n_927),
.B(n_924),
.Y(n_1150)
);

INVx4_ASAP7_75t_L g1151 ( 
.A(n_997),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_933),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_897),
.B(n_957),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_918),
.B(n_961),
.Y(n_1154)
);

INVxp67_ASAP7_75t_SL g1155 ( 
.A(n_894),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1006),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1014),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_968),
.B(n_948),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_988),
.Y(n_1159)
);

O2A1O1Ixp5_ASAP7_75t_SL g1160 ( 
.A1(n_873),
.A2(n_939),
.B(n_1012),
.C(n_917),
.Y(n_1160)
);

INVx5_ASAP7_75t_L g1161 ( 
.A(n_954),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_848),
.A2(n_863),
.B(n_869),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_978),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_979),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_875),
.A2(n_895),
.B(n_900),
.Y(n_1165)
);

OAI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_910),
.A2(n_885),
.B1(n_883),
.B2(n_998),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1008),
.Y(n_1167)
);

AND2x6_ASAP7_75t_SL g1168 ( 
.A(n_1009),
.B(n_932),
.Y(n_1168)
);

BUFx2_ASAP7_75t_L g1169 ( 
.A(n_1054),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1030),
.A2(n_903),
.B(n_904),
.Y(n_1170)
);

AO21x2_ASAP7_75t_L g1171 ( 
.A1(n_1162),
.A2(n_941),
.B(n_942),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1092),
.B(n_949),
.Y(n_1172)
);

AOI31xp67_ASAP7_75t_L g1173 ( 
.A1(n_1158),
.A2(n_859),
.A3(n_867),
.B(n_877),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_L g1174 ( 
.A(n_1095),
.B(n_981),
.C(n_993),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1030),
.A2(n_919),
.B(n_922),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1160),
.A2(n_943),
.B(n_958),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1106),
.A2(n_925),
.B1(n_935),
.B2(n_992),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1154),
.A2(n_946),
.B(n_984),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1093),
.A2(n_986),
.B1(n_1017),
.B2(n_1001),
.Y(n_1179)
);

AO31x2_ASAP7_75t_L g1180 ( 
.A1(n_1143),
.A2(n_1069),
.A3(n_1166),
.B(n_1162),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1153),
.A2(n_1069),
.B(n_1019),
.Y(n_1181)
);

AOI221x1_ASAP7_75t_L g1182 ( 
.A1(n_1048),
.A2(n_1060),
.B1(n_1047),
.B2(n_1117),
.C(n_1076),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1097),
.A2(n_1019),
.B(n_1132),
.Y(n_1183)
);

AO32x2_ASAP7_75t_L g1184 ( 
.A1(n_1042),
.A2(n_1126),
.A3(n_1090),
.B1(n_1086),
.B2(n_1080),
.Y(n_1184)
);

AOI221xp5_ASAP7_75t_SL g1185 ( 
.A1(n_1070),
.A2(n_1052),
.B1(n_1064),
.B2(n_1108),
.C(n_1073),
.Y(n_1185)
);

BUFx12f_ASAP7_75t_L g1186 ( 
.A(n_1018),
.Y(n_1186)
);

AO21x1_ASAP7_75t_L g1187 ( 
.A1(n_1070),
.A2(n_1048),
.B(n_1045),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1135),
.A2(n_1150),
.B(n_1165),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_SL g1189 ( 
.A1(n_1109),
.A2(n_1119),
.B1(n_1128),
.B2(n_1115),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1020),
.A2(n_1113),
.B(n_1138),
.C(n_1038),
.Y(n_1190)
);

CKINVDCx20_ASAP7_75t_R g1191 ( 
.A(n_1025),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1165),
.A2(n_1032),
.B(n_1040),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1040),
.A2(n_1150),
.B(n_1035),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1084),
.A2(n_1091),
.B(n_1130),
.C(n_1133),
.Y(n_1194)
);

INVx1_ASAP7_75t_SL g1195 ( 
.A(n_1056),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1078),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1026),
.A2(n_1024),
.B(n_1142),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1125),
.B(n_1044),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1079),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1072),
.B(n_1149),
.Y(n_1200)
);

OA21x2_ASAP7_75t_L g1201 ( 
.A1(n_1152),
.A2(n_1039),
.B(n_1029),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1039),
.A2(n_1164),
.B(n_1163),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1053),
.Y(n_1203)
);

NAND3xp33_ASAP7_75t_L g1204 ( 
.A(n_1052),
.B(n_1064),
.C(n_1045),
.Y(n_1204)
);

NOR2xp67_ASAP7_75t_L g1205 ( 
.A(n_1094),
.B(n_1034),
.Y(n_1205)
);

AO31x2_ASAP7_75t_L g1206 ( 
.A1(n_1147),
.A2(n_1096),
.A3(n_1050),
.B(n_1046),
.Y(n_1206)
);

AOI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1076),
.A2(n_1023),
.B1(n_1037),
.B2(n_1112),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1028),
.A2(n_1031),
.B(n_1094),
.Y(n_1208)
);

AOI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1131),
.A2(n_1102),
.B(n_1096),
.Y(n_1209)
);

INVx4_ASAP7_75t_SL g1210 ( 
.A(n_1098),
.Y(n_1210)
);

OA21x2_ASAP7_75t_L g1211 ( 
.A1(n_1155),
.A2(n_1081),
.B(n_1043),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_R g1212 ( 
.A(n_1145),
.B(n_1099),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1023),
.A2(n_1111),
.B1(n_1123),
.B2(n_1107),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1083),
.B(n_1033),
.Y(n_1214)
);

CKINVDCx20_ASAP7_75t_R g1215 ( 
.A(n_1127),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1140),
.A2(n_1046),
.B(n_1050),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1027),
.A2(n_1156),
.B(n_1068),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1104),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1065),
.B(n_1167),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_1127),
.Y(n_1220)
);

OR2x2_ASAP7_75t_L g1221 ( 
.A(n_1067),
.B(n_1059),
.Y(n_1221)
);

BUFx10_ASAP7_75t_L g1222 ( 
.A(n_1100),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1027),
.A2(n_1068),
.B(n_1129),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1055),
.B(n_1110),
.Y(n_1224)
);

AO31x2_ASAP7_75t_L g1225 ( 
.A1(n_1118),
.A2(n_1159),
.A3(n_1066),
.B(n_1136),
.Y(n_1225)
);

INVx4_ASAP7_75t_L g1226 ( 
.A(n_1094),
.Y(n_1226)
);

NAND3xp33_ASAP7_75t_SL g1227 ( 
.A(n_1122),
.B(n_1134),
.C(n_1073),
.Y(n_1227)
);

AO21x1_ASAP7_75t_L g1228 ( 
.A1(n_1049),
.A2(n_1118),
.B(n_1116),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1110),
.B(n_1100),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1094),
.A2(n_1146),
.B(n_1155),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1144),
.A2(n_1116),
.B(n_1105),
.C(n_1101),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1141),
.A2(n_1157),
.B(n_1161),
.Y(n_1232)
);

INVxp67_ASAP7_75t_L g1233 ( 
.A(n_1077),
.Y(n_1233)
);

NOR3xp33_ASAP7_75t_L g1234 ( 
.A(n_1057),
.B(n_1114),
.C(n_1071),
.Y(n_1234)
);

INVx1_ASAP7_75t_SL g1235 ( 
.A(n_1103),
.Y(n_1235)
);

INVx2_ASAP7_75t_SL g1236 ( 
.A(n_1124),
.Y(n_1236)
);

AO22x2_ASAP7_75t_L g1237 ( 
.A1(n_1021),
.A2(n_1087),
.B1(n_1088),
.B2(n_1082),
.Y(n_1237)
);

BUFx12f_ASAP7_75t_L g1238 ( 
.A(n_1089),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1034),
.B(n_1074),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1075),
.A2(n_1061),
.B(n_1161),
.Y(n_1240)
);

AO21x2_ASAP7_75t_L g1241 ( 
.A1(n_1148),
.A2(n_1161),
.B(n_1168),
.Y(n_1241)
);

A2O1A1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1161),
.A2(n_1120),
.B(n_1121),
.C(n_1041),
.Y(n_1242)
);

AOI221x1_ASAP7_75t_L g1243 ( 
.A1(n_1074),
.A2(n_1022),
.B1(n_1036),
.B2(n_1051),
.C(n_1058),
.Y(n_1243)
);

NAND2xp33_ASAP7_75t_SL g1244 ( 
.A(n_1022),
.B(n_1036),
.Y(n_1244)
);

NAND2x1_ASAP7_75t_L g1245 ( 
.A(n_1141),
.B(n_1151),
.Y(n_1245)
);

AOI211x1_ASAP7_75t_L g1246 ( 
.A1(n_1141),
.A2(n_1137),
.B(n_1151),
.C(n_1139),
.Y(n_1246)
);

INVxp67_ASAP7_75t_SL g1247 ( 
.A(n_1137),
.Y(n_1247)
);

O2A1O1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1098),
.A2(n_1063),
.B(n_1089),
.C(n_1051),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1139),
.A2(n_1062),
.B(n_1036),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1022),
.B(n_1051),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1058),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1058),
.A2(n_923),
.B(n_1154),
.Y(n_1252)
);

AO21x2_ASAP7_75t_L g1253 ( 
.A1(n_1062),
.A2(n_923),
.B(n_1162),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_1062),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1160),
.A2(n_923),
.B(n_874),
.Y(n_1255)
);

AO31x2_ASAP7_75t_L g1256 ( 
.A1(n_1158),
.A2(n_948),
.A3(n_923),
.B(n_1143),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1022),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1085),
.Y(n_1258)
);

BUFx3_ASAP7_75t_L g1259 ( 
.A(n_1054),
.Y(n_1259)
);

INVxp67_ASAP7_75t_L g1260 ( 
.A(n_1059),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_1022),
.Y(n_1261)
);

A2O1A1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1095),
.A2(n_874),
.B(n_923),
.C(n_1106),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_1054),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1085),
.Y(n_1264)
);

O2A1O1Ixp33_ASAP7_75t_SL g1265 ( 
.A1(n_1031),
.A2(n_923),
.B(n_1020),
.C(n_1092),
.Y(n_1265)
);

AO31x2_ASAP7_75t_L g1266 ( 
.A1(n_1158),
.A2(n_948),
.A3(n_923),
.B(n_1143),
.Y(n_1266)
);

AO31x2_ASAP7_75t_L g1267 ( 
.A1(n_1158),
.A2(n_948),
.A3(n_923),
.B(n_1143),
.Y(n_1267)
);

AOI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1095),
.A2(n_874),
.B1(n_1048),
.B2(n_1106),
.Y(n_1268)
);

BUFx6f_ASAP7_75t_L g1269 ( 
.A(n_1022),
.Y(n_1269)
);

AOI221x1_ASAP7_75t_L g1270 ( 
.A1(n_1048),
.A2(n_923),
.B1(n_1095),
.B2(n_874),
.C(n_1092),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1154),
.A2(n_923),
.B(n_1153),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1030),
.A2(n_1162),
.B(n_1069),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1154),
.A2(n_923),
.B(n_1153),
.Y(n_1273)
);

OA21x2_ASAP7_75t_L g1274 ( 
.A1(n_1097),
.A2(n_1158),
.B(n_1150),
.Y(n_1274)
);

INVxp67_ASAP7_75t_SL g1275 ( 
.A(n_1137),
.Y(n_1275)
);

A2O1A1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1095),
.A2(n_874),
.B(n_923),
.C(n_1106),
.Y(n_1276)
);

AO31x2_ASAP7_75t_L g1277 ( 
.A1(n_1158),
.A2(n_948),
.A3(n_923),
.B(n_1143),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1154),
.A2(n_923),
.B(n_1153),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1154),
.A2(n_923),
.B(n_1153),
.Y(n_1279)
);

AO32x2_ASAP7_75t_L g1280 ( 
.A1(n_1042),
.A2(n_794),
.A3(n_1126),
.B1(n_1166),
.B2(n_1090),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1022),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1085),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1092),
.B(n_874),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1154),
.A2(n_923),
.B(n_1153),
.Y(n_1284)
);

NAND2x1p5_ASAP7_75t_L g1285 ( 
.A(n_1094),
.B(n_853),
.Y(n_1285)
);

AO31x2_ASAP7_75t_L g1286 ( 
.A1(n_1158),
.A2(n_948),
.A3(n_923),
.B(n_1143),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1056),
.Y(n_1287)
);

A2O1A1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1095),
.A2(n_874),
.B(n_923),
.C(n_1106),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1154),
.A2(n_923),
.B(n_1153),
.Y(n_1289)
);

AO32x2_ASAP7_75t_L g1290 ( 
.A1(n_1042),
.A2(n_794),
.A3(n_1126),
.B1(n_1166),
.B2(n_1090),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1160),
.A2(n_923),
.B(n_874),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1154),
.A2(n_923),
.B(n_1153),
.Y(n_1292)
);

AO32x2_ASAP7_75t_L g1293 ( 
.A1(n_1042),
.A2(n_794),
.A3(n_1126),
.B1(n_1166),
.B2(n_1090),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1095),
.A2(n_874),
.B1(n_1048),
.B2(n_1106),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1030),
.A2(n_1162),
.B(n_1069),
.Y(n_1295)
);

NAND2x1_ASAP7_75t_L g1296 ( 
.A(n_1141),
.B(n_853),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1022),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1030),
.A2(n_1162),
.B(n_1069),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1037),
.B(n_527),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1085),
.Y(n_1300)
);

AO31x2_ASAP7_75t_L g1301 ( 
.A1(n_1158),
.A2(n_948),
.A3(n_923),
.B(n_1143),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1022),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1112),
.B(n_1100),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1154),
.A2(n_923),
.B(n_1153),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1154),
.A2(n_923),
.B(n_1153),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1154),
.A2(n_923),
.B(n_1153),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1092),
.B(n_874),
.Y(n_1307)
);

BUFx3_ASAP7_75t_L g1308 ( 
.A(n_1054),
.Y(n_1308)
);

NAND2x1p5_ASAP7_75t_L g1309 ( 
.A(n_1094),
.B(n_853),
.Y(n_1309)
);

CKINVDCx8_ASAP7_75t_R g1310 ( 
.A(n_1025),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_SL g1311 ( 
.A1(n_1118),
.A2(n_1070),
.B(n_837),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1037),
.B(n_527),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1154),
.A2(n_923),
.B(n_1153),
.Y(n_1313)
);

AOI221x1_ASAP7_75t_L g1314 ( 
.A1(n_1048),
.A2(n_923),
.B1(n_1095),
.B2(n_874),
.C(n_1092),
.Y(n_1314)
);

NOR2x1_ASAP7_75t_R g1315 ( 
.A(n_1018),
.B(n_671),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_SL g1316 ( 
.A(n_1092),
.B(n_527),
.Y(n_1316)
);

NOR2xp67_ASAP7_75t_L g1317 ( 
.A(n_1094),
.B(n_531),
.Y(n_1317)
);

AO21x1_ASAP7_75t_L g1318 ( 
.A1(n_1070),
.A2(n_874),
.B(n_1092),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1030),
.A2(n_1162),
.B(n_1069),
.Y(n_1319)
);

AO31x2_ASAP7_75t_L g1320 ( 
.A1(n_1158),
.A2(n_948),
.A3(n_923),
.B(n_1143),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1154),
.A2(n_923),
.B(n_1153),
.Y(n_1321)
);

OR2x6_ASAP7_75t_L g1322 ( 
.A(n_1141),
.B(n_716),
.Y(n_1322)
);

AO31x2_ASAP7_75t_L g1323 ( 
.A1(n_1158),
.A2(n_948),
.A3(n_923),
.B(n_1143),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1160),
.A2(n_923),
.B(n_874),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1259),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1294),
.A2(n_1268),
.B1(n_1187),
.B2(n_1204),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1196),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1258),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_1263),
.Y(n_1329)
);

CKINVDCx11_ASAP7_75t_R g1330 ( 
.A(n_1310),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_1257),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_SL g1332 ( 
.A1(n_1268),
.A2(n_1189),
.B1(n_1215),
.B2(n_1307),
.Y(n_1332)
);

BUFx4f_ASAP7_75t_SL g1333 ( 
.A(n_1238),
.Y(n_1333)
);

CKINVDCx11_ASAP7_75t_R g1334 ( 
.A(n_1186),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1283),
.B(n_1198),
.Y(n_1335)
);

AOI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1189),
.A2(n_1227),
.B1(n_1276),
.B2(n_1288),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_SL g1337 ( 
.A1(n_1204),
.A2(n_1311),
.B1(n_1212),
.B2(n_1229),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1199),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_SL g1339 ( 
.A1(n_1200),
.A2(n_1312),
.B1(n_1299),
.B2(n_1224),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1264),
.Y(n_1340)
);

INVx2_ASAP7_75t_SL g1341 ( 
.A(n_1308),
.Y(n_1341)
);

OAI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1270),
.A2(n_1314),
.B1(n_1182),
.B2(n_1207),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1282),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1300),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1318),
.A2(n_1234),
.B1(n_1324),
.B2(n_1255),
.Y(n_1345)
);

OAI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1207),
.A2(n_1213),
.B1(n_1219),
.B2(n_1316),
.Y(n_1346)
);

INVx4_ASAP7_75t_L g1347 ( 
.A(n_1210),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1324),
.A2(n_1255),
.B1(n_1291),
.B2(n_1213),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1169),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1262),
.A2(n_1194),
.B1(n_1190),
.B2(n_1195),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1195),
.A2(n_1231),
.B1(n_1235),
.B2(n_1260),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1214),
.Y(n_1352)
);

BUFx12f_ASAP7_75t_L g1353 ( 
.A(n_1220),
.Y(n_1353)
);

INVx3_ASAP7_75t_L g1354 ( 
.A(n_1239),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1237),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1251),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1291),
.A2(n_1228),
.B1(n_1278),
.B2(n_1305),
.Y(n_1357)
);

INVx1_ASAP7_75t_SL g1358 ( 
.A(n_1221),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1235),
.A2(n_1233),
.B1(n_1303),
.B2(n_1203),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1303),
.A2(n_1287),
.B1(n_1322),
.B2(n_1174),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_SL g1361 ( 
.A1(n_1241),
.A2(n_1174),
.B1(n_1275),
.B2(n_1247),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_1257),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1322),
.A2(n_1252),
.B1(n_1321),
.B2(n_1313),
.Y(n_1363)
);

CKINVDCx11_ASAP7_75t_R g1364 ( 
.A(n_1191),
.Y(n_1364)
);

CKINVDCx11_ASAP7_75t_R g1365 ( 
.A(n_1210),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1271),
.A2(n_1279),
.B1(n_1304),
.B2(n_1273),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1250),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1284),
.A2(n_1306),
.B1(n_1289),
.B2(n_1292),
.Y(n_1368)
);

NAND2x1p5_ASAP7_75t_L g1369 ( 
.A(n_1226),
.B(n_1296),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1254),
.Y(n_1370)
);

CKINVDCx11_ASAP7_75t_R g1371 ( 
.A(n_1222),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_SL g1372 ( 
.A1(n_1241),
.A2(n_1222),
.B1(n_1183),
.B2(n_1185),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1243),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_1257),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1236),
.Y(n_1375)
);

CKINVDCx6p67_ASAP7_75t_R g1376 ( 
.A(n_1322),
.Y(n_1376)
);

CKINVDCx20_ASAP7_75t_R g1377 ( 
.A(n_1218),
.Y(n_1377)
);

INVx6_ASAP7_75t_L g1378 ( 
.A(n_1239),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1253),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1261),
.B(n_1269),
.Y(n_1380)
);

INVx3_ASAP7_75t_SL g1381 ( 
.A(n_1261),
.Y(n_1381)
);

OAI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1172),
.A2(n_1185),
.B1(n_1183),
.B2(n_1181),
.Y(n_1382)
);

BUFx2_ASAP7_75t_SL g1383 ( 
.A(n_1205),
.Y(n_1383)
);

AOI22xp5_ASAP7_75t_SL g1384 ( 
.A1(n_1232),
.A2(n_1230),
.B1(n_1315),
.B2(n_1249),
.Y(n_1384)
);

BUFx3_ASAP7_75t_L g1385 ( 
.A(n_1269),
.Y(n_1385)
);

BUFx4_ASAP7_75t_SL g1386 ( 
.A(n_1315),
.Y(n_1386)
);

AOI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1265),
.A2(n_1317),
.B1(n_1177),
.B2(n_1179),
.Y(n_1387)
);

CKINVDCx11_ASAP7_75t_R g1388 ( 
.A(n_1269),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1281),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1246),
.A2(n_1317),
.B1(n_1242),
.B2(n_1240),
.Y(n_1390)
);

BUFx12f_ASAP7_75t_L g1391 ( 
.A(n_1281),
.Y(n_1391)
);

BUFx12f_ASAP7_75t_L g1392 ( 
.A(n_1281),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1188),
.A2(n_1178),
.B(n_1202),
.Y(n_1393)
);

CKINVDCx11_ASAP7_75t_R g1394 ( 
.A(n_1297),
.Y(n_1394)
);

OAI21xp5_ASAP7_75t_SL g1395 ( 
.A1(n_1248),
.A2(n_1209),
.B(n_1197),
.Y(n_1395)
);

AOI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1244),
.A2(n_1245),
.B1(n_1211),
.B2(n_1205),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1297),
.Y(n_1397)
);

OAI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1184),
.A2(n_1211),
.B1(n_1274),
.B2(n_1293),
.Y(n_1398)
);

CKINVDCx20_ASAP7_75t_R g1399 ( 
.A(n_1297),
.Y(n_1399)
);

CKINVDCx11_ASAP7_75t_R g1400 ( 
.A(n_1302),
.Y(n_1400)
);

INVx6_ASAP7_75t_L g1401 ( 
.A(n_1302),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1246),
.A2(n_1309),
.B1(n_1285),
.B2(n_1208),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1274),
.A2(n_1184),
.B1(n_1201),
.B2(n_1280),
.Y(n_1403)
);

BUFx10_ASAP7_75t_L g1404 ( 
.A(n_1173),
.Y(n_1404)
);

BUFx12f_ASAP7_75t_L g1405 ( 
.A(n_1225),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_1176),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_1216),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1184),
.A2(n_1201),
.B1(n_1176),
.B2(n_1280),
.Y(n_1408)
);

BUFx12f_ASAP7_75t_L g1409 ( 
.A(n_1225),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1256),
.Y(n_1410)
);

INVx1_ASAP7_75t_SL g1411 ( 
.A(n_1171),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1280),
.A2(n_1293),
.B1(n_1290),
.B2(n_1323),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1290),
.A2(n_1293),
.B1(n_1171),
.B2(n_1272),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1290),
.A2(n_1295),
.B1(n_1319),
.B2(n_1298),
.Y(n_1414)
);

INVx6_ASAP7_75t_L g1415 ( 
.A(n_1206),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1256),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1256),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_SL g1418 ( 
.A1(n_1193),
.A2(n_1266),
.B1(n_1320),
.B2(n_1301),
.Y(n_1418)
);

CKINVDCx11_ASAP7_75t_R g1419 ( 
.A(n_1266),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1266),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_SL g1421 ( 
.A1(n_1267),
.A2(n_1323),
.B1(n_1320),
.B2(n_1301),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1217),
.A2(n_1223),
.B1(n_1170),
.B2(n_1175),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1192),
.A2(n_1267),
.B1(n_1277),
.B2(n_1286),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1301),
.B(n_1277),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1277),
.B(n_1286),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1180),
.A2(n_1095),
.B1(n_1294),
.B2(n_874),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1180),
.A2(n_1095),
.B1(n_1294),
.B2(n_874),
.Y(n_1427)
);

BUFx8_ASAP7_75t_L g1428 ( 
.A(n_1206),
.Y(n_1428)
);

CKINVDCx11_ASAP7_75t_R g1429 ( 
.A(n_1180),
.Y(n_1429)
);

INVx1_ASAP7_75t_SL g1430 ( 
.A(n_1195),
.Y(n_1430)
);

CKINVDCx20_ASAP7_75t_R g1431 ( 
.A(n_1191),
.Y(n_1431)
);

BUFx12f_ASAP7_75t_L g1432 ( 
.A(n_1238),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_SL g1433 ( 
.A1(n_1189),
.A2(n_1095),
.B1(n_980),
.B2(n_1092),
.Y(n_1433)
);

INVx3_ASAP7_75t_L g1434 ( 
.A(n_1239),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1294),
.A2(n_1095),
.B1(n_874),
.B2(n_1268),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1294),
.A2(n_1095),
.B1(n_874),
.B2(n_1268),
.Y(n_1436)
);

BUFx10_ASAP7_75t_L g1437 ( 
.A(n_1220),
.Y(n_1437)
);

OAI22xp33_ASAP7_75t_SL g1438 ( 
.A1(n_1268),
.A2(n_1092),
.B1(n_1095),
.B2(n_1060),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1268),
.A2(n_1048),
.B1(n_874),
.B2(n_1095),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1294),
.A2(n_1268),
.B1(n_1092),
.B2(n_1262),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1294),
.A2(n_1095),
.B1(n_874),
.B2(n_1268),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1294),
.A2(n_1268),
.B1(n_1092),
.B2(n_1262),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1294),
.A2(n_1095),
.B1(n_874),
.B2(n_1268),
.Y(n_1443)
);

BUFx8_ASAP7_75t_L g1444 ( 
.A(n_1238),
.Y(n_1444)
);

BUFx3_ASAP7_75t_L g1445 ( 
.A(n_1259),
.Y(n_1445)
);

INVx3_ASAP7_75t_SL g1446 ( 
.A(n_1210),
.Y(n_1446)
);

CKINVDCx14_ASAP7_75t_R g1447 ( 
.A(n_1215),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1169),
.Y(n_1448)
);

INVx6_ASAP7_75t_L g1449 ( 
.A(n_1210),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1283),
.B(n_1307),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1294),
.A2(n_1095),
.B1(n_874),
.B2(n_1268),
.Y(n_1451)
);

OA21x2_ASAP7_75t_L g1452 ( 
.A1(n_1393),
.A2(n_1348),
.B(n_1345),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1335),
.B(n_1450),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1355),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1417),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1420),
.Y(n_1456)
);

NOR2x1_ASAP7_75t_L g1457 ( 
.A(n_1395),
.B(n_1346),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1358),
.B(n_1332),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_SL g1459 ( 
.A1(n_1350),
.A2(n_1390),
.B(n_1336),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1351),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1424),
.B(n_1425),
.Y(n_1461)
);

AO21x2_ASAP7_75t_L g1462 ( 
.A1(n_1342),
.A2(n_1382),
.B(n_1398),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1422),
.A2(n_1363),
.B(n_1414),
.Y(n_1463)
);

AO21x2_ASAP7_75t_L g1464 ( 
.A1(n_1342),
.A2(n_1382),
.B(n_1398),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1431),
.B(n_1430),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1410),
.Y(n_1466)
);

BUFx12f_ASAP7_75t_L g1467 ( 
.A(n_1330),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1364),
.Y(n_1468)
);

INVxp67_ASAP7_75t_L g1469 ( 
.A(n_1448),
.Y(n_1469)
);

BUFx3_ASAP7_75t_L g1470 ( 
.A(n_1376),
.Y(n_1470)
);

CKINVDCx11_ASAP7_75t_R g1471 ( 
.A(n_1334),
.Y(n_1471)
);

INVxp67_ASAP7_75t_L g1472 ( 
.A(n_1349),
.Y(n_1472)
);

BUFx3_ASAP7_75t_L g1473 ( 
.A(n_1428),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1379),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1415),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1422),
.A2(n_1414),
.B(n_1366),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1416),
.B(n_1348),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1366),
.A2(n_1368),
.B(n_1357),
.Y(n_1478)
);

OAI222xp33_ASAP7_75t_L g1479 ( 
.A1(n_1439),
.A2(n_1433),
.B1(n_1435),
.B2(n_1443),
.C1(n_1441),
.C2(n_1451),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1421),
.Y(n_1480)
);

INVx2_ASAP7_75t_SL g1481 ( 
.A(n_1449),
.Y(n_1481)
);

INVx5_ASAP7_75t_L g1482 ( 
.A(n_1407),
.Y(n_1482)
);

BUFx2_ASAP7_75t_R g1483 ( 
.A(n_1446),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1345),
.B(n_1326),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1370),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1428),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1367),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1435),
.A2(n_1443),
.B1(n_1451),
.B2(n_1436),
.Y(n_1488)
);

CKINVDCx20_ASAP7_75t_R g1489 ( 
.A(n_1447),
.Y(n_1489)
);

AO21x2_ASAP7_75t_L g1490 ( 
.A1(n_1387),
.A2(n_1408),
.B(n_1412),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1405),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1409),
.Y(n_1492)
);

CKINVDCx14_ASAP7_75t_R g1493 ( 
.A(n_1447),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1338),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1377),
.B(n_1349),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1436),
.A2(n_1441),
.B1(n_1442),
.B2(n_1440),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1340),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1373),
.Y(n_1498)
);

BUFx12f_ASAP7_75t_L g1499 ( 
.A(n_1365),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1343),
.Y(n_1500)
);

INVx3_ASAP7_75t_L g1501 ( 
.A(n_1407),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1368),
.A2(n_1357),
.B(n_1423),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1396),
.B(n_1384),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1407),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1404),
.Y(n_1505)
);

CKINVDCx6p67_ASAP7_75t_R g1506 ( 
.A(n_1446),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1429),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1411),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1419),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1406),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1344),
.Y(n_1511)
);

INVx3_ASAP7_75t_SL g1512 ( 
.A(n_1449),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1419),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1418),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1354),
.B(n_1434),
.Y(n_1515)
);

OAI21x1_ASAP7_75t_L g1516 ( 
.A1(n_1423),
.A2(n_1413),
.B(n_1403),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1403),
.Y(n_1517)
);

A2O1A1Ixp33_ASAP7_75t_L g1518 ( 
.A1(n_1326),
.A2(n_1426),
.B(n_1427),
.C(n_1372),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1327),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1352),
.B(n_1339),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1328),
.Y(n_1521)
);

BUFx2_ASAP7_75t_L g1522 ( 
.A(n_1360),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1413),
.B(n_1427),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_1386),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1386),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1359),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1346),
.Y(n_1527)
);

AOI21xp33_ASAP7_75t_L g1528 ( 
.A1(n_1438),
.A2(n_1426),
.B(n_1337),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1356),
.Y(n_1529)
);

INVxp67_ASAP7_75t_L g1530 ( 
.A(n_1325),
.Y(n_1530)
);

INVxp67_ASAP7_75t_L g1531 ( 
.A(n_1325),
.Y(n_1531)
);

OAI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1361),
.A2(n_1402),
.B(n_1369),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1380),
.B(n_1354),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1369),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1383),
.Y(n_1535)
);

OA21x2_ASAP7_75t_L g1536 ( 
.A1(n_1397),
.A2(n_1341),
.B(n_1331),
.Y(n_1536)
);

OAI21x1_ASAP7_75t_L g1537 ( 
.A1(n_1434),
.A2(n_1449),
.B(n_1371),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1371),
.A2(n_1378),
.B(n_1381),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1529),
.Y(n_1539)
);

NOR2x1_ASAP7_75t_SL g1540 ( 
.A(n_1473),
.B(n_1347),
.Y(n_1540)
);

OR2x6_ASAP7_75t_L g1541 ( 
.A(n_1503),
.B(n_1347),
.Y(n_1541)
);

CKINVDCx20_ASAP7_75t_R g1542 ( 
.A(n_1471),
.Y(n_1542)
);

AND2x2_ASAP7_75t_SL g1543 ( 
.A(n_1452),
.B(n_1374),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1455),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1517),
.B(n_1389),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1491),
.B(n_1385),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1490),
.B(n_1374),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1491),
.B(n_1385),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1453),
.B(n_1445),
.Y(n_1549)
);

OAI211xp5_ASAP7_75t_L g1550 ( 
.A1(n_1528),
.A2(n_1388),
.B(n_1400),
.C(n_1394),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1492),
.B(n_1486),
.Y(n_1551)
);

BUFx3_ASAP7_75t_L g1552 ( 
.A(n_1512),
.Y(n_1552)
);

INVx11_ASAP7_75t_L g1553 ( 
.A(n_1467),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1467),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1490),
.B(n_1523),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1492),
.B(n_1331),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1487),
.B(n_1445),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1514),
.B(n_1362),
.Y(n_1558)
);

A2O1A1Ixp33_ASAP7_75t_L g1559 ( 
.A1(n_1457),
.A2(n_1329),
.B(n_1399),
.C(n_1331),
.Y(n_1559)
);

INVx2_ASAP7_75t_SL g1560 ( 
.A(n_1536),
.Y(n_1560)
);

A2O1A1Ixp33_ASAP7_75t_L g1561 ( 
.A1(n_1457),
.A2(n_1329),
.B(n_1374),
.C(n_1362),
.Y(n_1561)
);

AOI21xp5_ASAP7_75t_L g1562 ( 
.A1(n_1452),
.A2(n_1378),
.B(n_1375),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1475),
.B(n_1388),
.Y(n_1563)
);

NOR4xp25_ASAP7_75t_SL g1564 ( 
.A(n_1528),
.B(n_1444),
.C(n_1333),
.D(n_1432),
.Y(n_1564)
);

A2O1A1Ixp33_ASAP7_75t_L g1565 ( 
.A1(n_1518),
.A2(n_1437),
.B(n_1391),
.C(n_1392),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1520),
.B(n_1401),
.Y(n_1566)
);

O2A1O1Ixp33_ASAP7_75t_L g1567 ( 
.A1(n_1479),
.A2(n_1333),
.B(n_1437),
.C(n_1444),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1465),
.B(n_1353),
.Y(n_1568)
);

INVx11_ASAP7_75t_L g1569 ( 
.A(n_1467),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1510),
.B(n_1495),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1516),
.B(n_1494),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1461),
.B(n_1498),
.Y(n_1572)
);

NOR2x1_ASAP7_75t_L g1573 ( 
.A(n_1535),
.B(n_1470),
.Y(n_1573)
);

OAI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1496),
.A2(n_1488),
.B(n_1527),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1516),
.B(n_1494),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1488),
.A2(n_1458),
.B1(n_1460),
.B2(n_1477),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_SL g1577 ( 
.A(n_1483),
.B(n_1468),
.Y(n_1577)
);

A2O1A1Ixp33_ASAP7_75t_L g1578 ( 
.A1(n_1527),
.A2(n_1484),
.B(n_1503),
.C(n_1532),
.Y(n_1578)
);

AO21x1_ASAP7_75t_L g1579 ( 
.A1(n_1484),
.A2(n_1480),
.B(n_1477),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1510),
.B(n_1526),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1497),
.B(n_1500),
.Y(n_1581)
);

AOI211xp5_ASAP7_75t_L g1582 ( 
.A1(n_1503),
.A2(n_1532),
.B(n_1507),
.C(n_1522),
.Y(n_1582)
);

OA21x2_ASAP7_75t_L g1583 ( 
.A1(n_1476),
.A2(n_1463),
.B(n_1502),
.Y(n_1583)
);

O2A1O1Ixp33_ASAP7_75t_SL g1584 ( 
.A1(n_1489),
.A2(n_1481),
.B(n_1507),
.C(n_1480),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1497),
.B(n_1500),
.Y(n_1585)
);

AOI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1503),
.A2(n_1522),
.B1(n_1493),
.B2(n_1513),
.Y(n_1586)
);

OA21x2_ASAP7_75t_L g1587 ( 
.A1(n_1463),
.A2(n_1502),
.B(n_1478),
.Y(n_1587)
);

INVxp67_ASAP7_75t_L g1588 ( 
.A(n_1485),
.Y(n_1588)
);

OR2x6_ASAP7_75t_L g1589 ( 
.A(n_1478),
.B(n_1473),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1461),
.B(n_1498),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1506),
.A2(n_1513),
.B1(n_1509),
.B2(n_1530),
.Y(n_1591)
);

NOR2x1_ASAP7_75t_SL g1592 ( 
.A(n_1473),
.B(n_1462),
.Y(n_1592)
);

AO21x2_ASAP7_75t_L g1593 ( 
.A1(n_1462),
.A2(n_1464),
.B(n_1505),
.Y(n_1593)
);

AO21x2_ASAP7_75t_L g1594 ( 
.A1(n_1462),
.A2(n_1464),
.B(n_1505),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1536),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1464),
.B(n_1454),
.Y(n_1596)
);

A2O1A1Ixp33_ASAP7_75t_L g1597 ( 
.A1(n_1509),
.A2(n_1513),
.B(n_1470),
.C(n_1459),
.Y(n_1597)
);

AOI21xp33_ASAP7_75t_L g1598 ( 
.A1(n_1576),
.A2(n_1459),
.B(n_1464),
.Y(n_1598)
);

INVxp67_ASAP7_75t_L g1599 ( 
.A(n_1580),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1544),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1549),
.B(n_1531),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1539),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1572),
.B(n_1474),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1572),
.B(n_1474),
.Y(n_1604)
);

BUFx3_ASAP7_75t_L g1605 ( 
.A(n_1552),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1555),
.B(n_1509),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1590),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1574),
.A2(n_1452),
.B1(n_1499),
.B2(n_1515),
.Y(n_1608)
);

INVx2_ASAP7_75t_SL g1609 ( 
.A(n_1551),
.Y(n_1609)
);

NOR2x1_ASAP7_75t_L g1610 ( 
.A(n_1573),
.B(n_1536),
.Y(n_1610)
);

AOI21xp33_ASAP7_75t_L g1611 ( 
.A1(n_1579),
.A2(n_1452),
.B(n_1508),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1579),
.A2(n_1499),
.B1(n_1515),
.B2(n_1470),
.Y(n_1612)
);

INVxp67_ASAP7_75t_L g1613 ( 
.A(n_1557),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1582),
.B(n_1515),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1581),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1571),
.B(n_1504),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1575),
.B(n_1504),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1541),
.A2(n_1499),
.B1(n_1515),
.B2(n_1534),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1575),
.B(n_1501),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1581),
.Y(n_1620)
);

AND2x4_ASAP7_75t_SL g1621 ( 
.A(n_1541),
.B(n_1563),
.Y(n_1621)
);

AOI222xp33_ASAP7_75t_L g1622 ( 
.A1(n_1578),
.A2(n_1469),
.B1(n_1525),
.B2(n_1524),
.C1(n_1472),
.C2(n_1511),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1560),
.Y(n_1623)
);

INVxp67_ASAP7_75t_L g1624 ( 
.A(n_1595),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1541),
.A2(n_1534),
.B1(n_1535),
.B2(n_1533),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1590),
.B(n_1529),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1585),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1596),
.B(n_1466),
.Y(n_1628)
);

NAND2x1p5_ASAP7_75t_L g1629 ( 
.A(n_1543),
.B(n_1482),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1547),
.B(n_1456),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1547),
.B(n_1456),
.Y(n_1631)
);

INVx3_ASAP7_75t_L g1632 ( 
.A(n_1619),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1613),
.B(n_1591),
.Y(n_1633)
);

AOI222xp33_ASAP7_75t_L g1634 ( 
.A1(n_1608),
.A2(n_1550),
.B1(n_1565),
.B2(n_1570),
.C1(n_1599),
.C2(n_1612),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1623),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1598),
.A2(n_1541),
.B1(n_1586),
.B2(n_1551),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1600),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1610),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1607),
.B(n_1626),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1600),
.Y(n_1640)
);

OAI21xp5_ASAP7_75t_SL g1641 ( 
.A1(n_1622),
.A2(n_1567),
.B(n_1559),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1606),
.B(n_1583),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1626),
.B(n_1588),
.Y(n_1643)
);

AOI21x1_ASAP7_75t_L g1644 ( 
.A1(n_1610),
.A2(n_1562),
.B(n_1589),
.Y(n_1644)
);

INVx1_ASAP7_75t_SL g1645 ( 
.A(n_1603),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_SL g1646 ( 
.A(n_1598),
.B(n_1561),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1624),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1628),
.Y(n_1648)
);

BUFx3_ASAP7_75t_L g1649 ( 
.A(n_1629),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1614),
.A2(n_1597),
.B1(n_1564),
.B2(n_1566),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1603),
.B(n_1593),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1602),
.Y(n_1652)
);

AOI221xp5_ASAP7_75t_L g1653 ( 
.A1(n_1611),
.A2(n_1584),
.B1(n_1551),
.B2(n_1519),
.C(n_1521),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1630),
.B(n_1592),
.Y(n_1654)
);

NAND4xp25_ASAP7_75t_L g1655 ( 
.A(n_1622),
.B(n_1577),
.C(n_1568),
.D(n_1545),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1631),
.B(n_1592),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1619),
.B(n_1589),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_SL g1658 ( 
.A(n_1629),
.B(n_1563),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1602),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1631),
.B(n_1587),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1604),
.B(n_1594),
.Y(n_1661)
);

INVx3_ASAP7_75t_L g1662 ( 
.A(n_1619),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1647),
.B(n_1615),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1635),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1651),
.B(n_1604),
.Y(n_1665)
);

AND2x2_ASAP7_75t_SL g1666 ( 
.A(n_1646),
.B(n_1621),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1652),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1635),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1651),
.B(n_1615),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1647),
.B(n_1645),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1651),
.B(n_1620),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1645),
.B(n_1620),
.Y(n_1672)
);

INVx3_ASAP7_75t_L g1673 ( 
.A(n_1657),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1652),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1660),
.B(n_1619),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1657),
.B(n_1632),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1635),
.Y(n_1677)
);

NAND3xp33_ASAP7_75t_L g1678 ( 
.A(n_1646),
.B(n_1611),
.C(n_1601),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1648),
.B(n_1627),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1652),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1648),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1635),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1637),
.B(n_1627),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1652),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1659),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1642),
.B(n_1616),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1642),
.B(n_1616),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1642),
.B(n_1654),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_SL g1689 ( 
.A(n_1650),
.B(n_1605),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1654),
.B(n_1616),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1659),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1654),
.B(n_1656),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1637),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1656),
.B(n_1617),
.Y(n_1694)
);

NOR3xp33_ASAP7_75t_SL g1695 ( 
.A(n_1641),
.B(n_1554),
.C(n_1553),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1640),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1640),
.Y(n_1697)
);

NOR2x1_ASAP7_75t_L g1698 ( 
.A(n_1689),
.B(n_1542),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1693),
.Y(n_1699)
);

INVx1_ASAP7_75t_SL g1700 ( 
.A(n_1666),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1693),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1678),
.B(n_1633),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_1666),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1693),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1681),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1676),
.B(n_1649),
.Y(n_1706)
);

INVxp67_ASAP7_75t_L g1707 ( 
.A(n_1689),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1678),
.B(n_1633),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1666),
.B(n_1657),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1696),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1664),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1696),
.Y(n_1712)
);

NAND2x1p5_ASAP7_75t_L g1713 ( 
.A(n_1666),
.B(n_1644),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1696),
.Y(n_1714)
);

NOR2x1_ASAP7_75t_L g1715 ( 
.A(n_1670),
.B(n_1542),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1697),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1681),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1670),
.B(n_1643),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1697),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1665),
.B(n_1661),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1697),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1692),
.B(n_1657),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1665),
.B(n_1661),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1692),
.B(n_1657),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1685),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1692),
.B(n_1632),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1673),
.B(n_1632),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1685),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1663),
.B(n_1643),
.Y(n_1729)
);

BUFx3_ASAP7_75t_L g1730 ( 
.A(n_1663),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1685),
.Y(n_1731)
);

INVx2_ASAP7_75t_SL g1732 ( 
.A(n_1673),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1672),
.B(n_1639),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1691),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1691),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1691),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1683),
.Y(n_1737)
);

NAND2x1_ASAP7_75t_L g1738 ( 
.A(n_1673),
.B(n_1632),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1672),
.B(n_1639),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1664),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1702),
.B(n_1695),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1709),
.B(n_1676),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1705),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1717),
.B(n_1665),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1704),
.Y(n_1745)
);

BUFx2_ASAP7_75t_L g1746 ( 
.A(n_1715),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1708),
.B(n_1695),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1729),
.B(n_1669),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1709),
.B(n_1673),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1707),
.B(n_1698),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1730),
.B(n_1718),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1704),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_SL g1753 ( 
.A(n_1700),
.B(n_1703),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_L g1754 ( 
.A(n_1733),
.B(n_1554),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1730),
.B(n_1669),
.Y(n_1755)
);

CKINVDCx16_ASAP7_75t_R g1756 ( 
.A(n_1706),
.Y(n_1756)
);

INVx4_ASAP7_75t_L g1757 ( 
.A(n_1713),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1722),
.B(n_1673),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1739),
.B(n_1737),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1712),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1722),
.B(n_1673),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1712),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1732),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1737),
.B(n_1656),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1724),
.B(n_1676),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1714),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1714),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1716),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1706),
.B(n_1553),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1732),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1726),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1706),
.B(n_1569),
.Y(n_1772)
);

NAND2x1_ASAP7_75t_L g1773 ( 
.A(n_1724),
.B(n_1676),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1720),
.B(n_1669),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1720),
.B(n_1671),
.Y(n_1775)
);

OAI21xp33_ASAP7_75t_L g1776 ( 
.A1(n_1713),
.A2(n_1641),
.B(n_1655),
.Y(n_1776)
);

OAI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1746),
.A2(n_1650),
.B1(n_1713),
.B2(n_1636),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1745),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1752),
.Y(n_1779)
);

OAI321xp33_ASAP7_75t_L g1780 ( 
.A1(n_1776),
.A2(n_1753),
.A3(n_1750),
.B1(n_1747),
.B2(n_1741),
.C(n_1655),
.Y(n_1780)
);

AOI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1753),
.A2(n_1772),
.B(n_1769),
.Y(n_1781)
);

AOI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1756),
.A2(n_1634),
.B1(n_1658),
.B2(n_1653),
.Y(n_1782)
);

AO22x1_ASAP7_75t_L g1783 ( 
.A1(n_1757),
.A2(n_1638),
.B1(n_1649),
.B2(n_1676),
.Y(n_1783)
);

NAND2xp33_ASAP7_75t_L g1784 ( 
.A(n_1751),
.B(n_1658),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1742),
.Y(n_1785)
);

AOI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1742),
.A2(n_1634),
.B1(n_1653),
.B2(n_1636),
.Y(n_1786)
);

AOI211x1_ASAP7_75t_L g1787 ( 
.A1(n_1743),
.A2(n_1644),
.B(n_1726),
.C(n_1727),
.Y(n_1787)
);

OAI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1751),
.A2(n_1649),
.B1(n_1638),
.B2(n_1618),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1760),
.Y(n_1789)
);

INVx3_ASAP7_75t_L g1790 ( 
.A(n_1773),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_L g1791 ( 
.A(n_1754),
.B(n_1569),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1762),
.Y(n_1792)
);

OAI31xp33_ASAP7_75t_L g1793 ( 
.A1(n_1749),
.A2(n_1649),
.A3(n_1727),
.B(n_1676),
.Y(n_1793)
);

NOR2xp33_ASAP7_75t_L g1794 ( 
.A(n_1757),
.B(n_1506),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1766),
.Y(n_1795)
);

OAI221xp5_ASAP7_75t_L g1796 ( 
.A1(n_1757),
.A2(n_1738),
.B1(n_1721),
.B2(n_1699),
.C(n_1701),
.Y(n_1796)
);

BUFx3_ASAP7_75t_L g1797 ( 
.A(n_1763),
.Y(n_1797)
);

INVxp67_ASAP7_75t_SL g1798 ( 
.A(n_1763),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1742),
.B(n_1690),
.Y(n_1799)
);

A2O1A1Ixp33_ASAP7_75t_L g1800 ( 
.A1(n_1755),
.A2(n_1744),
.B(n_1759),
.C(n_1749),
.Y(n_1800)
);

OAI21xp33_ASAP7_75t_SL g1801 ( 
.A1(n_1765),
.A2(n_1688),
.B(n_1710),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1759),
.B(n_1723),
.Y(n_1802)
);

OAI21xp5_ASAP7_75t_SL g1803 ( 
.A1(n_1782),
.A2(n_1765),
.B(n_1761),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1798),
.Y(n_1804)
);

AOI322xp5_ASAP7_75t_L g1805 ( 
.A1(n_1786),
.A2(n_1764),
.A3(n_1771),
.B1(n_1758),
.B2(n_1761),
.C1(n_1688),
.C2(n_1767),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1790),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1800),
.B(n_1744),
.Y(n_1807)
);

AOI32xp33_ASAP7_75t_L g1808 ( 
.A1(n_1780),
.A2(n_1771),
.A3(n_1758),
.B1(n_1755),
.B2(n_1770),
.Y(n_1808)
);

OAI221xp5_ASAP7_75t_L g1809 ( 
.A1(n_1777),
.A2(n_1748),
.B1(n_1768),
.B2(n_1770),
.C(n_1738),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1781),
.A2(n_1748),
.B1(n_1589),
.B2(n_1621),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1798),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1800),
.B(n_1774),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1778),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1779),
.B(n_1716),
.Y(n_1814)
);

INVxp67_ASAP7_75t_L g1815 ( 
.A(n_1794),
.Y(n_1815)
);

AOI21xp33_ASAP7_75t_L g1816 ( 
.A1(n_1794),
.A2(n_1725),
.B(n_1719),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1789),
.B(n_1719),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1785),
.B(n_1675),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1792),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1799),
.B(n_1675),
.Y(n_1820)
);

AO22x1_ASAP7_75t_L g1821 ( 
.A1(n_1790),
.A2(n_1512),
.B1(n_1734),
.B2(n_1728),
.Y(n_1821)
);

OR2x6_ASAP7_75t_L g1822 ( 
.A(n_1797),
.B(n_1481),
.Y(n_1822)
);

INVxp67_ASAP7_75t_L g1823 ( 
.A(n_1807),
.Y(n_1823)
);

O2A1O1Ixp33_ASAP7_75t_L g1824 ( 
.A1(n_1812),
.A2(n_1784),
.B(n_1788),
.C(n_1797),
.Y(n_1824)
);

AOI21xp33_ASAP7_75t_L g1825 ( 
.A1(n_1815),
.A2(n_1802),
.B(n_1796),
.Y(n_1825)
);

XNOR2xp5_ASAP7_75t_L g1826 ( 
.A(n_1809),
.B(n_1563),
.Y(n_1826)
);

O2A1O1Ixp33_ASAP7_75t_L g1827 ( 
.A1(n_1804),
.A2(n_1795),
.B(n_1801),
.C(n_1793),
.Y(n_1827)
);

XOR2x2_ASAP7_75t_L g1828 ( 
.A(n_1811),
.B(n_1791),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1806),
.B(n_1787),
.Y(n_1829)
);

OAI221xp5_ASAP7_75t_L g1830 ( 
.A1(n_1803),
.A2(n_1791),
.B1(n_1774),
.B2(n_1775),
.C(n_1734),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1813),
.B(n_1783),
.Y(n_1831)
);

INVx3_ASAP7_75t_L g1832 ( 
.A(n_1822),
.Y(n_1832)
);

INVxp67_ASAP7_75t_L g1833 ( 
.A(n_1822),
.Y(n_1833)
);

INVx1_ASAP7_75t_SL g1834 ( 
.A(n_1822),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1823),
.B(n_1808),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_SL g1836 ( 
.A(n_1824),
.B(n_1834),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1828),
.B(n_1818),
.Y(n_1837)
);

AOI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1826),
.A2(n_1810),
.B1(n_1819),
.B2(n_1820),
.Y(n_1838)
);

AOI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1829),
.A2(n_1816),
.B(n_1821),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1832),
.Y(n_1840)
);

NAND4xp25_ASAP7_75t_L g1841 ( 
.A(n_1825),
.B(n_1805),
.C(n_1816),
.D(n_1814),
.Y(n_1841)
);

CKINVDCx20_ASAP7_75t_R g1842 ( 
.A(n_1833),
.Y(n_1842)
);

AOI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1831),
.A2(n_1817),
.B1(n_1814),
.B2(n_1731),
.Y(n_1843)
);

OAI222xp33_ASAP7_75t_L g1844 ( 
.A1(n_1830),
.A2(n_1817),
.B1(n_1775),
.B2(n_1644),
.C1(n_1723),
.C2(n_1735),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1832),
.B(n_1675),
.Y(n_1845)
);

NAND4xp25_ASAP7_75t_L g1846 ( 
.A(n_1827),
.B(n_1625),
.C(n_1552),
.D(n_1605),
.Y(n_1846)
);

AOI211xp5_ASAP7_75t_L g1847 ( 
.A1(n_1841),
.A2(n_1512),
.B(n_1736),
.C(n_1735),
.Y(n_1847)
);

AOI221xp5_ASAP7_75t_L g1848 ( 
.A1(n_1835),
.A2(n_1736),
.B1(n_1731),
.B2(n_1728),
.C(n_1725),
.Y(n_1848)
);

NAND3xp33_ASAP7_75t_SL g1849 ( 
.A(n_1839),
.B(n_1740),
.C(n_1711),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1837),
.B(n_1840),
.Y(n_1850)
);

AOI221xp5_ASAP7_75t_L g1851 ( 
.A1(n_1846),
.A2(n_1740),
.B1(n_1711),
.B2(n_1688),
.C(n_1668),
.Y(n_1851)
);

OAI221xp5_ASAP7_75t_L g1852 ( 
.A1(n_1836),
.A2(n_1605),
.B1(n_1589),
.B2(n_1679),
.C(n_1609),
.Y(n_1852)
);

AOI31xp33_ASAP7_75t_L g1853 ( 
.A1(n_1843),
.A2(n_1546),
.A3(n_1548),
.B(n_1556),
.Y(n_1853)
);

OAI311xp33_ASAP7_75t_L g1854 ( 
.A1(n_1848),
.A2(n_1838),
.A3(n_1850),
.B1(n_1852),
.C1(n_1851),
.Y(n_1854)
);

AOI221xp5_ASAP7_75t_L g1855 ( 
.A1(n_1849),
.A2(n_1844),
.B1(n_1842),
.B2(n_1845),
.C(n_1664),
.Y(n_1855)
);

OAI22xp5_ASAP7_75t_L g1856 ( 
.A1(n_1847),
.A2(n_1632),
.B1(n_1662),
.B2(n_1671),
.Y(n_1856)
);

AOI32xp33_ASAP7_75t_L g1857 ( 
.A1(n_1853),
.A2(n_1694),
.A3(n_1690),
.B1(n_1687),
.B2(n_1686),
.Y(n_1857)
);

AOI211xp5_ASAP7_75t_L g1858 ( 
.A1(n_1849),
.A2(n_1538),
.B(n_1548),
.C(n_1546),
.Y(n_1858)
);

OAI221xp5_ASAP7_75t_L g1859 ( 
.A1(n_1847),
.A2(n_1679),
.B1(n_1609),
.B2(n_1668),
.C(n_1664),
.Y(n_1859)
);

AOI21xp33_ASAP7_75t_SL g1860 ( 
.A1(n_1850),
.A2(n_1538),
.B(n_1682),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1859),
.Y(n_1861)
);

NAND4xp75_ASAP7_75t_L g1862 ( 
.A(n_1855),
.B(n_1680),
.C(n_1667),
.D(n_1674),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1858),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1856),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1860),
.Y(n_1865)
);

AND4x1_ASAP7_75t_L g1866 ( 
.A(n_1864),
.B(n_1854),
.C(n_1857),
.D(n_1558),
.Y(n_1866)
);

CKINVDCx12_ASAP7_75t_R g1867 ( 
.A(n_1861),
.Y(n_1867)
);

NAND3xp33_ASAP7_75t_L g1868 ( 
.A(n_1865),
.B(n_1682),
.C(n_1677),
.Y(n_1868)
);

OAI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1868),
.A2(n_1863),
.B1(n_1862),
.B2(n_1668),
.Y(n_1869)
);

OAI22x1_ASAP7_75t_L g1870 ( 
.A1(n_1869),
.A2(n_1866),
.B1(n_1867),
.B2(n_1862),
.Y(n_1870)
);

OAI22xp5_ASAP7_75t_L g1871 ( 
.A1(n_1870),
.A2(n_1677),
.B1(n_1682),
.B2(n_1668),
.Y(n_1871)
);

AOI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1870),
.A2(n_1548),
.B1(n_1546),
.B2(n_1677),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1872),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1871),
.Y(n_1874)
);

AOI22xp33_ASAP7_75t_L g1875 ( 
.A1(n_1873),
.A2(n_1677),
.B1(n_1682),
.B2(n_1556),
.Y(n_1875)
);

OAI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1874),
.A2(n_1537),
.B(n_1667),
.Y(n_1876)
);

AOI22xp5_ASAP7_75t_L g1877 ( 
.A1(n_1875),
.A2(n_1876),
.B1(n_1667),
.B2(n_1674),
.Y(n_1877)
);

OA21x2_ASAP7_75t_L g1878 ( 
.A1(n_1877),
.A2(n_1684),
.B(n_1674),
.Y(n_1878)
);

XOR2xp5_ASAP7_75t_L g1879 ( 
.A(n_1878),
.B(n_1540),
.Y(n_1879)
);

OAI221xp5_ASAP7_75t_R g1880 ( 
.A1(n_1879),
.A2(n_1540),
.B1(n_1680),
.B2(n_1684),
.C(n_1671),
.Y(n_1880)
);

AOI211xp5_ASAP7_75t_L g1881 ( 
.A1(n_1880),
.A2(n_1680),
.B(n_1684),
.C(n_1537),
.Y(n_1881)
);


endmodule