module real_jpeg_6695_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_0),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_0),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_0),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_0),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_0),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_0),
.B(n_289),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_0),
.B(n_118),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_0),
.B(n_428),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_1),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_1),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_1),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_1),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_1),
.B(n_171),
.Y(n_170)
);

AND2x2_ASAP7_75t_SL g196 ( 
.A(n_1),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_1),
.B(n_199),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_1),
.B(n_234),
.Y(n_233)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_2),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g278 ( 
.A(n_2),
.Y(n_278)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_2),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_2),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_2),
.Y(n_385)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_3),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_3),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_4),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_5),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_5),
.B(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_5),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_5),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_5),
.B(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_5),
.B(n_177),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_5),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_6),
.B(n_114),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_6),
.B(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_6),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_6),
.B(n_307),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_6),
.B(n_341),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_6),
.B(n_289),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_6),
.B(n_421),
.Y(n_420)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_7),
.Y(n_115)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_7),
.Y(n_246)
);

BUFx5_ASAP7_75t_L g412 ( 
.A(n_7),
.Y(n_412)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_9),
.Y(n_121)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_9),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g382 ( 
.A(n_9),
.Y(n_382)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_11),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_11),
.Y(n_290)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_13),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_13),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_13),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_13),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_13),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_13),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_13),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_13),
.B(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_14),
.B(n_49),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_14),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_14),
.B(n_321),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_14),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_14),
.B(n_363),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_14),
.B(n_105),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_14),
.B(n_408),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_15),
.B(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_15),
.B(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_15),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_15),
.B(n_350),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_15),
.B(n_232),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_15),
.B(n_33),
.Y(n_397)
);

AND2x6_ASAP7_75t_SL g411 ( 
.A(n_15),
.B(n_412),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_16),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_16),
.B(n_203),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_16),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_16),
.B(n_47),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_16),
.B(n_304),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_16),
.B(n_323),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_16),
.B(n_388),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_16),
.B(n_382),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_17),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_17),
.B(n_98),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_17),
.B(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_17),
.B(n_323),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_17),
.B(n_289),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_17),
.B(n_369),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_17),
.B(n_225),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_17),
.B(n_232),
.Y(n_418)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_19),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_19),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_19),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_19),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_19),
.B(n_228),
.Y(n_227)
);

AND2x2_ASAP7_75t_SL g301 ( 
.A(n_19),
.B(n_120),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_19),
.B(n_385),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_19),
.B(n_426),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_23),
.B(n_537),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx13_ASAP7_75t_L g539 ( 
.A(n_22),
.Y(n_539)
);

O2A1O1Ixp33_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_45),
.B(n_80),
.C(n_536),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_50),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_26),
.B(n_50),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_43),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_32),
.C(n_36),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_28),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_28),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_28),
.A2(n_32),
.B1(n_44),
.B2(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_30),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_32),
.A2(n_54),
.B1(n_59),
.B2(n_60),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_32),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_32),
.B(n_54),
.C(n_61),
.Y(n_77)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_34),
.Y(n_282)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_35),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_35),
.Y(n_308)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_35),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_36),
.B(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_76),
.C(n_78),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_51),
.B(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_63),
.C(n_68),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_52),
.B(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_61),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_54),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_54),
.A2(n_60),
.B1(n_72),
.B2(n_122),
.Y(n_126)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_57),
.Y(n_220)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_58),
.Y(n_150)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_58),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_69),
.C(n_72),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_63),
.B(n_68),
.Y(n_129)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_69),
.A2(n_70),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_72),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_72),
.A2(n_116),
.B1(n_117),
.B2(n_122),
.Y(n_509)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_75),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g235 ( 
.A(n_75),
.Y(n_235)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_75),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_76),
.A2(n_77),
.B1(n_78),
.B2(n_132),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

AO21x1_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_133),
.B(n_535),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_130),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_82),
.B(n_130),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_127),
.C(n_128),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_83),
.A2(n_84),
.B1(n_531),
.B2(n_532),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_110),
.C(n_123),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_85),
.A2(n_86),
.B1(n_513),
.B2(n_515),
.Y(n_512)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_96),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_91),
.C(n_96),
.Y(n_127)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_94),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_101),
.C(n_106),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_97),
.B(n_504),
.Y(n_503)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_99),
.Y(n_182)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_101),
.A2(n_102),
.B1(n_106),
.B2(n_107),
.Y(n_504)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_104),
.B(n_292),
.Y(n_291)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_109),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_110),
.A2(n_123),
.B1(n_124),
.B2(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_110),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_116),
.C(n_122),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g508 ( 
.A(n_111),
.B(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_115),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_116),
.A2(n_117),
.B1(n_212),
.B2(n_215),
.Y(n_211)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_117),
.B(n_208),
.C(n_212),
.Y(n_510)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx5_ASAP7_75t_L g347 ( 
.A(n_121),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_121),
.Y(n_370)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g532 ( 
.A(n_127),
.B(n_128),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_529),
.B(n_534),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_497),
.B(n_526),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_309),
.B(n_496),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_263),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_137),
.B(n_263),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_205),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_138),
.B(n_206),
.C(n_238),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_179),
.C(n_189),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_139),
.B(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_152),
.C(n_166),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_140),
.B(n_482),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_146),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_141),
.B(n_147),
.C(n_151),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_145),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_145),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_152),
.A2(n_153),
.B1(n_166),
.B2(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.C(n_162),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_154),
.B(n_162),
.Y(n_472)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_157),
.B(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx5_ASAP7_75t_L g365 ( 
.A(n_161),
.Y(n_365)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_161),
.Y(n_421)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_166),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_167),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_175),
.B2(n_176),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_170),
.B(n_175),
.C(n_249),
.Y(n_248)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_174),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_174),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_174),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_175),
.A2(n_176),
.B1(n_212),
.B2(n_215),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_175),
.B(n_212),
.C(n_242),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_178),
.Y(n_332)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_178),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_179),
.B(n_189),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_188),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_183),
.B1(n_186),
.B2(n_187),
.Y(n_180)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_181),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_183),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_183),
.A2(n_187),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_183),
.B(n_186),
.C(n_262),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_183),
.B(n_255),
.C(n_259),
.Y(n_505)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_188),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_198),
.C(n_202),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_190),
.B(n_295),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.C(n_196),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_191),
.B(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_193),
.B(n_196),
.Y(n_275)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_198),
.B(n_202),
.Y(n_295)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_201),
.Y(n_327)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_238),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_216),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_207),
.B(n_217),
.C(n_237),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_212),
.Y(n_215)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_214),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_226),
.B1(n_236),
.B2(n_237),
.Y(n_216)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_217),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.C(n_222),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_222),
.Y(n_251)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_226),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_230),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_227),
.B(n_231),
.C(n_233),
.Y(n_511)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_252),
.B2(n_253),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_239),
.B(n_254),
.C(n_261),
.Y(n_522)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_248),
.C(n_250),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_241),
.B(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_247),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_250),
.Y(n_269)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_261),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_257),
.B2(n_258),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_259),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_267),
.C(n_270),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_265),
.B(n_268),
.Y(n_492)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_270),
.B(n_492),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_293),
.C(n_296),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_272),
.B(n_485),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_276),
.C(n_283),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_273),
.A2(n_274),
.B1(n_463),
.B2(n_464),
.Y(n_462)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_276),
.A2(n_277),
.B(n_279),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_276),
.B(n_283),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

MAJx2_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_287),
.C(n_291),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_284),
.A2(n_285),
.B1(n_287),
.B2(n_288),
.Y(n_440)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx8_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_291),
.B(n_440),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_292),
.B(n_381),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_L g485 ( 
.A1(n_293),
.A2(n_294),
.B1(n_296),
.B2(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_296),
.Y(n_486)
);

MAJx2_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_305),
.C(n_306),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_298),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_298),
.B(n_474),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.C(n_302),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_299),
.B(n_452),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_301),
.A2(n_302),
.B1(n_303),
.B2(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_301),
.Y(n_453)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_305),
.B(n_306),
.Y(n_474)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

AOI21x1_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_490),
.B(n_495),
.Y(n_309)
);

OAI21x1_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_477),
.B(n_489),
.Y(n_310)
);

AOI21x1_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_459),
.B(n_476),
.Y(n_311)
);

OAI21x1_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_433),
.B(n_458),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_314),
.A2(n_402),
.B(n_432),
.Y(n_313)
);

OAI21x1_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_373),
.B(n_401),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_354),
.B(n_372),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_334),
.B(n_353),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_328),
.B(n_333),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_325),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_319),
.B(n_325),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_322),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_329),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_320),
.B(n_322),
.Y(n_335)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_336),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_337),
.A2(n_338),
.B1(n_342),
.B2(n_343),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_337),
.B(n_345),
.C(n_348),
.Y(n_371)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_339),
.B(n_340),
.Y(n_360)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_344),
.A2(n_345),
.B1(n_348),
.B2(n_349),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_355),
.B(n_371),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_355),
.B(n_371),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_361),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_360),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_357),
.B(n_360),
.C(n_375),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_358),
.B(n_359),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_361),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_366),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_362),
.B(n_392),
.C(n_393),
.Y(n_391)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_368),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_367),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_368),
.Y(n_393)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_376),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_374),
.B(n_376),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_390),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_377),
.B(n_391),
.C(n_394),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_378),
.B(n_380),
.C(n_383),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_383),
.Y(n_379)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_384),
.A2(n_386),
.B1(n_387),
.B2(n_389),
.Y(n_383)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_384),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_386),
.B(n_389),
.Y(n_413)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_394),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_396),
.Y(n_394)
);

MAJx2_ASAP7_75t_L g430 ( 
.A(n_395),
.B(n_398),
.C(n_399),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_397),
.A2(n_398),
.B1(n_399),
.B2(n_400),
.Y(n_396)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_397),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_398),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_403),
.B(n_431),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_403),
.B(n_431),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_404),
.B(n_415),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_414),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_405),
.B(n_414),
.C(n_457),
.Y(n_456)
);

XNOR2x1_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_413),
.Y(n_405)
);

XNOR2x1_ASAP7_75t_SL g406 ( 
.A(n_407),
.B(n_411),
.Y(n_406)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_407),
.Y(n_447)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx6_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

CKINVDCx14_ASAP7_75t_R g448 ( 
.A(n_411),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_413),
.B(n_447),
.C(n_448),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_415),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_422),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_416),
.B(n_424),
.C(n_429),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_420),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_419),
.Y(n_417)
);

MAJx2_ASAP7_75t_L g444 ( 
.A(n_418),
.B(n_419),
.C(n_420),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_424),
.B1(n_429),
.B2(n_430),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_427),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_425),
.B(n_427),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_430),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_434),
.B(n_456),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_434),
.B(n_456),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_445),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_437),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_436),
.B(n_437),
.C(n_445),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_438),
.A2(n_439),
.B1(n_441),
.B2(n_442),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_438),
.B(n_468),
.C(n_469),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_444),
.Y(n_442)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_443),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_444),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_446),
.B(n_449),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_446),
.B(n_450),
.C(n_455),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_450),
.A2(n_451),
.B1(n_454),
.B2(n_455),
.Y(n_449)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_450),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_451),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_460),
.B(n_475),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_460),
.B(n_475),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_SL g460 ( 
.A(n_461),
.B(n_466),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_465),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_462),
.B(n_465),
.C(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_463),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_466),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_467),
.B(n_470),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_467),
.B(n_471),
.C(n_473),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_473),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_478),
.B(n_487),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_478),
.B(n_487),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_480),
.Y(n_478)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_479),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_484),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_481),
.B(n_484),
.C(n_494),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_491),
.B(n_493),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_491),
.B(n_493),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_523),
.Y(n_497)
);

OAI21xp33_ASAP7_75t_L g526 ( 
.A1(n_498),
.A2(n_527),
.B(n_528),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_499),
.B(n_517),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_499),
.B(n_517),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_500),
.A2(n_501),
.B1(n_506),
.B2(n_516),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_500),
.B(n_507),
.C(n_512),
.Y(n_533)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_503),
.C(n_505),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_502),
.B(n_519),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_503),
.B(n_505),
.Y(n_519)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_506),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_512),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_510),
.C(n_511),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_508),
.B(n_521),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_510),
.B(n_511),
.Y(n_521)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_513),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_518),
.B(n_520),
.C(n_522),
.Y(n_517)
);

FAx1_ASAP7_75t_SL g524 ( 
.A(n_518),
.B(n_520),
.CI(n_522),
.CON(n_524),
.SN(n_524)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_524),
.B(n_525),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_524),
.B(n_525),
.Y(n_527)
);

BUFx24_ASAP7_75t_SL g541 ( 
.A(n_524),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_SL g529 ( 
.A(n_530),
.B(n_533),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_530),
.B(n_533),
.Y(n_534)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_538),
.B(n_540),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);


endmodule