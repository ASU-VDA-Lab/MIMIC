module fake_jpeg_24422_n_179 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_35),
.B(n_38),
.Y(n_44)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_0),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_1),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

NOR2x1_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_25),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_51),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_31),
.B1(n_22),
.B2(n_25),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_52),
.B1(n_54),
.B2(n_40),
.Y(n_63)
);

NOR2x1_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_25),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_32),
.A2(n_31),
.B1(n_40),
.B2(n_22),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_32),
.A2(n_31),
.B1(n_25),
.B2(n_27),
.Y(n_54)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_59),
.B(n_23),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_29),
.B1(n_27),
.B2(n_20),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_62),
.A2(n_63),
.B1(n_29),
.B2(n_15),
.Y(n_87)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_68),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_66),
.B(n_71),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_67),
.Y(n_99)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVxp67_ASAP7_75t_SL g85 ( 
.A(n_69),
.Y(n_85)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_72),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_56),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_53),
.Y(n_73)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_21),
.Y(n_75)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_77),
.Y(n_94)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_21),
.Y(n_78)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_48),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_49),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_45),
.C(n_44),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_84),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_70),
.B(n_59),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_96),
.B1(n_98),
.B2(n_67),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_80),
.A2(n_72),
.B1(n_71),
.B2(n_63),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_91),
.A2(n_76),
.B1(n_68),
.B2(n_64),
.Y(n_107)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_45),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_93),
.B(n_65),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_33),
.B1(n_42),
.B2(n_50),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_74),
.A2(n_33),
.B1(n_36),
.B2(n_54),
.Y(n_98)
);

OA21x2_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_20),
.B(n_49),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_99),
.B(n_101),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_84),
.B(n_34),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_90),
.C(n_97),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_67),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_105),
.B(n_109),
.Y(n_127)
);

NOR3xp33_ASAP7_75t_SL g106 ( 
.A(n_86),
.B(n_28),
.C(n_26),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_114),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_107),
.A2(n_100),
.B(n_83),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_89),
.B(n_23),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_101),
.A2(n_81),
.B1(n_77),
.B2(n_79),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_110),
.A2(n_98),
.B1(n_96),
.B2(n_92),
.Y(n_120)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_111),
.B(n_2),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_119),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_113),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_15),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_115),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_28),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_117),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_26),
.Y(n_118)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_118),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_82),
.B(n_1),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_120),
.A2(n_124),
.B1(n_129),
.B2(n_131),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_126),
.B1(n_110),
.B2(n_109),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_87),
.B1(n_82),
.B2(n_100),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_103),
.Y(n_125)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_90),
.B1(n_69),
.B2(n_43),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_108),
.Y(n_136)
);

AO22x1_ASAP7_75t_SL g131 ( 
.A1(n_102),
.A2(n_107),
.B1(n_113),
.B2(n_104),
.Y(n_131)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_142),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_115),
.Y(n_138)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_135),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_141),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_108),
.C(n_112),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_127),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_144),
.A2(n_121),
.B(n_133),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_145),
.A2(n_147),
.B(n_131),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_121),
.B(n_119),
.Y(n_146)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_146),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_106),
.B1(n_115),
.B2(n_16),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_149),
.A2(n_151),
.B(n_153),
.Y(n_158)
);

OAI321xp33_ASAP7_75t_L g150 ( 
.A1(n_137),
.A2(n_131),
.A3(n_124),
.B1(n_126),
.B2(n_125),
.C(n_120),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_156),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_139),
.B(n_131),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_129),
.B(n_132),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_156),
.A2(n_139),
.B1(n_142),
.B2(n_143),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_160),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_154),
.A2(n_143),
.B1(n_134),
.B2(n_136),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_148),
.A2(n_122),
.B1(n_13),
.B2(n_12),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_162),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_122),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_34),
.C(n_18),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_2),
.Y(n_168)
);

OAI322xp33_ASAP7_75t_L g164 ( 
.A1(n_159),
.A2(n_152),
.A3(n_16),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_167),
.B(n_18),
.Y(n_169)
);

OAI322xp33_ASAP7_75t_L g167 ( 
.A1(n_160),
.A2(n_157),
.A3(n_158),
.B1(n_163),
.B2(n_161),
.C1(n_34),
.C2(n_18),
.Y(n_167)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_168),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_170),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_165),
.A2(n_157),
.B(n_4),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_164),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_166),
.B1(n_6),
.B2(n_7),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_173),
.A2(n_7),
.B(n_8),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_5),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_175),
.A2(n_9),
.B(n_174),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_177),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_178),
.B(n_173),
.Y(n_179)
);


endmodule