module real_jpeg_23708_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_0),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_1),
.B(n_37),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_2),
.B(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_2),
.B(n_23),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_2),
.B(n_32),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_3),
.B(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_3),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_3),
.B(n_32),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_3),
.B(n_29),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_6),
.B(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_6),
.B(n_23),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_6),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_6),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_7),
.B(n_19),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_7),
.B(n_23),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_10),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_10),
.B(n_23),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_10),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_10),
.B(n_29),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_10),
.B(n_67),
.Y(n_80)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_72),
.Y(n_12)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_51),
.C(n_52),
.Y(n_13)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_34),
.C(n_41),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_17),
.B1(n_26),
.B2(n_27),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_16),
.B(n_28),
.C(n_31),
.Y(n_51)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_21),
.B1(n_22),
.B2(n_25),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_21),
.B(n_25),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_39),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_36),
.B1(n_39),
.B2(n_40),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.C(n_46),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_62),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_57),
.C(n_62),
.Y(n_73)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_58),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_59),
.B(n_61),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_65),
.B2(n_71),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_63),
.Y(n_71)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_66),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_70),
.C(n_71),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_85),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_90),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);


endmodule