module fake_netlist_1_4326_n_12 (n_1, n_2, n_0, n_12);
input n_1;
input n_2;
input n_0;
output n_12;
wire n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx1_ASAP7_75t_L g3 ( .A(n_2), .Y(n_3) );
INVx2_ASAP7_75t_L g4 ( .A(n_1), .Y(n_4) );
OAI22xp5_ASAP7_75t_L g5 ( .A1(n_3), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_5) );
OAI21x1_ASAP7_75t_L g6 ( .A1(n_4), .A2(n_0), .B(n_1), .Y(n_6) );
CKINVDCx20_ASAP7_75t_R g7 ( .A(n_5), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
O2A1O1Ixp5_ASAP7_75t_L g9 ( .A1(n_8), .A2(n_4), .B(n_6), .C(n_2), .Y(n_9) );
OAI31xp33_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_8), .A3(n_1), .B(n_2), .Y(n_10) );
OAI21xp5_ASAP7_75t_L g11 ( .A1(n_10), .A2(n_9), .B(n_6), .Y(n_11) );
AOI22xp5_ASAP7_75t_SL g12 ( .A1(n_11), .A2(n_0), .B1(n_10), .B2(n_7), .Y(n_12) );
endmodule