module fake_jpeg_30623_n_421 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_421);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_421;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx3_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_12),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_45),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_7),
.B(n_13),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_44),
.C(n_32),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_21),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_48),
.B(n_51),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_8),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_71),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_22),
.B(n_8),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_52),
.B(n_57),
.Y(n_106)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_56),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_22),
.B(n_8),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_21),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_58),
.B(n_59),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_21),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_21),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_60),
.B(n_63),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_21),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_65),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_33),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_67),
.B(n_69),
.Y(n_129)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_33),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_70),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_19),
.B(n_6),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_33),
.B(n_6),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_76),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_73),
.Y(n_139)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_33),
.B(n_9),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_78),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_33),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_81),
.B(n_83),
.Y(n_90)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_19),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_19),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_84),
.B(n_85),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_30),
.B(n_9),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_86),
.A2(n_87),
.B1(n_42),
.B2(n_35),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_88),
.B(n_44),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_46),
.A2(n_36),
.B1(n_25),
.B2(n_34),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_89),
.A2(n_100),
.B1(n_103),
.B2(n_113),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_94),
.B(n_98),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_96),
.A2(n_131),
.B1(n_61),
.B2(n_78),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_65),
.A2(n_28),
.B1(n_17),
.B2(n_25),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_97),
.A2(n_108),
.B1(n_114),
.B2(n_116),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_50),
.A2(n_25),
.B1(n_34),
.B2(n_31),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_64),
.A2(n_39),
.B1(n_32),
.B2(n_27),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_47),
.A2(n_17),
.B1(n_28),
.B2(n_86),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_72),
.B(n_31),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_112),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_26),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_56),
.A2(n_26),
.B1(n_43),
.B2(n_41),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_62),
.A2(n_28),
.B1(n_17),
.B2(n_42),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_88),
.A2(n_43),
.B1(n_41),
.B2(n_30),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_66),
.A2(n_28),
.B1(n_39),
.B2(n_23),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_117),
.A2(n_123),
.B1(n_124),
.B2(n_127),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_71),
.B(n_45),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_133),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_73),
.A2(n_28),
.B1(n_80),
.B2(n_87),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_54),
.A2(n_23),
.B1(n_35),
.B2(n_19),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_77),
.A2(n_79),
.B1(n_81),
.B2(n_58),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_48),
.A2(n_23),
.B1(n_35),
.B2(n_40),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_71),
.B(n_74),
.Y(n_133)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_140),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_105),
.B(n_70),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_141),
.B(n_160),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_143),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_99),
.B(n_84),
.C(n_83),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_144),
.B(n_115),
.C(n_134),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_129),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_145),
.B(n_151),
.Y(n_207)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_146),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_147),
.A2(n_117),
.B1(n_115),
.B2(n_126),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_149),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_118),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_106),
.B(n_138),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_152),
.B(n_162),
.Y(n_214)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_154),
.Y(n_226)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_155),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_99),
.B(n_67),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_157),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_112),
.B(n_59),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_93),
.B(n_60),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_158),
.B(n_172),
.Y(n_208)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_159),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_109),
.B(n_63),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_68),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_90),
.B(n_53),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_163),
.B(n_164),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_120),
.B(n_78),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_133),
.B(n_78),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_166),
.B(n_168),
.Y(n_223)
);

A2O1A1O1Ixp25_ASAP7_75t_L g167 ( 
.A1(n_89),
.A2(n_61),
.B(n_75),
.C(n_82),
.D(n_49),
.Y(n_167)
);

A2O1A1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_167),
.A2(n_52),
.B(n_40),
.C(n_137),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_121),
.B(n_61),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_102),
.Y(n_170)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_170),
.Y(n_210)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_171),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_93),
.B(n_23),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_174),
.Y(n_216)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_121),
.Y(n_175)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_175),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_101),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_104),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_177),
.B(n_181),
.Y(n_224)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_104),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_178),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_100),
.A2(n_55),
.B1(n_23),
.B2(n_3),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_179),
.A2(n_135),
.B1(n_130),
.B2(n_125),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_93),
.B(n_11),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_180),
.B(n_13),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_94),
.B(n_132),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_91),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_182),
.B(n_186),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_111),
.A2(n_40),
.B1(n_52),
.B2(n_3),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_183),
.A2(n_125),
.B1(n_139),
.B2(n_128),
.Y(n_189)
);

BUFx24_ASAP7_75t_L g185 ( 
.A(n_110),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_185),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_116),
.Y(n_186)
);

OAI21xp33_ASAP7_75t_L g259 ( 
.A1(n_189),
.A2(n_176),
.B(n_154),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_173),
.B(n_156),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_190),
.B(n_202),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_184),
.A2(n_98),
.B1(n_139),
.B2(n_128),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_191),
.A2(n_193),
.B1(n_201),
.B2(n_219),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_111),
.B(n_113),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_196),
.A2(n_199),
.B(n_164),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_184),
.A2(n_136),
.B1(n_130),
.B2(n_135),
.Y(n_201)
);

MAJx2_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_126),
.C(n_95),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_148),
.B(n_95),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_203),
.B(n_206),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_136),
.B1(n_135),
.B2(n_134),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_213),
.A2(n_140),
.B1(n_161),
.B2(n_169),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_218),
.B(n_220),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_157),
.A2(n_136),
.B1(n_110),
.B2(n_137),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_187),
.B(n_142),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_227),
.B(n_238),
.Y(n_266)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_228),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_225),
.A2(n_153),
.B1(n_150),
.B2(n_175),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_229),
.A2(n_255),
.B1(n_213),
.B2(n_222),
.Y(n_267)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_192),
.Y(n_230)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_230),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_232),
.A2(n_234),
.B1(n_242),
.B2(n_212),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_233),
.A2(n_241),
.B(n_215),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_187),
.A2(n_196),
.B1(n_199),
.B2(n_191),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_195),
.Y(n_235)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_235),
.Y(n_277)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_237),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_142),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_190),
.B(n_208),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_239),
.B(n_247),
.Y(n_284)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_197),
.Y(n_240)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_240),
.Y(n_273)
);

NAND2xp33_ASAP7_75t_SL g241 ( 
.A(n_208),
.B(n_158),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_224),
.A2(n_144),
.B1(n_167),
.B2(n_148),
.Y(n_242)
);

O2A1O1Ixp33_ASAP7_75t_L g243 ( 
.A1(n_188),
.A2(n_151),
.B(n_174),
.C(n_180),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_243),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_207),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_245),
.B(n_246),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_145),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_206),
.B(n_160),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_194),
.B(n_141),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_252),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_195),
.B(n_172),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_251),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_205),
.Y(n_250)
);

INVx13_ASAP7_75t_L g292 ( 
.A(n_250),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_165),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_194),
.B(n_223),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_218),
.B(n_165),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_253),
.B(n_198),
.Y(n_282)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_200),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_254),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_201),
.A2(n_178),
.B1(n_177),
.B2(n_171),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_222),
.B(n_165),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_257),
.Y(n_268)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_197),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_155),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_221),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_259),
.A2(n_261),
.B1(n_210),
.B2(n_209),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_205),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_260),
.B(n_202),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_263),
.B(n_281),
.C(n_244),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_267),
.A2(n_269),
.B1(n_278),
.B2(n_285),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_231),
.A2(n_220),
.B1(n_193),
.B2(n_212),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_270),
.A2(n_40),
.B(n_11),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_245),
.B(n_188),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_272),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_276),
.A2(n_279),
.B1(n_286),
.B2(n_287),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_231),
.A2(n_216),
.B1(n_200),
.B2(n_149),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_234),
.A2(n_216),
.B1(n_226),
.B2(n_211),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_204),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_280),
.B(n_288),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_185),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_282),
.B(n_290),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_247),
.A2(n_170),
.B1(n_226),
.B2(n_198),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_233),
.A2(n_204),
.B1(n_210),
.B2(n_209),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_255),
.A2(n_209),
.B1(n_215),
.B2(n_146),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_232),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_267),
.A2(n_242),
.B1(n_243),
.B2(n_235),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_293),
.A2(n_294),
.B(n_296),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_230),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_269),
.A2(n_228),
.B1(n_236),
.B2(n_254),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_253),
.Y(n_297)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_297),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_298),
.B(n_308),
.C(n_311),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_263),
.B(n_244),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_301),
.B(n_303),
.Y(n_323)
);

OR2x6_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_241),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_302),
.A2(n_310),
.B(n_276),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_284),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_264),
.Y(n_304)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_304),
.Y(n_336)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_264),
.Y(n_305)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_265),
.B(n_227),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_306),
.B(n_315),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_284),
.B(n_239),
.Y(n_308)
);

OA21x2_ASAP7_75t_L g310 ( 
.A1(n_283),
.A2(n_249),
.B(n_238),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_266),
.B(n_240),
.C(n_257),
.Y(n_311)
);

XNOR2x1_ASAP7_75t_L g312 ( 
.A(n_266),
.B(n_282),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_312),
.B(n_313),
.Y(n_332)
);

MAJx2_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_185),
.C(n_237),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_262),
.B(n_261),
.C(n_250),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_314),
.B(n_317),
.C(n_285),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_289),
.B(n_159),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_286),
.B(n_261),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_316),
.A2(n_319),
.B(n_273),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_262),
.B(n_250),
.C(n_185),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_288),
.A2(n_11),
.B1(n_14),
.B2(n_4),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_318),
.A2(n_268),
.B1(n_277),
.B2(n_275),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_300),
.B(n_274),
.Y(n_320)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_320),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_321),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_309),
.Y(n_325)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_325),
.Y(n_356)
);

NOR2x1_ASAP7_75t_L g326 ( 
.A(n_302),
.B(n_279),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_326),
.B(n_302),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_295),
.A2(n_316),
.B1(n_278),
.B2(n_294),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_327),
.A2(n_299),
.B1(n_293),
.B2(n_296),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_329),
.B(n_331),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_298),
.B(n_301),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_330),
.B(n_338),
.Y(n_346)
);

AOI21xp33_ASAP7_75t_L g331 ( 
.A1(n_302),
.A2(n_277),
.B(n_275),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_313),
.Y(n_333)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_333),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_311),
.B(n_274),
.Y(n_337)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_337),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_303),
.B(n_291),
.C(n_287),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_339),
.B(n_341),
.C(n_299),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_340),
.A2(n_273),
.B(n_292),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_314),
.B(n_307),
.C(n_317),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_312),
.B(n_291),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_342),
.B(n_308),
.Y(n_348)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_344),
.Y(n_364)
);

FAx1_ASAP7_75t_SL g347 ( 
.A(n_321),
.B(n_307),
.CI(n_302),
.CON(n_347),
.SN(n_347)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_347),
.B(n_332),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_348),
.B(n_353),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_334),
.B(n_310),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_349),
.B(n_358),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_352),
.A2(n_326),
.B1(n_360),
.B2(n_328),
.Y(n_368)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_320),
.Y(n_354)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_354),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_330),
.B(n_310),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_355),
.B(n_357),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_335),
.B(n_292),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_324),
.B(n_292),
.C(n_2),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_359),
.B(n_362),
.C(n_341),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_339),
.B(n_4),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_361),
.B(n_322),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_324),
.B(n_1),
.C(n_2),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_343),
.A2(n_333),
.B1(n_328),
.B2(n_327),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_363),
.B(n_371),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_345),
.B(n_337),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_365),
.B(n_368),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_356),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_366),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_370),
.A2(n_377),
.B(n_357),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_352),
.A2(n_340),
.B1(n_332),
.B2(n_342),
.Y(n_371)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_372),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_373),
.B(n_376),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_360),
.A2(n_338),
.B1(n_322),
.B2(n_336),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_351),
.A2(n_323),
.B1(n_1),
.B2(n_5),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_374),
.B(n_346),
.C(n_353),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_378),
.B(n_381),
.C(n_383),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_369),
.B(n_343),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_379),
.B(n_368),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_380),
.B(n_389),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_374),
.B(n_346),
.C(n_351),
.Y(n_381)
);

OAI21x1_ASAP7_75t_SL g382 ( 
.A1(n_364),
.A2(n_344),
.B(n_347),
.Y(n_382)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_382),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_376),
.B(n_355),
.C(n_359),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_375),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_387),
.B(n_366),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_388),
.A2(n_367),
.B(n_363),
.Y(n_390)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_390),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_391),
.B(n_393),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_384),
.B(n_356),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_389),
.A2(n_350),
.B1(n_354),
.B2(n_367),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_394),
.B(n_397),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_386),
.B(n_377),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_395),
.B(n_396),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_378),
.B(n_373),
.C(n_371),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_398),
.B(n_381),
.C(n_385),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_400),
.B(n_404),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_399),
.A2(n_385),
.B(n_383),
.Y(n_403)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_403),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_394),
.A2(n_370),
.B1(n_362),
.B2(n_347),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_392),
.B(n_323),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_406),
.B(n_4),
.C(n_5),
.Y(n_409)
);

A2O1A1O1Ixp25_ASAP7_75t_L g408 ( 
.A1(n_401),
.A2(n_392),
.B(n_398),
.C(n_397),
.D(n_348),
.Y(n_408)
);

O2A1O1Ixp33_ASAP7_75t_SL g415 ( 
.A1(n_408),
.A2(n_411),
.B(n_407),
.C(n_400),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_409),
.B(n_405),
.Y(n_414)
);

O2A1O1Ixp33_ASAP7_75t_SL g411 ( 
.A1(n_402),
.A2(n_14),
.B(n_5),
.C(n_12),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_410),
.Y(n_413)
);

OAI21x1_ASAP7_75t_L g417 ( 
.A1(n_413),
.A2(n_415),
.B(n_407),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_414),
.Y(n_416)
);

O2A1O1Ixp33_ASAP7_75t_SL g418 ( 
.A1(n_417),
.A2(n_412),
.B(n_12),
.C(n_13),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_418),
.B(n_416),
.Y(n_419)
);

NOR3xp33_ASAP7_75t_L g420 ( 
.A(n_419),
.B(n_13),
.C(n_14),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_420),
.B(n_1),
.Y(n_421)
);


endmodule