module real_jpeg_25711_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_173;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_113;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_1),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_2),
.A2(n_25),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_4),
.A2(n_37),
.B1(n_38),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_4),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_4),
.A2(n_52),
.B1(n_53),
.B2(n_59),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_4),
.A2(n_25),
.B1(n_31),
.B2(n_59),
.Y(n_160)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_6),
.A2(n_25),
.B1(n_31),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_9),
.A2(n_37),
.B1(n_38),
.B2(n_62),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_9),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_9),
.A2(n_52),
.B1(n_53),
.B2(n_62),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_9),
.A2(n_47),
.B1(n_62),
.B2(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_9),
.A2(n_25),
.B1(n_31),
.B2(n_62),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_10),
.A2(n_37),
.B1(n_38),
.B2(n_81),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_10),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_10),
.A2(n_52),
.B1(n_53),
.B2(n_81),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_10),
.A2(n_25),
.B1(n_31),
.B2(n_81),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_11),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_11),
.B(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_11),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_11),
.B(n_53),
.C(n_55),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_11),
.A2(n_37),
.B1(n_38),
.B2(n_97),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_11),
.B(n_79),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_11),
.A2(n_52),
.B1(n_53),
.B2(n_97),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_11),
.B(n_25),
.C(n_87),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_11),
.A2(n_24),
.B(n_148),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_13),
.A2(n_25),
.B1(n_31),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_13),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_13),
.A2(n_52),
.B1(n_53),
.B2(n_71),
.Y(n_84)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_14),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_14),
.B(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_14),
.Y(n_162)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_14),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_123),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_121),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_103),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_18),
.B(n_103),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_74),
.B2(n_75),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_49),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_36),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_23),
.A2(n_159),
.B1(n_161),
.B2(n_163),
.Y(n_158)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_24),
.A2(n_30),
.B1(n_70),
.B2(n_72),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_24),
.B(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_24),
.A2(n_147),
.B(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_25),
.A2(n_31),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_31),
.B(n_173),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_33),
.A2(n_118),
.B(n_119),
.Y(n_117)
);

AOI32xp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.A3(n_43),
.B1(n_45),
.B2(n_48),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_37),
.A2(n_38),
.B1(n_55),
.B2(n_56),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_37),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_68)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp33_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_44),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_38),
.B(n_116),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp33_ASAP7_75t_L g96 ( 
.A1(n_41),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_42),
.A2(n_43),
.B1(n_44),
.B2(n_47),
.Y(n_94)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVxp33_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_66),
.C(n_69),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_50),
.B(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_57),
.B(n_60),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_52),
.A2(n_53),
.B1(n_86),
.B2(n_87),
.Y(n_90)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_53),
.B(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_63),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_63),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_61),
.B(n_79),
.Y(n_133)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g131 ( 
.A1(n_64),
.A2(n_132),
.B(n_133),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_66),
.A2(n_67),
.B1(n_69),
.B2(n_107),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_92),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_82),
.B2(n_83),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B(n_88),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_85),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_85),
.A2(n_88),
.B(n_129),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_85),
.B(n_97),
.Y(n_168)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_91),
.Y(n_88)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_89),
.A2(n_111),
.B1(n_113),
.B2(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_96),
.B(n_99),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_97),
.B(n_174),
.Y(n_173)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_108),
.C(n_114),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_104),
.A2(n_105),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_114),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_110),
.B(n_112),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_109),
.A2(n_112),
.B(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_117),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_115),
.B(n_117),
.Y(n_126)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_137),
.B(n_185),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_134),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_125),
.B(n_134),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.C(n_130),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_126),
.B(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_127),
.A2(n_130),
.B1(n_131),
.B2(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_127),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_179),
.B(n_184),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_156),
.B(n_178),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_150),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_150),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_146),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_142),
.B(n_145),
.C(n_146),
.Y(n_183)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_152),
.B1(n_154),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_154),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_166),
.B(n_177),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_164),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_164),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_160),
.A2(n_162),
.B(n_170),
.Y(n_169)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_171),
.B(n_176),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_169),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_175),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_183),
.Y(n_184)
);


endmodule