module fake_jpeg_7697_n_304 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_304);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_304;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_303;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_19),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_35),
.A2(n_27),
.B1(n_29),
.B2(n_33),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_44),
.Y(n_46)
);

CKINVDCx9p33_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_51),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_64),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_28),
.Y(n_48)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_28),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_20),
.B1(n_25),
.B2(n_17),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_55),
.B1(n_59),
.B2(n_18),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_20),
.B1(n_25),
.B2(n_26),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_38),
.B(n_32),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_70),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_62),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_25),
.B1(n_18),
.B2(n_31),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_29),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_31),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_69),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_35),
.B(n_22),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_27),
.B1(n_65),
.B2(n_54),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_71),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_33),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_42),
.B(n_22),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_68),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_76),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_68),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_68),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_82),
.Y(n_115)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_61),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_83),
.A2(n_63),
.B1(n_70),
.B2(n_58),
.Y(n_112)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_10),
.Y(n_102)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_91),
.Y(n_96)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

NAND2x1p5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_0),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_93),
.A2(n_48),
.B(n_21),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_71),
.B1(n_46),
.B2(n_45),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_99),
.A2(n_111),
.B1(n_112),
.B2(n_116),
.Y(n_133)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_106),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_102),
.A2(n_23),
.B(n_34),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_46),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_108),
.Y(n_123)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_107),
.B(n_110),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_80),
.B(n_64),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_61),
.B1(n_52),
.B2(n_56),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_69),
.C(n_57),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_94),
.C(n_72),
.Y(n_125)
);

BUFx24_ASAP7_75t_SL g114 ( 
.A(n_94),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_117),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_61),
.B1(n_56),
.B2(n_52),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_91),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_51),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_118),
.B(n_43),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_21),
.B(n_24),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_74),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_125),
.C(n_138),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_121),
.B(n_124),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_115),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_74),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_127),
.A2(n_129),
.B(n_137),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_0),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_92),
.Y(n_130)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_92),
.Y(n_131)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_136),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_82),
.B1(n_91),
.B2(n_90),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_135),
.A2(n_97),
.B1(n_103),
.B2(n_87),
.Y(n_151)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_76),
.C(n_73),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_77),
.Y(n_139)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_99),
.A2(n_81),
.B(n_43),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_140),
.A2(n_97),
.B(n_98),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_43),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_143),
.C(n_144),
.Y(n_160)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_143),
.Y(n_153)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_108),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_145),
.A2(n_119),
.B(n_24),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_147),
.A2(n_140),
.B(n_127),
.Y(n_181)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_162),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_151),
.A2(n_124),
.B1(n_134),
.B2(n_44),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_132),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_106),
.Y(n_154)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_132),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_155),
.B(n_159),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_142),
.A2(n_103),
.B1(n_117),
.B2(n_96),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_158),
.A2(n_170),
.B1(n_172),
.B2(n_87),
.Y(n_192)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_163),
.C(n_165),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_161),
.A2(n_167),
.B(n_145),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_136),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_102),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_138),
.C(n_125),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_98),
.C(n_96),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_137),
.C(n_128),
.Y(n_196)
);

AND2x4_ASAP7_75t_L g167 ( 
.A(n_121),
.B(n_102),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_133),
.A2(n_103),
.B1(n_60),
.B2(n_100),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_122),
.B(n_109),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_129),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_133),
.A2(n_60),
.B1(n_79),
.B2(n_75),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_152),
.Y(n_203)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_168),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_175),
.B(n_176),
.Y(n_220)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_171),
.Y(n_178)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_179),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_135),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_196),
.C(n_42),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_181),
.A2(n_190),
.B(n_197),
.Y(n_215)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_182),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_185),
.B1(n_188),
.B2(n_195),
.Y(n_217)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_184),
.Y(n_218)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_186),
.A2(n_194),
.B(n_44),
.Y(n_212)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_154),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_189),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_147),
.A2(n_127),
.B(n_129),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_149),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_191),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_192),
.A2(n_167),
.B1(n_156),
.B2(n_170),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_151),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_33),
.Y(n_197)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_192),
.A2(n_167),
.B1(n_172),
.B2(n_150),
.Y(n_200)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_173),
.A2(n_167),
.B1(n_146),
.B2(n_165),
.Y(n_201)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_201),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_173),
.A2(n_146),
.B1(n_164),
.B2(n_161),
.Y(n_202)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_202),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_205),
.C(n_208),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_163),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_181),
.A2(n_148),
.B1(n_169),
.B2(n_75),
.Y(n_206)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_206),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_169),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_1),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_189),
.B(n_197),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_190),
.A2(n_44),
.B1(n_81),
.B2(n_84),
.Y(n_211)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_9),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_219),
.C(n_196),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_191),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_183),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_1),
.C(n_2),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_221),
.A2(n_225),
.B(n_233),
.Y(n_246)
);

BUFx24_ASAP7_75t_SL g222 ( 
.A(n_220),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_227),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_210),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_231),
.Y(n_243)
);

OA21x2_ASAP7_75t_SL g225 ( 
.A1(n_202),
.A2(n_186),
.B(n_208),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_239),
.C(n_215),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_217),
.B(n_177),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_187),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_240),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_215),
.A2(n_195),
.B(n_3),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_219),
.B(n_9),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_236),
.B(n_14),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_237),
.A2(n_207),
.B1(n_199),
.B2(n_200),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_1),
.C(n_3),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_9),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_244),
.C(n_254),
.Y(n_257)
);

OA21x2_ASAP7_75t_L g242 ( 
.A1(n_235),
.A2(n_204),
.B(n_206),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_242),
.A2(n_238),
.B(n_226),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_205),
.C(n_201),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_232),
.B(n_218),
.Y(n_245)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_216),
.Y(n_249)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_252),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_211),
.Y(n_252)
);

INVxp33_ASAP7_75t_SL g253 ( 
.A(n_233),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_253),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_203),
.C(n_209),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_209),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_221),
.Y(n_261)
);

XNOR2x1_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_8),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_256),
.A2(n_239),
.B(n_4),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_260),
.B(n_265),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_6),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_246),
.A2(n_230),
.B(n_238),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_262),
.A2(n_256),
.B(n_242),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_242),
.A2(n_234),
.B1(n_229),
.B2(n_227),
.Y(n_263)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_263),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_251),
.B(n_234),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_247),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_253),
.A2(n_229),
.B1(n_3),
.B2(n_5),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_6),
.C(n_8),
.Y(n_279)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_264),
.A2(n_241),
.B1(n_243),
.B2(n_255),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_271),
.B(n_278),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_273),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_254),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_262),
.A2(n_4),
.B(n_5),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_277),
.C(n_268),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_5),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_258),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_269),
.A2(n_6),
.B(n_7),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_8),
.Y(n_285)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_259),
.Y(n_283)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_283),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_288),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_260),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_274),
.B(n_263),
.Y(n_288)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_289),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_257),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_280),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_281),
.A2(n_257),
.B(n_280),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_284),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_295),
.A2(n_298),
.B(n_292),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_296),
.Y(n_300)
);

AOI31xp67_ASAP7_75t_L g298 ( 
.A1(n_293),
.A2(n_287),
.A3(n_12),
.B(n_13),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_299),
.B(n_300),
.Y(n_301)
);

AOI321xp33_ASAP7_75t_L g302 ( 
.A1(n_301),
.A2(n_290),
.A3(n_13),
.B1(n_15),
.B2(n_16),
.C(n_11),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_15),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_15),
.Y(n_304)
);


endmodule