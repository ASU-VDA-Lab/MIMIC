module fake_jpeg_20874_n_301 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_282;
wire n_258;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_8),
.B(n_5),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_40),
.Y(n_49)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_20),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_44),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_32),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_20),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_42),
.A2(n_18),
.B1(n_15),
.B2(n_21),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_56),
.B1(n_60),
.B2(n_39),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_44),
.A2(n_18),
.B1(n_17),
.B2(n_15),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_44),
.B1(n_33),
.B2(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_59),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_27),
.Y(n_54)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_18),
.B1(n_15),
.B2(n_17),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_18),
.B1(n_15),
.B2(n_21),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_34),
.B1(n_40),
.B2(n_38),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_32),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_17),
.B1(n_26),
.B2(n_21),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_62),
.B(n_66),
.Y(n_109)
);

FAx1_ASAP7_75t_SL g65 ( 
.A(n_52),
.B(n_28),
.CI(n_39),
.CON(n_65),
.SN(n_65)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_65),
.B(n_84),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_19),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_67),
.A2(n_69),
.B1(n_30),
.B2(n_24),
.Y(n_126)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_45),
.A2(n_56),
.B1(n_51),
.B2(n_47),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_70),
.B(n_74),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_71),
.A2(n_85),
.B1(n_92),
.B2(n_99),
.Y(n_115)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_35),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_29),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_49),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_75),
.A2(n_30),
.B(n_24),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_60),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_76),
.B(n_82),
.Y(n_129)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_55),
.A2(n_26),
.B1(n_25),
.B2(n_23),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_81),
.A2(n_91),
.B1(n_95),
.B2(n_97),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_53),
.Y(n_82)
);

CKINVDCx5p33_ASAP7_75t_R g83 ( 
.A(n_55),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_93),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_54),
.B(n_23),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_58),
.A2(n_38),
.B1(n_34),
.B2(n_33),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_93),
.Y(n_134)
);

MAJx2_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_35),
.C(n_31),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_35),
.C(n_53),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_54),
.A2(n_31),
.B(n_19),
.C(n_28),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_48),
.B(n_29),
.C(n_43),
.Y(n_111)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_55),
.A2(n_25),
.B1(n_23),
.B2(n_19),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_59),
.A2(n_25),
.B1(n_19),
.B2(n_31),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_94),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_96),
.B(n_100),
.Y(n_105)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_35),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_101),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_47),
.A2(n_19),
.B1(n_31),
.B2(n_16),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_56),
.B(n_35),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_53),
.A2(n_31),
.B1(n_22),
.B2(n_16),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_85),
.B1(n_101),
.B2(n_79),
.Y(n_119)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_103),
.A2(n_24),
.B1(n_22),
.B2(n_16),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_98),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_48),
.B1(n_57),
.B2(n_43),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_110),
.A2(n_80),
.B1(n_90),
.B2(n_83),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_113),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_63),
.A2(n_57),
.B1(n_48),
.B2(n_29),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_112),
.A2(n_127),
.B(n_63),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_114),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_119),
.A2(n_130),
.B1(n_69),
.B2(n_68),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_73),
.B(n_30),
.C(n_24),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_75),
.C(n_67),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_131),
.Y(n_147)
);

AND2x4_ASAP7_75t_SL g127 ( 
.A(n_65),
.B(n_30),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_78),
.B1(n_97),
.B2(n_103),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_100),
.A2(n_22),
.B1(n_1),
.B2(n_2),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_88),
.A2(n_22),
.B(n_1),
.C(n_2),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_86),
.B1(n_129),
.B2(n_105),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_137),
.A2(n_139),
.B1(n_144),
.B2(n_154),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_142),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_72),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_148),
.Y(n_173)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_151),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_65),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_135),
.B(n_64),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_150),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_105),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_134),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_64),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_157),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_153),
.A2(n_111),
.B1(n_131),
.B2(n_121),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_119),
.A2(n_75),
.B1(n_87),
.B2(n_77),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_108),
.B(n_89),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_155),
.B(n_164),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_104),
.B(n_106),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_133),
.Y(n_158)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_106),
.B(n_75),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_159),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_120),
.A2(n_95),
.B1(n_94),
.B2(n_61),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_110),
.B1(n_130),
.B2(n_133),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_120),
.A2(n_0),
.B(n_1),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_116),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_129),
.B(n_2),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_165),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_113),
.B(n_2),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_3),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_123),
.B1(n_115),
.B2(n_127),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_166),
.A2(n_192),
.B1(n_183),
.B2(n_169),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_143),
.A2(n_123),
.B1(n_115),
.B2(n_126),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_170),
.A2(n_183),
.B1(n_188),
.B2(n_193),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_158),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_187),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_155),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_109),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_178),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_179),
.A2(n_182),
.B1(n_190),
.B2(n_162),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_139),
.A2(n_114),
.B1(n_107),
.B2(n_109),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_147),
.A2(n_118),
.B1(n_112),
.B2(n_116),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_137),
.B(n_132),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_185),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_160),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_145),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_159),
.A2(n_136),
.B1(n_111),
.B2(n_131),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_189),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_154),
.A2(n_136),
.B1(n_132),
.B2(n_125),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_147),
.A2(n_125),
.B1(n_117),
.B2(n_122),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_144),
.Y(n_194)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_193),
.B(n_148),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_195),
.A2(n_200),
.B(n_205),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_196),
.B(n_175),
.Y(n_226)
);

BUFx24_ASAP7_75t_SL g198 ( 
.A(n_178),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_215),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_191),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_201),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_150),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_189),
.A2(n_151),
.B1(n_122),
.B2(n_146),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_204),
.A2(n_208),
.B1(n_216),
.B2(n_219),
.Y(n_222)
);

NAND3xp33_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_141),
.C(n_165),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_138),
.Y(n_207)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_194),
.A2(n_141),
.B1(n_149),
.B2(n_153),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_209),
.A2(n_210),
.B1(n_195),
.B2(n_211),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_172),
.A2(n_152),
.B1(n_163),
.B2(n_142),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_168),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_212),
.B(n_214),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_164),
.Y(n_213)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_117),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_3),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_170),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_176),
.C(n_177),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_225),
.C(n_232),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_176),
.C(n_177),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_230),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_212),
.B(n_173),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_228),
.B(n_215),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_182),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_186),
.B(n_167),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_231),
.A2(n_235),
.B(n_202),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_172),
.C(n_184),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_167),
.C(n_166),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_202),
.C(n_209),
.Y(n_244)
);

O2A1O1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_211),
.A2(n_174),
.B(n_169),
.C(n_180),
.Y(n_234)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

AND2x4_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_186),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_236),
.A2(n_179),
.B1(n_197),
.B2(n_216),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_200),
.B(n_171),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_239),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_180),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_223),
.B(n_203),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_249),
.Y(n_258)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_253),
.C(n_238),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_222),
.A2(n_218),
.B1(n_195),
.B2(n_217),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_247),
.Y(n_262)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_219),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_227),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_250),
.B(n_220),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_251),
.A2(n_236),
.B(n_233),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_252),
.A2(n_255),
.B1(n_234),
.B2(n_235),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_199),
.C(n_197),
.Y(n_253)
);

INVxp33_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_254),
.A2(n_229),
.B1(n_237),
.B2(n_8),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_239),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_4),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_257),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_5),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_259),
.B(n_260),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_224),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_261),
.A2(n_245),
.B1(n_255),
.B2(n_253),
.Y(n_272)
);

NOR2x1_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_235),
.Y(n_265)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_265),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_266),
.A2(n_13),
.B(n_9),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_267),
.A2(n_257),
.B1(n_8),
.B2(n_9),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_269),
.C(n_241),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_243),
.B(n_13),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_244),
.B(n_6),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_270),
.B(n_7),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_272),
.A2(n_274),
.B1(n_264),
.B2(n_269),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_273),
.B(n_276),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_265),
.A2(n_249),
.B(n_248),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_275),
.A2(n_260),
.B(n_266),
.Y(n_280)
);

AOI322xp5_ASAP7_75t_L g276 ( 
.A1(n_262),
.A2(n_256),
.A3(n_248),
.B1(n_243),
.B2(n_241),
.C1(n_7),
.C2(n_11),
.Y(n_276)
);

MAJx2_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_10),
.C(n_11),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_278),
.B(n_10),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_282),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_268),
.C(n_258),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_279),
.A2(n_261),
.B(n_263),
.Y(n_283)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_283),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_284),
.A2(n_286),
.B1(n_287),
.B2(n_279),
.Y(n_289)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_285),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_277),
.A2(n_258),
.B1(n_264),
.B2(n_13),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_289),
.B(n_291),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_281),
.A2(n_271),
.B(n_275),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_282),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_294),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_283),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_295),
.B(n_292),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_297),
.A2(n_296),
.B(n_290),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_293),
.C(n_286),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_10),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_11),
.Y(n_301)
);


endmodule