module real_aes_6978_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_0), .B(n_108), .C(n_109), .Y(n_107) );
INVx1_ASAP7_75t_L g463 ( .A(n_0), .Y(n_463) );
INVx1_ASAP7_75t_L g497 ( .A(n_1), .Y(n_497) );
INVx1_ASAP7_75t_L g204 ( .A(n_2), .Y(n_204) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_3), .A2(n_37), .B1(n_165), .B2(n_527), .Y(n_542) );
AOI21xp33_ASAP7_75t_L g172 ( .A1(n_4), .A2(n_146), .B(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_5), .B(n_139), .Y(n_510) );
AND2x6_ASAP7_75t_L g151 ( .A(n_6), .B(n_152), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_7), .A2(n_254), .B(n_255), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_8), .B(n_38), .Y(n_113) );
INVx1_ASAP7_75t_L g179 ( .A(n_9), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_10), .B(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g144 ( .A(n_11), .Y(n_144) );
INVx1_ASAP7_75t_L g491 ( .A(n_12), .Y(n_491) );
INVx1_ASAP7_75t_L g260 ( .A(n_13), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_14), .B(n_187), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_15), .B(n_140), .Y(n_568) );
AO32x2_ASAP7_75t_L g540 ( .A1(n_16), .A2(n_139), .A3(n_184), .B1(n_519), .B2(n_541), .Y(n_540) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_17), .A2(n_63), .B1(n_128), .B2(n_129), .Y(n_127) );
INVx1_ASAP7_75t_L g129 ( .A(n_17), .Y(n_129) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_18), .B(n_165), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_19), .B(n_160), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_20), .B(n_140), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_21), .A2(n_51), .B1(n_165), .B2(n_527), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_22), .B(n_146), .Y(n_216) );
AOI22xp33_ASAP7_75t_SL g528 ( .A1(n_23), .A2(n_80), .B1(n_165), .B2(n_187), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_24), .B(n_165), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_25), .B(n_168), .Y(n_167) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_26), .A2(n_258), .B(n_259), .C(n_261), .Y(n_257) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_27), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_28), .B(n_181), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_29), .B(n_177), .Y(n_206) );
INVx1_ASAP7_75t_L g193 ( .A(n_30), .Y(n_193) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_31), .A2(n_32), .B1(n_122), .B2(n_123), .Y(n_121) );
INVx1_ASAP7_75t_L g123 ( .A(n_31), .Y(n_123) );
INVxp67_ASAP7_75t_L g122 ( .A(n_32), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_32), .B(n_181), .Y(n_557) );
INVx2_ASAP7_75t_L g149 ( .A(n_33), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_34), .B(n_165), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_35), .B(n_181), .Y(n_539) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_36), .A2(n_151), .B(n_155), .C(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g191 ( .A(n_39), .Y(n_191) );
OAI22xp5_ASAP7_75t_SL g470 ( .A1(n_40), .A2(n_471), .B1(n_474), .B2(n_475), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_40), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_41), .B(n_177), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_42), .B(n_165), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_43), .A2(n_90), .B1(n_223), .B2(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_44), .B(n_165), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_45), .B(n_165), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_46), .A2(n_105), .B1(n_114), .B2(n_776), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g194 ( .A(n_47), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_48), .A2(n_70), .B1(n_472), .B2(n_473), .Y(n_471) );
CKINVDCx16_ASAP7_75t_R g473 ( .A(n_48), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_49), .B(n_496), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_50), .B(n_146), .Y(n_248) );
AOI22xp33_ASAP7_75t_SL g566 ( .A1(n_52), .A2(n_61), .B1(n_165), .B2(n_187), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_53), .A2(n_155), .B1(n_187), .B2(n_189), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_54), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_55), .B(n_165), .Y(n_518) );
CKINVDCx16_ASAP7_75t_R g201 ( .A(n_56), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_57), .B(n_165), .Y(n_533) );
A2O1A1Ixp33_ASAP7_75t_L g175 ( .A1(n_58), .A2(n_164), .B(n_176), .C(n_178), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_59), .Y(n_236) );
INVx1_ASAP7_75t_L g174 ( .A(n_60), .Y(n_174) );
INVx1_ASAP7_75t_L g152 ( .A(n_62), .Y(n_152) );
INVx1_ASAP7_75t_L g128 ( .A(n_63), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_64), .B(n_165), .Y(n_498) );
INVx1_ASAP7_75t_L g143 ( .A(n_65), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_66), .Y(n_118) );
AO32x2_ASAP7_75t_L g524 ( .A1(n_67), .A2(n_139), .A3(n_240), .B1(n_519), .B2(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g517 ( .A(n_68), .Y(n_517) );
INVx1_ASAP7_75t_L g552 ( .A(n_69), .Y(n_552) );
INVx1_ASAP7_75t_L g472 ( .A(n_70), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_SL g159 ( .A1(n_71), .A2(n_160), .B(n_161), .C(n_164), .Y(n_159) );
INVxp67_ASAP7_75t_L g162 ( .A(n_72), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_73), .B(n_187), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_74), .A2(n_469), .B1(n_470), .B2(n_476), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_74), .Y(n_469) );
INVx1_ASAP7_75t_L g111 ( .A(n_75), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_76), .B(n_459), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_77), .A2(n_461), .B1(n_467), .B2(n_771), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g197 ( .A(n_78), .Y(n_197) );
INVx1_ASAP7_75t_L g229 ( .A(n_79), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_81), .A2(n_151), .B(n_155), .C(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_82), .B(n_527), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_83), .B(n_187), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_84), .B(n_205), .Y(n_219) );
INVx2_ASAP7_75t_L g141 ( .A(n_85), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_86), .B(n_160), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_87), .B(n_187), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_88), .A2(n_151), .B(n_155), .C(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g108 ( .A(n_89), .Y(n_108) );
OR2x2_ASAP7_75t_L g460 ( .A(n_89), .B(n_461), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_91), .A2(n_103), .B1(n_187), .B2(n_188), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_92), .B(n_181), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g209 ( .A(n_93), .Y(n_209) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_94), .A2(n_151), .B(n_155), .C(n_243), .Y(n_242) );
CKINVDCx20_ASAP7_75t_R g250 ( .A(n_95), .Y(n_250) );
INVx1_ASAP7_75t_L g158 ( .A(n_96), .Y(n_158) );
CKINVDCx16_ASAP7_75t_R g256 ( .A(n_97), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_98), .B(n_205), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_99), .B(n_187), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_100), .B(n_139), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_101), .B(n_111), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_102), .A2(n_146), .B(n_153), .Y(n_145) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_106), .Y(n_778) );
OR2x2_ASAP7_75t_SL g106 ( .A(n_107), .B(n_112), .Y(n_106) );
AOI22xp5_ASAP7_75t_SL g477 ( .A1(n_108), .A2(n_130), .B1(n_478), .B2(n_770), .Y(n_477) );
INVx2_ASAP7_75t_L g770 ( .A(n_108), .Y(n_770) );
NOR2x2_ASAP7_75t_L g773 ( .A(n_108), .B(n_461), .Y(n_773) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVxp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_L g462 ( .A(n_113), .B(n_463), .Y(n_462) );
AO21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_119), .B(n_465), .Y(n_114) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g775 ( .A(n_118), .Y(n_775) );
OAI21xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_457), .B(n_464), .Y(n_119) );
AOI22xp33_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_124), .B1(n_125), .B2(n_456), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_121), .Y(n_456) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI22xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_127), .B1(n_130), .B2(n_455), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g455 ( .A(n_130), .Y(n_455) );
INVx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND4x1_ASAP7_75t_L g131 ( .A(n_132), .B(n_373), .C(n_420), .D(n_440), .Y(n_131) );
NOR3xp33_ASAP7_75t_SL g132 ( .A(n_133), .B(n_303), .C(n_328), .Y(n_132) );
OAI211xp5_ASAP7_75t_SL g133 ( .A1(n_134), .A2(n_211), .B(n_263), .C(n_293), .Y(n_133) );
INVxp67_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_136), .B(n_182), .Y(n_135) );
INVx3_ASAP7_75t_SL g345 ( .A(n_136), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_136), .B(n_276), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_136), .B(n_198), .Y(n_426) );
AND2x2_ASAP7_75t_L g449 ( .A(n_136), .B(n_315), .Y(n_449) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_170), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g267 ( .A(n_138), .B(n_171), .Y(n_267) );
INVx3_ASAP7_75t_L g280 ( .A(n_138), .Y(n_280) );
AND2x2_ASAP7_75t_L g285 ( .A(n_138), .B(n_170), .Y(n_285) );
OR2x2_ASAP7_75t_L g336 ( .A(n_138), .B(n_277), .Y(n_336) );
BUFx2_ASAP7_75t_L g356 ( .A(n_138), .Y(n_356) );
AND2x2_ASAP7_75t_L g366 ( .A(n_138), .B(n_277), .Y(n_366) );
AND2x2_ASAP7_75t_L g372 ( .A(n_138), .B(n_183), .Y(n_372) );
OA21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_145), .B(n_167), .Y(n_138) );
INVx4_ASAP7_75t_L g169 ( .A(n_139), .Y(n_169) );
OA21x2_ASAP7_75t_L g502 ( .A1(n_139), .A2(n_503), .B(n_510), .Y(n_502) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g184 ( .A(n_140), .Y(n_184) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x2_ASAP7_75t_SL g181 ( .A(n_141), .B(n_142), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
BUFx2_ASAP7_75t_L g254 ( .A(n_146), .Y(n_254) );
AND2x4_ASAP7_75t_L g146 ( .A(n_147), .B(n_151), .Y(n_146) );
NAND2x1p5_ASAP7_75t_L g195 ( .A(n_147), .B(n_151), .Y(n_195) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_150), .Y(n_147) );
INVx1_ASAP7_75t_L g496 ( .A(n_148), .Y(n_496) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g156 ( .A(n_149), .Y(n_156) );
INVx1_ASAP7_75t_L g188 ( .A(n_149), .Y(n_188) );
INVx1_ASAP7_75t_L g157 ( .A(n_150), .Y(n_157) );
INVx1_ASAP7_75t_L g160 ( .A(n_150), .Y(n_160) );
INVx3_ASAP7_75t_L g163 ( .A(n_150), .Y(n_163) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_150), .Y(n_177) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_150), .Y(n_190) );
INVx4_ASAP7_75t_SL g166 ( .A(n_151), .Y(n_166) );
OAI21xp5_ASAP7_75t_L g489 ( .A1(n_151), .A2(n_490), .B(n_494), .Y(n_489) );
OAI21xp5_ASAP7_75t_L g503 ( .A1(n_151), .A2(n_504), .B(n_507), .Y(n_503) );
BUFx3_ASAP7_75t_L g519 ( .A(n_151), .Y(n_519) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_151), .A2(n_532), .B(n_536), .Y(n_531) );
OAI21xp5_ASAP7_75t_L g550 ( .A1(n_151), .A2(n_551), .B(n_554), .Y(n_550) );
O2A1O1Ixp33_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_158), .B(n_159), .C(n_166), .Y(n_153) );
O2A1O1Ixp33_ASAP7_75t_L g173 ( .A1(n_154), .A2(n_166), .B(n_174), .C(n_175), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_L g255 ( .A1(n_154), .A2(n_166), .B(n_256), .C(n_257), .Y(n_255) );
INVx5_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AND2x6_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_156), .Y(n_165) );
BUFx3_ASAP7_75t_L g223 ( .A(n_156), .Y(n_223) );
INVx1_ASAP7_75t_L g527 ( .A(n_156), .Y(n_527) );
INVx1_ASAP7_75t_L g535 ( .A(n_160), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_162), .B(n_163), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_163), .B(n_179), .Y(n_178) );
INVx5_ASAP7_75t_L g205 ( .A(n_163), .Y(n_205) );
OAI22xp5_ASAP7_75t_SL g525 ( .A1(n_163), .A2(n_177), .B1(n_526), .B2(n_528), .Y(n_525) );
O2A1O1Ixp5_ASAP7_75t_SL g551 ( .A1(n_164), .A2(n_205), .B(n_552), .C(n_553), .Y(n_551) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_165), .Y(n_247) );
OAI22xp33_ASAP7_75t_L g185 ( .A1(n_166), .A2(n_186), .B1(n_194), .B2(n_195), .Y(n_185) );
OA21x2_ASAP7_75t_L g171 ( .A1(n_168), .A2(n_172), .B(n_180), .Y(n_171) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_SL g225 ( .A(n_169), .B(n_226), .Y(n_225) );
AO21x1_ASAP7_75t_L g563 ( .A1(n_169), .A2(n_564), .B(n_567), .Y(n_563) );
NAND3xp33_ASAP7_75t_L g582 ( .A(n_169), .B(n_519), .C(n_564), .Y(n_582) );
INVx1_ASAP7_75t_SL g170 ( .A(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_171), .B(n_277), .Y(n_291) );
INVx2_ASAP7_75t_L g301 ( .A(n_171), .Y(n_301) );
AND2x2_ASAP7_75t_L g314 ( .A(n_171), .B(n_280), .Y(n_314) );
OR2x2_ASAP7_75t_L g325 ( .A(n_171), .B(n_277), .Y(n_325) );
AND2x2_ASAP7_75t_SL g371 ( .A(n_171), .B(n_372), .Y(n_371) );
BUFx2_ASAP7_75t_L g383 ( .A(n_171), .Y(n_383) );
AND2x2_ASAP7_75t_L g429 ( .A(n_171), .B(n_183), .Y(n_429) );
O2A1O1Ixp5_ASAP7_75t_L g516 ( .A1(n_176), .A2(n_495), .B(n_517), .C(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_176), .A2(n_537), .B(n_538), .Y(n_536) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx4_ASAP7_75t_L g246 ( .A(n_177), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_177), .A2(n_499), .B1(n_542), .B2(n_543), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_177), .A2(n_499), .B1(n_565), .B2(n_566), .Y(n_564) );
INVx1_ASAP7_75t_L g210 ( .A(n_181), .Y(n_210) );
INVx2_ASAP7_75t_L g240 ( .A(n_181), .Y(n_240) );
OA21x2_ASAP7_75t_L g252 ( .A1(n_181), .A2(n_253), .B(n_262), .Y(n_252) );
OA21x2_ASAP7_75t_L g530 ( .A1(n_181), .A2(n_531), .B(n_539), .Y(n_530) );
OA21x2_ASAP7_75t_L g549 ( .A1(n_181), .A2(n_550), .B(n_557), .Y(n_549) );
INVx3_ASAP7_75t_SL g302 ( .A(n_182), .Y(n_302) );
OR2x2_ASAP7_75t_L g355 ( .A(n_182), .B(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_198), .Y(n_182) );
INVx3_ASAP7_75t_L g277 ( .A(n_183), .Y(n_277) );
AND2x2_ASAP7_75t_L g344 ( .A(n_183), .B(n_199), .Y(n_344) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_183), .Y(n_412) );
AOI33xp33_ASAP7_75t_L g416 ( .A1(n_183), .A2(n_345), .A3(n_352), .B1(n_361), .B2(n_417), .B3(n_418), .Y(n_416) );
AO21x2_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_196), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_184), .B(n_197), .Y(n_196) );
AO21x2_ASAP7_75t_L g199 ( .A1(n_184), .A2(n_200), .B(n_208), .Y(n_199) );
INVx2_ASAP7_75t_L g224 ( .A(n_184), .Y(n_224) );
INVx2_ASAP7_75t_L g207 ( .A(n_187), .Y(n_207) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
OAI22xp5_ASAP7_75t_SL g189 ( .A1(n_190), .A2(n_191), .B1(n_192), .B2(n_193), .Y(n_189) );
INVx2_ASAP7_75t_L g192 ( .A(n_190), .Y(n_192) );
INVx4_ASAP7_75t_L g258 ( .A(n_190), .Y(n_258) );
OAI21xp5_ASAP7_75t_L g200 ( .A1(n_195), .A2(n_201), .B(n_202), .Y(n_200) );
OAI21xp5_ASAP7_75t_L g228 ( .A1(n_195), .A2(n_229), .B(n_230), .Y(n_228) );
INVx1_ASAP7_75t_L g265 ( .A(n_198), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_198), .B(n_280), .Y(n_279) );
NOR3xp33_ASAP7_75t_L g339 ( .A(n_198), .B(n_340), .C(n_342), .Y(n_339) );
AND2x2_ASAP7_75t_L g365 ( .A(n_198), .B(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_198), .B(n_372), .Y(n_375) );
AND2x2_ASAP7_75t_L g428 ( .A(n_198), .B(n_429), .Y(n_428) );
INVx3_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx3_ASAP7_75t_L g284 ( .A(n_199), .Y(n_284) );
OR2x2_ASAP7_75t_L g378 ( .A(n_199), .B(n_277), .Y(n_378) );
O2A1O1Ixp33_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_206), .C(n_207), .Y(n_203) );
INVx2_ASAP7_75t_L g499 ( .A(n_205), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_205), .A2(n_505), .B(n_506), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_205), .A2(n_514), .B(n_515), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_207), .A2(n_491), .B(n_492), .C(n_493), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_210), .B(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_210), .B(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_237), .Y(n_211) );
AOI32xp33_ASAP7_75t_L g329 ( .A1(n_212), .A2(n_330), .A3(n_332), .B1(n_334), .B2(n_337), .Y(n_329) );
NOR2xp67_ASAP7_75t_L g402 ( .A(n_212), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g432 ( .A(n_212), .Y(n_432) );
INVx4_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g364 ( .A(n_213), .B(n_348), .Y(n_364) );
AND2x2_ASAP7_75t_L g384 ( .A(n_213), .B(n_310), .Y(n_384) );
AND2x2_ASAP7_75t_L g452 ( .A(n_213), .B(n_370), .Y(n_452) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_227), .Y(n_213) );
INVx3_ASAP7_75t_L g273 ( .A(n_214), .Y(n_273) );
AND2x2_ASAP7_75t_L g287 ( .A(n_214), .B(n_271), .Y(n_287) );
OR2x2_ASAP7_75t_L g292 ( .A(n_214), .B(n_270), .Y(n_292) );
INVx1_ASAP7_75t_L g299 ( .A(n_214), .Y(n_299) );
AND2x2_ASAP7_75t_L g307 ( .A(n_214), .B(n_281), .Y(n_307) );
AND2x2_ASAP7_75t_L g309 ( .A(n_214), .B(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_214), .B(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g362 ( .A(n_214), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_214), .B(n_447), .Y(n_446) );
OR2x6_ASAP7_75t_L g214 ( .A(n_215), .B(n_225), .Y(n_214) );
AOI21xp5_ASAP7_75t_SL g215 ( .A1(n_216), .A2(n_217), .B(n_224), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_221), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_221), .A2(n_232), .B(n_233), .Y(n_231) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g261 ( .A(n_223), .Y(n_261) );
INVx1_ASAP7_75t_L g234 ( .A(n_224), .Y(n_234) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_224), .A2(n_489), .B(n_500), .Y(n_488) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_224), .A2(n_512), .B(n_520), .Y(n_511) );
INVx2_ASAP7_75t_L g271 ( .A(n_227), .Y(n_271) );
AND2x2_ASAP7_75t_L g317 ( .A(n_227), .B(n_238), .Y(n_317) );
AND2x2_ASAP7_75t_L g327 ( .A(n_227), .B(n_252), .Y(n_327) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_234), .B(n_235), .Y(n_227) );
INVx2_ASAP7_75t_L g447 ( .A(n_237), .Y(n_447) );
OR2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_251), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_238), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g288 ( .A(n_238), .Y(n_288) );
AND2x2_ASAP7_75t_L g332 ( .A(n_238), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g348 ( .A(n_238), .B(n_311), .Y(n_348) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g296 ( .A(n_239), .Y(n_296) );
AND2x2_ASAP7_75t_L g310 ( .A(n_239), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g361 ( .A(n_239), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_239), .B(n_271), .Y(n_393) );
AO21x2_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B(n_249), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_248), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_247), .Y(n_243) );
AND2x2_ASAP7_75t_L g272 ( .A(n_251), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g333 ( .A(n_251), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_251), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g370 ( .A(n_251), .Y(n_370) );
INVx1_ASAP7_75t_L g403 ( .A(n_251), .Y(n_403) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g281 ( .A(n_252), .B(n_271), .Y(n_281) );
INVx1_ASAP7_75t_L g311 ( .A(n_252), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_258), .B(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g493 ( .A(n_258), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_258), .A2(n_555), .B(n_556), .Y(n_554) );
AOI221xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_268), .B1(n_274), .B2(n_281), .C(n_282), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_265), .B(n_285), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_265), .B(n_348), .Y(n_425) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_267), .B(n_315), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_267), .B(n_276), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_267), .B(n_290), .Y(n_419) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_272), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g341 ( .A(n_271), .Y(n_341) );
AND2x2_ASAP7_75t_L g316 ( .A(n_272), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g394 ( .A(n_272), .Y(n_394) );
AND2x2_ASAP7_75t_L g326 ( .A(n_273), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_273), .B(n_296), .Y(n_342) );
AND2x2_ASAP7_75t_L g406 ( .A(n_273), .B(n_332), .Y(n_406) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
BUFx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g315 ( .A(n_277), .B(n_284), .Y(n_315) );
AND2x2_ASAP7_75t_L g411 ( .A(n_278), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_280), .B(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_281), .B(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_281), .B(n_288), .Y(n_376) );
AND2x2_ASAP7_75t_L g396 ( .A(n_281), .B(n_296), .Y(n_396) );
AND2x2_ASAP7_75t_L g417 ( .A(n_281), .B(n_361), .Y(n_417) );
OAI32xp33_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_286), .A3(n_288), .B1(n_289), .B2(n_292), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx1_ASAP7_75t_SL g290 ( .A(n_284), .Y(n_290) );
NAND2x1_ASAP7_75t_L g331 ( .A(n_284), .B(n_314), .Y(n_331) );
OR2x2_ASAP7_75t_L g335 ( .A(n_284), .B(n_336), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_284), .B(n_383), .Y(n_436) );
INVx1_ASAP7_75t_L g304 ( .A(n_285), .Y(n_304) );
OAI221xp5_ASAP7_75t_SL g422 ( .A1(n_286), .A2(n_377), .B1(n_423), .B2(n_426), .C(n_427), .Y(n_422) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g294 ( .A(n_287), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g337 ( .A(n_287), .B(n_310), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_287), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g415 ( .A(n_287), .B(n_348), .Y(n_415) );
INVxp67_ASAP7_75t_L g351 ( .A(n_288), .Y(n_351) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
AND2x2_ASAP7_75t_L g421 ( .A(n_290), .B(n_408), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_290), .B(n_371), .Y(n_444) );
INVx1_ASAP7_75t_L g319 ( .A(n_292), .Y(n_319) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_292), .B(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g437 ( .A(n_292), .B(n_438), .Y(n_437) );
OAI21xp5_ASAP7_75t_SL g293 ( .A1(n_294), .A2(n_297), .B(n_300), .Y(n_293) );
AND2x2_ASAP7_75t_L g306 ( .A(n_295), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g390 ( .A(n_299), .B(n_310), .Y(n_390) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
AND2x2_ASAP7_75t_L g408 ( .A(n_301), .B(n_366), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_301), .B(n_365), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_302), .B(n_314), .Y(n_388) );
OAI211xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_305), .B(n_308), .C(n_318), .Y(n_303) );
AOI221xp5_ASAP7_75t_L g338 ( .A1(n_304), .A2(n_339), .B1(n_343), .B2(n_346), .C(n_349), .Y(n_338) );
AOI31xp33_ASAP7_75t_L g433 ( .A1(n_304), .A2(n_434), .A3(n_435), .B(n_437), .Y(n_433) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_312), .B1(n_314), .B2(n_316), .Y(n_308) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx1_ASAP7_75t_L g434 ( .A(n_314), .Y(n_434) );
INVx1_ASAP7_75t_L g397 ( .A(n_315), .Y(n_397) );
O2A1O1Ixp33_ASAP7_75t_L g440 ( .A1(n_317), .A2(n_441), .B(n_443), .C(n_445), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_320), .B1(n_322), .B2(n_326), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_323), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OAI221xp5_ASAP7_75t_SL g413 ( .A1(n_325), .A2(n_359), .B1(n_378), .B2(n_414), .C(n_416), .Y(n_413) );
INVx1_ASAP7_75t_L g409 ( .A(n_326), .Y(n_409) );
INVx1_ASAP7_75t_L g363 ( .A(n_327), .Y(n_363) );
NAND3xp33_ASAP7_75t_SL g328 ( .A(n_329), .B(n_338), .C(n_353), .Y(n_328) );
OAI21xp33_ASAP7_75t_L g379 ( .A1(n_330), .A2(n_380), .B(n_384), .Y(n_379) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_332), .B(n_432), .Y(n_431) );
INVxp67_ASAP7_75t_L g439 ( .A(n_333), .Y(n_439) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g377 ( .A(n_340), .B(n_360), .Y(n_377) );
INVx1_ASAP7_75t_L g352 ( .A(n_341), .Y(n_352) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_L g350 ( .A(n_344), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_344), .B(n_382), .Y(n_381) );
NOR4xp25_ASAP7_75t_L g349 ( .A(n_345), .B(n_350), .C(n_351), .D(n_352), .Y(n_349) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AOI222xp33_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_358), .B1(n_364), .B2(n_365), .C1(n_367), .C2(n_371), .Y(n_353) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_355), .B(n_357), .Y(n_354) );
INVx1_ASAP7_75t_L g451 ( .A(n_355), .Y(n_451) );
INVx1_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_363), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_367), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OAI21xp5_ASAP7_75t_SL g427 ( .A1(n_372), .A2(n_428), .B(n_430), .Y(n_427) );
NOR4xp25_ASAP7_75t_L g373 ( .A(n_374), .B(n_385), .C(n_398), .D(n_413), .Y(n_373) );
OAI221xp5_ASAP7_75t_SL g374 ( .A1(n_375), .A2(n_376), .B1(n_377), .B2(n_378), .C(n_379), .Y(n_374) );
INVx1_ASAP7_75t_L g454 ( .A(n_375), .Y(n_454) );
INVx1_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_382), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
OAI222xp33_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_389), .B1(n_391), .B2(n_392), .C1(n_395), .C2(n_397), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI211xp5_ASAP7_75t_L g420 ( .A1(n_390), .A2(n_421), .B(n_422), .C(n_433), .Y(n_420) );
OR2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx1_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
OAI222xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_404), .B1(n_405), .B2(n_407), .C1(n_409), .C2(n_410), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVxp67_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_415), .A2(n_418), .B1(n_451), .B2(n_452), .Y(n_450) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OAI211xp5_ASAP7_75t_SL g445 ( .A1(n_446), .A2(n_448), .B(n_450), .C(n_453), .Y(n_445) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_464), .A2(n_466), .B(n_774), .Y(n_465) );
XNOR2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_477), .Y(n_467) );
INVx1_ASAP7_75t_L g476 ( .A(n_470), .Y(n_476) );
INVx1_ASAP7_75t_L g474 ( .A(n_471), .Y(n_474) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_SL g479 ( .A(n_480), .B(n_736), .Y(n_479) );
NOR3xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_640), .C(n_724), .Y(n_480) );
NAND4xp25_ASAP7_75t_L g481 ( .A(n_482), .B(n_583), .C(n_605), .D(n_621), .Y(n_481) );
AOI221xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_521), .B1(n_544), .B2(n_562), .C(n_569), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_501), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_485), .B(n_562), .Y(n_595) );
NAND4xp25_ASAP7_75t_L g635 ( .A(n_485), .B(n_623), .C(n_636), .D(n_638), .Y(n_635) );
INVxp67_ASAP7_75t_L g752 ( .A(n_485), .Y(n_752) );
INVx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OR2x2_ASAP7_75t_L g634 ( .A(n_486), .B(n_572), .Y(n_634) );
AND2x2_ASAP7_75t_L g658 ( .A(n_486), .B(n_501), .Y(n_658) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g625 ( .A(n_487), .B(n_561), .Y(n_625) );
AND2x2_ASAP7_75t_L g665 ( .A(n_487), .B(n_646), .Y(n_665) );
AND2x2_ASAP7_75t_L g682 ( .A(n_487), .B(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_487), .B(n_502), .Y(n_706) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g560 ( .A(n_488), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g577 ( .A(n_488), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g589 ( .A(n_488), .B(n_502), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_488), .B(n_511), .Y(n_611) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_497), .B(n_498), .C(n_499), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_499), .A2(n_508), .B(n_509), .Y(n_507) );
AND2x2_ASAP7_75t_L g592 ( .A(n_501), .B(n_593), .Y(n_592) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_501), .A2(n_642), .B1(n_645), .B2(n_647), .C(n_651), .Y(n_641) );
AND2x2_ASAP7_75t_L g700 ( .A(n_501), .B(n_665), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_501), .B(n_682), .Y(n_734) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_511), .Y(n_501) );
INVx3_ASAP7_75t_L g561 ( .A(n_502), .Y(n_561) );
AND2x2_ASAP7_75t_L g609 ( .A(n_502), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g663 ( .A(n_502), .B(n_578), .Y(n_663) );
AND2x2_ASAP7_75t_L g721 ( .A(n_502), .B(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g562 ( .A(n_511), .B(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g578 ( .A(n_511), .Y(n_578) );
INVx1_ASAP7_75t_L g633 ( .A(n_511), .Y(n_633) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_511), .Y(n_639) );
AND2x2_ASAP7_75t_L g684 ( .A(n_511), .B(n_561), .Y(n_684) );
OR2x2_ASAP7_75t_L g723 ( .A(n_511), .B(n_563), .Y(n_723) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_516), .B(n_519), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_521), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_529), .Y(n_521) );
AND2x2_ASAP7_75t_L g719 ( .A(n_522), .B(n_716), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_522), .B(n_701), .Y(n_751) );
BUFx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g650 ( .A(n_523), .B(n_574), .Y(n_650) );
AND2x2_ASAP7_75t_L g699 ( .A(n_523), .B(n_547), .Y(n_699) );
INVx1_ASAP7_75t_L g745 ( .A(n_523), .Y(n_745) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_524), .Y(n_559) );
AND2x2_ASAP7_75t_L g600 ( .A(n_524), .B(n_574), .Y(n_600) );
INVx1_ASAP7_75t_L g617 ( .A(n_524), .Y(n_617) );
AND2x2_ASAP7_75t_L g623 ( .A(n_524), .B(n_540), .Y(n_623) );
AND2x2_ASAP7_75t_L g691 ( .A(n_529), .B(n_599), .Y(n_691) );
INVx2_ASAP7_75t_L g756 ( .A(n_529), .Y(n_756) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_540), .Y(n_529) );
AND2x2_ASAP7_75t_L g573 ( .A(n_530), .B(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g586 ( .A(n_530), .B(n_548), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_530), .B(n_547), .Y(n_614) );
INVx1_ASAP7_75t_L g620 ( .A(n_530), .Y(n_620) );
INVx1_ASAP7_75t_L g637 ( .A(n_530), .Y(n_637) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_530), .Y(n_649) );
INVx2_ASAP7_75t_L g717 ( .A(n_530), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_534), .B(n_535), .Y(n_532) );
INVx2_ASAP7_75t_L g574 ( .A(n_540), .Y(n_574) );
BUFx2_ASAP7_75t_L g671 ( .A(n_540), .Y(n_671) );
AND2x2_ASAP7_75t_L g716 ( .A(n_540), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_558), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_546), .B(n_653), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g739 ( .A1(n_546), .A2(n_715), .B(n_729), .Y(n_739) );
AND2x2_ASAP7_75t_L g764 ( .A(n_546), .B(n_650), .Y(n_764) );
BUFx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g686 ( .A(n_548), .Y(n_686) );
AND2x2_ASAP7_75t_L g715 ( .A(n_548), .B(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_549), .Y(n_599) );
INVx2_ASAP7_75t_L g618 ( .A(n_549), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_549), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
INVx2_ASAP7_75t_L g572 ( .A(n_559), .Y(n_572) );
OR2x2_ASAP7_75t_L g585 ( .A(n_559), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g653 ( .A(n_559), .B(n_649), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_559), .B(n_749), .Y(n_748) );
OR2x2_ASAP7_75t_L g754 ( .A(n_559), .B(n_755), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_559), .B(n_691), .Y(n_766) );
AND2x2_ASAP7_75t_L g645 ( .A(n_560), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g668 ( .A(n_560), .B(n_562), .Y(n_668) );
INVx2_ASAP7_75t_L g580 ( .A(n_561), .Y(n_580) );
AND2x2_ASAP7_75t_L g608 ( .A(n_561), .B(n_581), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_561), .B(n_633), .Y(n_689) );
AND2x2_ASAP7_75t_L g603 ( .A(n_562), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g750 ( .A(n_562), .Y(n_750) );
AND2x2_ASAP7_75t_L g762 ( .A(n_562), .B(n_625), .Y(n_762) );
AND2x2_ASAP7_75t_L g588 ( .A(n_563), .B(n_578), .Y(n_588) );
INVx1_ASAP7_75t_L g683 ( .A(n_563), .Y(n_683) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x4_ASAP7_75t_L g581 ( .A(n_568), .B(n_582), .Y(n_581) );
INVxp67_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_575), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_572), .B(n_619), .Y(n_628) );
OR2x2_ASAP7_75t_L g760 ( .A(n_572), .B(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g677 ( .A(n_573), .B(n_618), .Y(n_677) );
AND2x2_ASAP7_75t_L g685 ( .A(n_573), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g744 ( .A(n_573), .B(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_L g768 ( .A(n_573), .B(n_615), .Y(n_768) );
NOR2xp67_ASAP7_75t_L g726 ( .A(n_574), .B(n_727), .Y(n_726) );
OR2x2_ASAP7_75t_L g755 ( .A(n_574), .B(n_618), .Y(n_755) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND2x1p5_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
AND2x2_ASAP7_75t_L g607 ( .A(n_577), .B(n_608), .Y(n_607) );
INVxp67_ASAP7_75t_L g769 ( .A(n_577), .Y(n_769) );
NOR2x1_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
INVx1_ASAP7_75t_L g604 ( .A(n_580), .Y(n_604) );
AND2x2_ASAP7_75t_L g655 ( .A(n_580), .B(n_588), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_580), .B(n_723), .Y(n_749) );
INVx2_ASAP7_75t_L g594 ( .A(n_581), .Y(n_594) );
INVx3_ASAP7_75t_L g646 ( .A(n_581), .Y(n_646) );
OR2x2_ASAP7_75t_L g674 ( .A(n_581), .B(n_675), .Y(n_674) );
AOI311xp33_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_587), .A3(n_589), .B(n_590), .C(n_601), .Y(n_583) );
O2A1O1Ixp33_ASAP7_75t_L g621 ( .A1(n_584), .A2(n_622), .B(n_624), .C(n_626), .Y(n_621) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_SL g606 ( .A(n_586), .Y(n_606) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g624 ( .A(n_588), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_588), .B(n_604), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_588), .B(n_589), .Y(n_757) );
AND2x2_ASAP7_75t_L g679 ( .A(n_589), .B(n_593), .Y(n_679) );
AOI21xp33_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_595), .B(n_596), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g737 ( .A(n_593), .B(n_625), .Y(n_737) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_594), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g631 ( .A(n_594), .Y(n_631) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
AND2x2_ASAP7_75t_L g622 ( .A(n_598), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g667 ( .A(n_600), .Y(n_667) );
AND2x4_ASAP7_75t_L g729 ( .A(n_600), .B(n_698), .Y(n_729) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AOI222xp33_ASAP7_75t_L g680 ( .A1(n_603), .A2(n_669), .B1(n_681), .B2(n_685), .C1(n_687), .C2(n_691), .Y(n_680) );
A2O1A1Ixp33_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_607), .B(n_609), .C(n_612), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_606), .B(n_650), .Y(n_673) );
INVx1_ASAP7_75t_L g695 ( .A(n_608), .Y(n_695) );
INVx1_ASAP7_75t_L g629 ( .A(n_610), .Y(n_629) );
OR2x2_ASAP7_75t_L g694 ( .A(n_611), .B(n_695), .Y(n_694) );
OAI21xp33_ASAP7_75t_SL g612 ( .A1(n_613), .A2(n_615), .B(n_619), .Y(n_612) );
NAND3xp33_ASAP7_75t_L g630 ( .A(n_613), .B(n_631), .C(n_632), .Y(n_630) );
AOI21xp5_ASAP7_75t_L g728 ( .A1(n_613), .A2(n_650), .B(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_617), .Y(n_670) );
AND2x2_ASAP7_75t_SL g636 ( .A(n_618), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g727 ( .A(n_618), .Y(n_727) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_618), .Y(n_743) );
INVx2_ASAP7_75t_L g701 ( .A(n_619), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_623), .B(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g675 ( .A(n_625), .Y(n_675) );
OAI221xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_629), .B1(n_630), .B2(n_634), .C(n_635), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_629), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_SL g763 ( .A(n_629), .Y(n_763) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g644 ( .A(n_636), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_636), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g702 ( .A(n_636), .B(n_650), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_636), .B(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g735 ( .A(n_636), .B(n_670), .Y(n_735) );
BUFx3_ASAP7_75t_L g698 ( .A(n_637), .Y(n_698) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND5xp2_ASAP7_75t_L g640 ( .A(n_641), .B(n_659), .C(n_680), .D(n_692), .E(n_707), .Y(n_640) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AOI32xp33_ASAP7_75t_L g732 ( .A1(n_644), .A2(n_671), .A3(n_687), .B1(n_733), .B2(n_735), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_646), .B(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_SL g656 ( .A(n_650), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_654), .B1(n_656), .B2(n_657), .Y(n_651) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_666), .B1(n_668), .B2(n_669), .C(n_672), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OR2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g731 ( .A(n_663), .B(n_682), .Y(n_731) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AOI221xp5_ASAP7_75t_L g746 ( .A1(n_668), .A2(n_729), .B1(n_747), .B2(n_752), .C(n_753), .Y(n_746) );
AND2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
INVx2_ASAP7_75t_L g712 ( .A(n_671), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_674), .B1(n_676), .B2(n_678), .Y(n_672) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_684), .Y(n_681) );
INVx1_ASAP7_75t_L g690 ( .A(n_682), .Y(n_690) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
OR2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
AOI222xp33_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_696), .B1(n_700), .B2(n_701), .C1(n_702), .C2(n_703), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_699), .Y(n_696) );
INVxp67_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OAI22xp33_ASAP7_75t_L g747 ( .A1(n_701), .A2(n_748), .B1(n_750), .B2(n_751), .Y(n_747) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_710), .B(n_713), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AOI21xp33_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_718), .B(n_720), .Y(n_713) );
INVx2_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g761 ( .A(n_716), .Y(n_761) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
A2O1A1Ixp33_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_728), .B(n_730), .C(n_732), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
AOI211xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_738), .B(n_740), .C(n_765), .Y(n_736) );
CKINVDCx16_ASAP7_75t_R g741 ( .A(n_737), .Y(n_741) );
INVxp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
OAI211xp5_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_742), .B(n_746), .C(n_758), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
AOI21xp33_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_756), .B(n_757), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_762), .B1(n_763), .B2(n_764), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
AOI21xp33_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_767), .B(n_769), .Y(n_765) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
BUFx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_SL g777 ( .A(n_778), .Y(n_777) );
endmodule