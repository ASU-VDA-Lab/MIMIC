module real_jpeg_24024_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_347, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_347;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_1),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_1),
.A2(n_56),
.B1(n_118),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_118),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_1),
.A2(n_48),
.B1(n_49),
.B2(n_118),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_4),
.A2(n_10),
.B1(n_57),
.B2(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_4),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_130),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_130),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_4),
.A2(n_48),
.B1(n_49),
.B2(n_130),
.Y(n_225)
);

INVx8_ASAP7_75t_SL g65 ( 
.A(n_5),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_6),
.A2(n_71),
.B(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_6),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_6),
.B(n_62),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_L g198 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_127),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_6),
.B(n_44),
.C(n_49),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_6),
.B(n_29),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_6),
.A2(n_101),
.B1(n_219),
.B2(n_225),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_7),
.A2(n_39),
.B1(n_56),
.B2(n_57),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_39),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_7),
.A2(n_39),
.B1(n_48),
.B2(n_49),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_8),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_8),
.A2(n_28),
.B1(n_57),
.B2(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_8),
.A2(n_28),
.B1(n_48),
.B2(n_49),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_11),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_11),
.A2(n_48),
.B1(n_49),
.B2(n_69),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_69),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_69),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_12),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_120),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_12),
.A2(n_48),
.B1(n_49),
.B2(n_120),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_12),
.A2(n_70),
.B1(n_71),
.B2(n_120),
.Y(n_261)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_14),
.A2(n_55),
.B1(n_58),
.B2(n_59),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_58),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_14),
.A2(n_48),
.B1(n_49),
.B2(n_58),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_58),
.Y(n_288)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_15),
.Y(n_104)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_15),
.Y(n_110)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_15),
.Y(n_156)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_15),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_86),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_85),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_78),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_19),
.B(n_78),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_73),
.C(n_74),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_20),
.B(n_342),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_40),
.C(n_52),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_21),
.A2(n_22),
.B1(n_40),
.B2(n_326),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_35),
.Y(n_22)
);

OAI21xp33_ASAP7_75t_L g140 ( 
.A1(n_23),
.A2(n_116),
.B(n_119),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_24),
.A2(n_29),
.B(n_36),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_24),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_25),
.A2(n_26),
.B1(n_30),
.B2(n_34),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_25),
.A2(n_26),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_25),
.A2(n_64),
.B(n_126),
.C(n_143),
.Y(n_142)
);

HAxp5_ASAP7_75t_SL g171 ( 
.A(n_25),
.B(n_127),
.CON(n_171),
.SN(n_171)
);

INVx3_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

NAND3xp33_ASAP7_75t_L g143 ( 
.A(n_26),
.B(n_63),
.C(n_84),
.Y(n_143)
);

OAI32xp33_ASAP7_75t_L g170 ( 
.A1(n_26),
.A2(n_30),
.A3(n_32),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_29),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_29),
.A2(n_36),
.B1(n_162),
.B2(n_171),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_29),
.B(n_38),
.Y(n_265)
);

AO22x1_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_29)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_32),
.B1(n_44),
.B2(n_46),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_31),
.B(n_34),
.Y(n_172)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_32),
.B(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_35),
.A2(n_121),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_36),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_36),
.A2(n_324),
.B(n_325),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_40),
.A2(n_322),
.B1(n_323),
.B2(n_326),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_40),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_47),
.B(n_50),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_42),
.B(n_98),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_42),
.A2(n_51),
.B(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_42),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_42),
.A2(n_180),
.B(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_42),
.A2(n_179),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_42),
.A2(n_178),
.B1(n_179),
.B2(n_199),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_42),
.A2(n_179),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_42),
.A2(n_114),
.B(n_255),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_47),
.Y(n_42)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_47),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_47),
.B(n_99),
.Y(n_114)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_47),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_47),
.B(n_50),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_47),
.B(n_127),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_48),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_48),
.B(n_230),
.Y(n_229)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_52),
.B(n_331),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_60),
.B1(n_62),
.B2(n_68),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_54),
.A2(n_61),
.B(n_79),
.Y(n_319)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_63),
.B1(n_64),
.B2(n_67),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_68),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_60),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_60),
.A2(n_62),
.B1(n_129),
.B2(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_60),
.A2(n_62),
.B1(n_137),
.B2(n_261),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_60),
.A2(n_82),
.B(n_261),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_60),
.A2(n_76),
.B(n_307),
.Y(n_306)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_66),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_61),
.A2(n_123),
.B1(n_124),
.B2(n_128),
.Y(n_122)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_73),
.A2(n_74),
.B1(n_75),
.B2(n_343),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_73),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_83),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_84),
.B(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_339),
.B(n_344),
.Y(n_86)
);

OAI321xp33_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_315),
.A3(n_334),
.B1(n_337),
.B2(n_338),
.C(n_347),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_293),
.B(n_314),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_270),
.B(n_292),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_163),
.B(n_245),
.C(n_269),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_148),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_92),
.B(n_148),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_133),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_111),
.B1(n_131),
.B2(n_132),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_94),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_94),
.B(n_132),
.C(n_133),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_100),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_95),
.B(n_100),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_96),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_97),
.B(n_300),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_105),
.B(n_107),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_101),
.A2(n_107),
.B(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_101),
.A2(n_209),
.B(n_210),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_101),
.A2(n_216),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_101),
.A2(n_174),
.B(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_102),
.A2(n_103),
.B1(n_106),
.B2(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_102),
.B(n_108),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_102),
.A2(n_215),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_104),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_115),
.C(n_122),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_112),
.A2(n_113),
.B1(n_115),
.B2(n_151),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_119),
.B2(n_121),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_116),
.A2(n_117),
.B1(n_121),
.B2(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_116),
.A2(n_264),
.B(n_265),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_116),
.A2(n_121),
.B1(n_288),
.B2(n_302),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_122),
.B(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_127),
.B(n_156),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_141),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_139),
.B2(n_140),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_136),
.B(n_139),
.C(n_141),
.Y(n_267)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_142),
.A2(n_144),
.B1(n_145),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_147),
.A2(n_156),
.B(n_157),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.C(n_154),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_149),
.B(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_152),
.B(n_154),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.C(n_160),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_155),
.A2(n_158),
.B1(n_159),
.B2(n_185),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_155),
.Y(n_185)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_156),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_156),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_157),
.B(n_210),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_240),
.B(n_244),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_193),
.B(n_239),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_181),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_168),
.B(n_181),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_176),
.C(n_177),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_169),
.B(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_173),
.Y(n_188)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_176),
.B(n_177),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_186),
.B2(n_187),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_182),
.B(n_189),
.C(n_192),
.Y(n_241)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_192),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_188),
.Y(n_192)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_191),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_234),
.B(n_238),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_212),
.B(n_233),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_202),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_196),
.B(n_202),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_200),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_208),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_207),
.C(n_208),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_206),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_209),
.Y(n_217)
);

AOI21xp33_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_221),
.B(n_232),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_220),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_220),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_227),
.B(n_231),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_223),
.B(n_224),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_235),
.B(n_236),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_241),
.B(n_242),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_247),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_267),
.B2(n_268),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_257),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_257),
.C(n_268),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_256),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_256),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_253),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_266),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_262),
.B2(n_263),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_260),
.B(n_262),
.C(n_266),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_265),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_267),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_271),
.B(n_272),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_291),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_281),
.B1(n_289),
.B2(n_290),
.Y(n_273)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_274),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_290),
.C(n_291),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_276),
.B(n_277),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_277),
.A2(n_278),
.B1(n_306),
.B2(n_308),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_277),
.A2(n_308),
.B(n_309),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_281),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_282),
.B(n_285),
.C(n_286),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_294),
.B(n_295),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_312),
.B2(n_313),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_304),
.B1(n_310),
.B2(n_311),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_298),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_298),
.B(n_311),
.C(n_313),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_301),
.B(n_303),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_301),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_302),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_317),
.C(n_327),
.Y(n_316)
);

FAx1_ASAP7_75t_SL g336 ( 
.A(n_303),
.B(n_317),
.CI(n_327),
.CON(n_336),
.SN(n_336)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_304),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_309),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_306),
.Y(n_308)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_312),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_328),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_316),
.B(n_328),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_319),
.B1(n_320),
.B2(n_321),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_318),
.A2(n_319),
.B1(n_330),
.B2(n_332),
.Y(n_329)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_319),
.B(n_323),
.C(n_326),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_319),
.B(n_332),
.C(n_333),
.Y(n_340)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_333),
.Y(n_328)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_330),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_335),
.B(n_336),
.Y(n_337)
);

BUFx24_ASAP7_75t_SL g346 ( 
.A(n_336),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_340),
.B(n_341),
.Y(n_344)
);


endmodule