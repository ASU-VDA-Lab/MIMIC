module fake_netlist_6_585_n_1689 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1689);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1689;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_55),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_19),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_27),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_10),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_129),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_74),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_138),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_70),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_119),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_57),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_93),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_53),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_117),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_135),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_122),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_21),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_30),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_9),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_50),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_125),
.Y(n_178)
);

BUFx10_ASAP7_75t_L g179 ( 
.A(n_139),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_128),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_154),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_46),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_27),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_9),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_47),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_11),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_107),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_145),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_8),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_84),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_127),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_148),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_21),
.Y(n_193)
);

BUFx10_ASAP7_75t_L g194 ( 
.A(n_114),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_47),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_65),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_26),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_153),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_109),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_16),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_118),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_56),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_46),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_113),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_142),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_68),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_131),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_100),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_150),
.Y(n_209)
);

BUFx10_ASAP7_75t_L g210 ( 
.A(n_49),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_40),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_98),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_0),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_7),
.Y(n_214)
);

BUFx8_ASAP7_75t_SL g215 ( 
.A(n_103),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_44),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_110),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_12),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_39),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g220 ( 
.A(n_38),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_11),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_75),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_120),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_14),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_81),
.Y(n_225)
);

INVx4_ASAP7_75t_R g226 ( 
.A(n_85),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_112),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_62),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_26),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_72),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_10),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_92),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_20),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_4),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_61),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_35),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_22),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_30),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_144),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_16),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_37),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_14),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_108),
.Y(n_243)
);

BUFx8_ASAP7_75t_SL g244 ( 
.A(n_97),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_141),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_104),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_22),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_66),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_40),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_137),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_99),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_126),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_77),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_39),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_51),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_82),
.Y(n_256)
);

BUFx8_ASAP7_75t_SL g257 ( 
.A(n_45),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_52),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_80),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_76),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_19),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_96),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_78),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_4),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_87),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_28),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_71),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_95),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_20),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_7),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_140),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_69),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_23),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_134),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_41),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_116),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_88),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_58),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_24),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_23),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_106),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_28),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_67),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_123),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_37),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_17),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_5),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_91),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_50),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_133),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_42),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_29),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_86),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_105),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_35),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_90),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_156),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_132),
.Y(n_298)
);

BUFx2_ASAP7_75t_SL g299 ( 
.A(n_38),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_29),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_73),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_64),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_17),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_33),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_94),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_8),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_48),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_49),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_149),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_36),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_124),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_237),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_220),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_300),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_215),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_169),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_244),
.Y(n_317)
);

BUFx6f_ASAP7_75t_SL g318 ( 
.A(n_179),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_220),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_220),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_257),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_220),
.B(n_0),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_210),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_161),
.B(n_190),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_228),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_175),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_192),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_199),
.B(n_283),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_178),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_251),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_253),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_188),
.Y(n_332)
);

NOR2xp67_ASAP7_75t_L g333 ( 
.A(n_160),
.B(n_1),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_220),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_220),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_243),
.B(n_157),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_220),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_198),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_201),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_220),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_202),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_204),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_209),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_252),
.Y(n_344)
);

OR2x2_ASAP7_75t_L g345 ( 
.A(n_186),
.B(n_1),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_174),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_174),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_212),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_296),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_217),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_243),
.B(n_2),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_188),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_174),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_222),
.Y(n_354)
);

INVxp33_ASAP7_75t_L g355 ( 
.A(n_189),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_225),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_159),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_223),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_232),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_174),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_245),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_246),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_174),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_254),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_254),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_254),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_254),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_248),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_250),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_254),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_259),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_225),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_256),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_264),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_260),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_264),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_262),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_263),
.Y(n_378)
);

CKINVDCx14_ASAP7_75t_R g379 ( 
.A(n_210),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_264),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_271),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_272),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_264),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_264),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_159),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_157),
.B(n_2),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_256),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_325),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_358),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_325),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_346),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_325),
.Y(n_392)
);

AND2x6_ASAP7_75t_L g393 ( 
.A(n_325),
.B(n_207),
.Y(n_393)
);

AND3x2_ASAP7_75t_L g394 ( 
.A(n_324),
.B(n_208),
.C(n_207),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_328),
.B(n_179),
.Y(n_395)
);

NAND2x1p5_ASAP7_75t_L g396 ( 
.A(n_386),
.B(n_165),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_346),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_359),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_347),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_325),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_325),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_332),
.B(n_175),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_313),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_361),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_313),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_352),
.B(n_195),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_347),
.B(n_208),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_336),
.B(n_163),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_319),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_319),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_353),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_353),
.B(n_255),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_360),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_372),
.B(n_195),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_373),
.B(n_163),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_320),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_360),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_363),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_320),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_387),
.B(n_200),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_334),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_368),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_363),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_351),
.B(n_164),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_364),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_364),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_365),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_365),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_327),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_334),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_366),
.B(n_164),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_331),
.B(n_314),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_366),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_356),
.B(n_326),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_367),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_367),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_370),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_370),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_374),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_374),
.Y(n_440)
);

INVx6_ASAP7_75t_L g441 ( 
.A(n_356),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_312),
.A2(n_182),
.B1(n_287),
.B2(n_197),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_356),
.B(n_200),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_376),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_335),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_335),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_326),
.B(n_255),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_376),
.B(n_166),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_337),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_380),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_337),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_380),
.Y(n_452)
);

XOR2x2_ASAP7_75t_SL g453 ( 
.A(n_322),
.B(n_214),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_383),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_340),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_383),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_384),
.B(n_166),
.Y(n_457)
);

OA21x2_ASAP7_75t_L g458 ( 
.A1(n_340),
.A2(n_219),
.B(n_160),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_441),
.B(n_338),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_427),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_395),
.B(n_339),
.Y(n_461)
);

NOR3xp33_ASAP7_75t_L g462 ( 
.A(n_395),
.B(n_323),
.C(n_357),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_441),
.B(n_424),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g464 ( 
.A1(n_396),
.A2(n_333),
.B1(n_345),
.B2(n_291),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_403),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_396),
.B(n_341),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_389),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_396),
.B(n_342),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_396),
.A2(n_333),
.B1(n_345),
.B2(n_219),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_443),
.B(n_384),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_396),
.A2(n_350),
.B1(n_382),
.B2(n_381),
.Y(n_471)
);

INVx4_ASAP7_75t_L g472 ( 
.A(n_421),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_441),
.B(n_343),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_427),
.Y(n_474)
);

BUFx10_ASAP7_75t_L g475 ( 
.A(n_429),
.Y(n_475)
);

NAND2xp33_ASAP7_75t_L g476 ( 
.A(n_424),
.B(n_228),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_390),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_458),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_458),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_403),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_390),
.Y(n_481)
);

BUFx10_ASAP7_75t_L g482 ( 
.A(n_429),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_441),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_415),
.B(n_348),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_458),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_403),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_441),
.B(n_408),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_403),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_458),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_458),
.Y(n_490)
);

NAND2xp33_ASAP7_75t_L g491 ( 
.A(n_393),
.B(n_228),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_458),
.Y(n_492)
);

INVx4_ASAP7_75t_L g493 ( 
.A(n_421),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_415),
.B(n_354),
.Y(n_494)
);

BUFx8_ASAP7_75t_SL g495 ( 
.A(n_389),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_390),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_442),
.B(n_316),
.Y(n_497)
);

NAND2xp33_ASAP7_75t_L g498 ( 
.A(n_393),
.B(n_228),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_408),
.B(n_362),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_441),
.B(n_369),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_432),
.A2(n_378),
.B1(n_377),
.B2(n_375),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_443),
.B(n_158),
.Y(n_502)
);

BUFx10_ASAP7_75t_L g503 ( 
.A(n_432),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_390),
.Y(n_504)
);

NAND2xp33_ASAP7_75t_L g505 ( 
.A(n_393),
.B(n_228),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_409),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_409),
.Y(n_507)
);

A2O1A1Ixp33_ASAP7_75t_L g508 ( 
.A1(n_405),
.A2(n_276),
.B(n_355),
.C(n_291),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_409),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_390),
.Y(n_510)
);

OA22x2_ASAP7_75t_L g511 ( 
.A1(n_394),
.A2(n_385),
.B1(n_216),
.B2(n_221),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_409),
.Y(n_512)
);

AND3x2_ASAP7_75t_L g513 ( 
.A(n_447),
.B(n_276),
.C(n_180),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_441),
.B(n_371),
.Y(n_514)
);

NAND3xp33_ASAP7_75t_SL g515 ( 
.A(n_442),
.B(n_269),
.C(n_183),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_453),
.B(n_434),
.Y(n_516)
);

BUFx6f_ASAP7_75t_SL g517 ( 
.A(n_407),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_410),
.Y(n_518)
);

NOR2x1p5_ASAP7_75t_L g519 ( 
.A(n_398),
.B(n_315),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_398),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_410),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_405),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_405),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_434),
.B(n_379),
.Y(n_524)
);

AOI21x1_ASAP7_75t_L g525 ( 
.A1(n_407),
.A2(n_187),
.B(n_171),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_402),
.A2(n_261),
.B1(n_249),
.B2(n_286),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_390),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_405),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_434),
.B(n_317),
.Y(n_529)
);

BUFx10_ASAP7_75t_L g530 ( 
.A(n_404),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_443),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_405),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_404),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_410),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_402),
.B(n_229),
.Y(n_535)
);

AND2x6_ASAP7_75t_L g536 ( 
.A(n_447),
.B(n_230),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_410),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_453),
.B(n_321),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_427),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_L g540 ( 
.A(n_393),
.B(n_230),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_427),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_390),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_421),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_416),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_430),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_390),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_430),
.Y(n_547)
);

AND2x6_ASAP7_75t_L g548 ( 
.A(n_447),
.B(n_230),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_421),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_416),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_416),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_416),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_402),
.B(n_206),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_421),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_421),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_416),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_430),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_419),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_430),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_419),
.Y(n_560)
);

CKINVDCx6p67_ASAP7_75t_R g561 ( 
.A(n_406),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_419),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_422),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_421),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_419),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_406),
.A2(n_233),
.B1(n_236),
.B2(n_273),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_446),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_419),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_406),
.B(n_318),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_446),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_421),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_446),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_414),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_414),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_393),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_422),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_400),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_400),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_446),
.Y(n_579)
);

OR2x6_ASAP7_75t_L g580 ( 
.A(n_420),
.B(n_299),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_449),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_453),
.B(n_179),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_420),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_449),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_445),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_400),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_407),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_431),
.B(n_194),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_407),
.A2(n_303),
.B1(n_242),
.B2(n_230),
.Y(n_589)
);

INVx6_ASAP7_75t_L g590 ( 
.A(n_407),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_445),
.Y(n_591)
);

OR2x6_ASAP7_75t_L g592 ( 
.A(n_431),
.B(n_196),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_445),
.Y(n_593)
);

AND2x6_ASAP7_75t_L g594 ( 
.A(n_445),
.B(n_230),
.Y(n_594)
);

NOR2x1p5_ASAP7_75t_L g595 ( 
.A(n_448),
.B(n_162),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_400),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_449),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_449),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_445),
.Y(n_599)
);

NOR2x1p5_ASAP7_75t_L g600 ( 
.A(n_448),
.B(n_162),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_457),
.B(n_194),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_400),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_451),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_SL g604 ( 
.A(n_407),
.B(n_318),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_451),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_412),
.Y(n_606)
);

AND2x2_ASAP7_75t_SL g607 ( 
.A(n_476),
.B(n_499),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_484),
.B(n_451),
.Y(n_608)
);

AOI22x1_ASAP7_75t_SL g609 ( 
.A1(n_576),
.A2(n_533),
.B1(n_563),
.B2(n_520),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_573),
.B(n_455),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_529),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_573),
.B(n_455),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_583),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_494),
.B(n_455),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_574),
.B(n_394),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_574),
.B(n_583),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_L g617 ( 
.A1(n_478),
.A2(n_392),
.B(n_388),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_531),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_470),
.B(n_601),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_465),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_470),
.B(n_412),
.Y(n_621)
);

OR2x2_ASAP7_75t_L g622 ( 
.A(n_553),
.B(n_176),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_587),
.B(n_412),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_531),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_601),
.B(n_412),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_465),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_580),
.B(n_176),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_599),
.Y(n_628)
);

NOR3xp33_ASAP7_75t_L g629 ( 
.A(n_582),
.B(n_203),
.C(n_193),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_L g630 ( 
.A(n_536),
.B(n_274),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_587),
.B(n_412),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_590),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_460),
.Y(n_633)
);

INVxp33_ASAP7_75t_L g634 ( 
.A(n_497),
.Y(n_634)
);

BUFx6f_ASAP7_75t_SL g635 ( 
.A(n_475),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_503),
.B(n_167),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_587),
.B(n_205),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_474),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_539),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_541),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_478),
.A2(n_265),
.B1(n_227),
.B2(n_258),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_590),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_479),
.B(n_485),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_479),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_587),
.B(n_267),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_485),
.B(n_397),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_535),
.Y(n_647)
);

INVx2_ASAP7_75t_SL g648 ( 
.A(n_535),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_595),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_600),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_502),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_489),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_590),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_561),
.B(n_329),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_489),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_590),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_516),
.A2(n_330),
.B1(n_344),
.B2(n_349),
.Y(n_657)
);

INVx8_ASAP7_75t_L g658 ( 
.A(n_580),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_502),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_490),
.B(n_397),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_490),
.B(n_399),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_587),
.B(n_268),
.Y(n_662)
);

NAND2x1p5_ASAP7_75t_L g663 ( 
.A(n_575),
.B(n_277),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_606),
.B(n_463),
.Y(n_664)
);

OR2x6_ASAP7_75t_L g665 ( 
.A(n_580),
.B(n_278),
.Y(n_665)
);

INVxp67_ASAP7_75t_SL g666 ( 
.A(n_492),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_492),
.B(n_399),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_522),
.Y(n_668)
);

NAND2xp33_ASAP7_75t_L g669 ( 
.A(n_536),
.B(n_284),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_487),
.B(n_411),
.Y(n_670)
);

O2A1O1Ixp33_ASAP7_75t_L g671 ( 
.A1(n_476),
.A2(n_435),
.B(n_454),
.C(n_452),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_522),
.B(n_411),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_606),
.B(n_281),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_599),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_523),
.B(n_413),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g676 ( 
.A1(n_523),
.A2(n_388),
.B(n_392),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_503),
.B(n_167),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_480),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_606),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_606),
.B(n_575),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_528),
.B(n_413),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_486),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_561),
.B(n_210),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_483),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_486),
.Y(n_685)
);

NOR2x1p5_ASAP7_75t_L g686 ( 
.A(n_515),
.B(n_177),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_577),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_528),
.B(n_425),
.Y(n_688)
);

NAND3x1_ASAP7_75t_L g689 ( 
.A(n_462),
.B(n_311),
.C(n_309),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_580),
.Y(n_690)
);

NOR2x1p5_ASAP7_75t_L g691 ( 
.A(n_520),
.B(n_177),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_575),
.B(n_293),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_592),
.A2(n_294),
.B1(n_290),
.B2(n_168),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_532),
.B(n_425),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_503),
.B(n_211),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_488),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_488),
.Y(n_697)
);

NAND3xp33_ASAP7_75t_L g698 ( 
.A(n_464),
.B(n_231),
.C(n_224),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_544),
.B(n_426),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_501),
.B(n_168),
.Y(n_700)
);

BUFx12f_ASAP7_75t_L g701 ( 
.A(n_530),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_550),
.B(n_551),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_550),
.B(n_426),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_R g704 ( 
.A(n_533),
.B(n_563),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_466),
.B(n_170),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_551),
.B(n_428),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_502),
.B(n_298),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_506),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_513),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_552),
.B(n_428),
.Y(n_710)
);

AO221x1_ASAP7_75t_L g711 ( 
.A1(n_577),
.A2(n_302),
.B1(n_318),
.B2(n_226),
.C(n_194),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_506),
.Y(n_712)
);

INVxp67_ASAP7_75t_L g713 ( 
.A(n_524),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_471),
.B(n_170),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_507),
.Y(n_715)
);

A2O1A1Ixp33_ASAP7_75t_L g716 ( 
.A1(n_469),
.A2(n_566),
.B(n_526),
.C(n_569),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_556),
.B(n_558),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_511),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_467),
.B(n_184),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_468),
.B(n_172),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_507),
.Y(n_721)
);

O2A1O1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_508),
.A2(n_436),
.B(n_454),
.C(n_452),
.Y(n_722)
);

A2O1A1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_556),
.A2(n_234),
.B(n_184),
.C(n_185),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_461),
.B(n_592),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_483),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_475),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_592),
.B(n_172),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_558),
.B(n_173),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_577),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_560),
.B(n_181),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_511),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_560),
.B(n_181),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_562),
.B(n_191),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_592),
.B(n_588),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_562),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_565),
.B(n_433),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_509),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_565),
.B(n_433),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_509),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_475),
.B(n_213),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_SL g741 ( 
.A(n_482),
.B(n_191),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_538),
.B(n_235),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_578),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_568),
.B(n_235),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_511),
.A2(n_239),
.B1(n_290),
.B2(n_294),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_568),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_585),
.B(n_435),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_585),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_593),
.B(n_239),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_SL g750 ( 
.A(n_482),
.B(n_288),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_512),
.Y(n_751)
);

NOR2xp67_ASAP7_75t_SL g752 ( 
.A(n_481),
.B(n_288),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_593),
.B(n_297),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_459),
.B(n_436),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_512),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_578),
.B(n_297),
.Y(n_756)
);

NAND3xp33_ASAP7_75t_L g757 ( 
.A(n_589),
.B(n_218),
.C(n_240),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_591),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_473),
.B(n_301),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_500),
.B(n_301),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_518),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_518),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_514),
.B(n_305),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_578),
.B(n_438),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_497),
.B(n_185),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_482),
.B(n_241),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_517),
.A2(n_305),
.B1(n_456),
.B2(n_444),
.Y(n_767)
);

O2A1O1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_491),
.A2(n_438),
.B(n_450),
.C(n_439),
.Y(n_768)
);

OAI221xp5_ASAP7_75t_L g769 ( 
.A1(n_604),
.A2(n_247),
.B1(n_266),
.B2(n_270),
.C(n_275),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_521),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_619),
.B(n_536),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_R g772 ( 
.A(n_701),
.B(n_576),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_719),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_611),
.B(n_586),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_680),
.A2(n_564),
.B(n_493),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_613),
.Y(n_776)
);

NAND3xp33_ASAP7_75t_L g777 ( 
.A(n_700),
.B(n_742),
.C(n_616),
.Y(n_777)
);

O2A1O1Ixp33_ASAP7_75t_SL g778 ( 
.A1(n_692),
.A2(n_605),
.B(n_586),
.C(n_602),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_668),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_680),
.A2(n_543),
.B(n_564),
.Y(n_780)
);

OAI21xp5_ASAP7_75t_L g781 ( 
.A1(n_643),
.A2(n_603),
.B(n_521),
.Y(n_781)
);

BUFx12f_ASAP7_75t_L g782 ( 
.A(n_649),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_L g783 ( 
.A1(n_617),
.A2(n_603),
.B(n_534),
.Y(n_783)
);

OAI21xp33_ASAP7_75t_L g784 ( 
.A1(n_700),
.A2(n_289),
.B(n_310),
.Y(n_784)
);

INVxp67_ASAP7_75t_SL g785 ( 
.A(n_644),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_664),
.A2(n_472),
.B(n_564),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_616),
.B(n_586),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_608),
.B(n_536),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_614),
.B(n_536),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_607),
.B(n_548),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_607),
.B(n_548),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_735),
.Y(n_792)
);

BUFx12f_ASAP7_75t_L g793 ( 
.A(n_650),
.Y(n_793)
);

INVx4_ASAP7_75t_L g794 ( 
.A(n_628),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_625),
.B(n_596),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_713),
.B(n_596),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_678),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_623),
.A2(n_472),
.B(n_543),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_647),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_623),
.A2(n_472),
.B(n_543),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_628),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_648),
.B(n_596),
.Y(n_802)
);

NOR3xp33_ASAP7_75t_L g803 ( 
.A(n_742),
.B(n_505),
.C(n_491),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_666),
.B(n_548),
.Y(n_804)
);

NOR2xp67_ASAP7_75t_SL g805 ( 
.A(n_726),
.B(n_628),
.Y(n_805)
);

AOI21xp33_ASAP7_75t_L g806 ( 
.A1(n_705),
.A2(n_720),
.B(n_727),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_631),
.A2(n_493),
.B(n_481),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_631),
.A2(n_493),
.B(n_481),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_670),
.A2(n_504),
.B(n_496),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_644),
.B(n_548),
.Y(n_810)
);

AO21x1_ASAP7_75t_L g811 ( 
.A1(n_705),
.A2(n_720),
.B(n_724),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_726),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_652),
.B(n_548),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_SL g814 ( 
.A(n_635),
.B(n_530),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_628),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_746),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_621),
.A2(n_504),
.B(n_496),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_754),
.B(n_602),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_646),
.A2(n_504),
.B(n_496),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_636),
.B(n_602),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_660),
.A2(n_504),
.B(n_496),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_674),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_661),
.A2(n_527),
.B(n_542),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_652),
.B(n_655),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_708),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_667),
.A2(n_527),
.B(n_542),
.Y(n_826)
);

NOR3xp33_ASAP7_75t_L g827 ( 
.A(n_714),
.B(n_498),
.C(n_505),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_610),
.A2(n_527),
.B(n_542),
.Y(n_828)
);

AND2x4_ASAP7_75t_L g829 ( 
.A(n_618),
.B(n_519),
.Y(n_829)
);

INVxp67_ASAP7_75t_L g830 ( 
.A(n_615),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_610),
.A2(n_527),
.B(n_542),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_655),
.B(n_548),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_612),
.A2(n_481),
.B(n_527),
.Y(n_833)
);

OAI22xp5_ASAP7_75t_L g834 ( 
.A1(n_641),
.A2(n_517),
.B1(n_554),
.B2(n_555),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_641),
.B(n_549),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_759),
.B(n_549),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_612),
.A2(n_481),
.B(n_542),
.Y(n_837)
);

AOI22x1_ASAP7_75t_L g838 ( 
.A1(n_687),
.A2(n_555),
.B1(n_554),
.B2(n_571),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_708),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_748),
.Y(n_840)
);

INVx3_ASAP7_75t_SL g841 ( 
.A(n_658),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_636),
.B(n_530),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_759),
.B(n_554),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_692),
.A2(n_555),
.B(n_571),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_663),
.A2(n_510),
.B(n_477),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_760),
.B(n_534),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_663),
.A2(n_676),
.B(n_754),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_760),
.B(n_537),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_763),
.B(n_545),
.Y(n_849)
);

OAI321xp33_ASAP7_75t_L g850 ( 
.A1(n_714),
.A2(n_525),
.A3(n_439),
.B1(n_450),
.B2(n_456),
.C(n_444),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_734),
.B(n_477),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_677),
.B(n_545),
.Y(n_852)
);

O2A1O1Ixp5_ASAP7_75t_L g853 ( 
.A1(n_637),
.A2(n_525),
.B(n_597),
.C(n_567),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_624),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_763),
.B(n_547),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_717),
.A2(n_598),
.B(n_597),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_718),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_712),
.Y(n_858)
);

NOR2x1p5_ASAP7_75t_L g859 ( 
.A(n_765),
.B(n_234),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_734),
.B(n_510),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_716),
.B(n_731),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_717),
.A2(n_559),
.B(n_584),
.Y(n_862)
);

OAI21xp5_ASAP7_75t_L g863 ( 
.A1(n_702),
.A2(n_559),
.B(n_584),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_642),
.A2(n_510),
.B(n_546),
.Y(n_864)
);

NAND3xp33_ASAP7_75t_L g865 ( 
.A(n_677),
.B(n_280),
.C(n_279),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_674),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_656),
.A2(n_546),
.B(n_540),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_724),
.B(n_546),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_651),
.A2(n_659),
.B1(n_727),
.B2(n_653),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_679),
.B(n_547),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_618),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_716),
.B(n_557),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_633),
.B(n_557),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_690),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_638),
.B(n_570),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_679),
.A2(n_540),
.B(n_498),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_622),
.B(n_572),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_654),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_764),
.A2(n_581),
.B(n_579),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_695),
.B(n_238),
.Y(n_880)
);

OR2x6_ASAP7_75t_L g881 ( 
.A(n_658),
.B(n_495),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_627),
.B(n_572),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_639),
.B(n_579),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_715),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_640),
.B(n_581),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_683),
.B(n_289),
.Y(n_886)
);

AO21x1_ASAP7_75t_L g887 ( 
.A1(n_637),
.A2(n_423),
.B(n_391),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_653),
.A2(n_392),
.B(n_388),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_740),
.B(n_766),
.Y(n_889)
);

OR2x2_ASAP7_75t_L g890 ( 
.A(n_657),
.B(n_238),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_741),
.B(n_517),
.Y(n_891)
);

AO21x1_ASAP7_75t_L g892 ( 
.A1(n_645),
.A2(n_423),
.B(n_456),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_721),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_753),
.B(n_391),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_758),
.B(n_391),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_687),
.B(n_444),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_750),
.B(n_282),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_684),
.A2(n_392),
.B(n_401),
.Y(n_898)
);

OAI22xp5_ASAP7_75t_L g899 ( 
.A1(n_632),
.A2(n_417),
.B1(n_440),
.B2(n_437),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_729),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_684),
.A2(n_401),
.B(n_440),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_684),
.A2(n_401),
.B(n_440),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_729),
.B(n_437),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_R g904 ( 
.A(n_635),
.B(n_658),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_743),
.Y(n_905)
);

O2A1O1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_723),
.A2(n_733),
.B(n_732),
.C(n_730),
.Y(n_906)
);

NAND3xp33_ASAP7_75t_L g907 ( 
.A(n_693),
.B(n_285),
.C(n_292),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_743),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_704),
.B(n_285),
.Y(n_909)
);

NOR2xp67_ASAP7_75t_L g910 ( 
.A(n_769),
.B(n_83),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_684),
.A2(n_401),
.B(n_423),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_674),
.B(n_417),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_704),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_698),
.B(n_292),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_721),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_761),
.Y(n_916)
);

OAI21xp33_ASAP7_75t_L g917 ( 
.A1(n_745),
.A2(n_295),
.B(n_304),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_709),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_725),
.A2(n_418),
.B(n_417),
.Y(n_919)
);

NOR2xp67_ASAP7_75t_L g920 ( 
.A(n_757),
.B(n_63),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_707),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_691),
.B(n_295),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_SL g923 ( 
.A(n_634),
.B(n_665),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_632),
.B(n_418),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_707),
.B(n_418),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_728),
.B(n_304),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_665),
.B(n_59),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_674),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_725),
.A2(n_594),
.B(n_393),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_686),
.B(n_306),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_665),
.Y(n_931)
);

INVx3_ASAP7_75t_L g932 ( 
.A(n_725),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_725),
.B(n_310),
.Y(n_933)
);

NOR2xp67_ASAP7_75t_L g934 ( 
.A(n_756),
.B(n_54),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_762),
.Y(n_935)
);

O2A1O1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_723),
.A2(n_308),
.B(n_307),
.C(n_306),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_756),
.A2(n_307),
.B1(n_308),
.B2(n_594),
.Y(n_937)
);

CKINVDCx10_ASAP7_75t_R g938 ( 
.A(n_609),
.Y(n_938)
);

NAND3xp33_ASAP7_75t_L g939 ( 
.A(n_629),
.B(n_3),
.C(n_5),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_770),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_728),
.B(n_152),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_770),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_730),
.B(n_151),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_672),
.Y(n_944)
);

A2O1A1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_732),
.A2(n_594),
.B(n_6),
.C(n_12),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_733),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_675),
.A2(n_393),
.B(n_147),
.Y(n_947)
);

OA21x2_ASAP7_75t_L g948 ( 
.A1(n_790),
.A2(n_706),
.B(n_681),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_871),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_944),
.B(n_744),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_857),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_782),
.Y(n_952)
);

AOI21x1_ASAP7_75t_L g953 ( 
.A1(n_868),
.A2(n_703),
.B(n_699),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_857),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_847),
.A2(n_630),
.B(n_669),
.Y(n_955)
);

AOI21x1_ASAP7_75t_L g956 ( 
.A1(n_868),
.A2(n_747),
.B(n_736),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_822),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_779),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_806),
.A2(n_749),
.B(n_744),
.C(n_662),
.Y(n_959)
);

NAND3xp33_ASAP7_75t_L g960 ( 
.A(n_777),
.B(n_914),
.C(n_926),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_830),
.A2(n_749),
.B(n_767),
.C(n_673),
.Y(n_961)
);

AOI21x1_ASAP7_75t_L g962 ( 
.A1(n_836),
.A2(n_688),
.B(n_694),
.Y(n_962)
);

INVxp67_ASAP7_75t_L g963 ( 
.A(n_773),
.Y(n_963)
);

OR2x6_ASAP7_75t_SL g964 ( 
.A(n_907),
.B(n_689),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_830),
.B(n_710),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_775),
.A2(n_738),
.B(n_755),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_842),
.B(n_620),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_942),
.Y(n_968)
);

A2O1A1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_906),
.A2(n_722),
.B(n_768),
.C(n_671),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_SL g970 ( 
.A1(n_842),
.A2(n_711),
.B1(n_682),
.B2(n_685),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_776),
.B(n_751),
.Y(n_971)
);

O2A1O1Ixp5_ASAP7_75t_L g972 ( 
.A1(n_811),
.A2(n_752),
.B(n_739),
.C(n_737),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_877),
.B(n_697),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_874),
.Y(n_974)
);

OAI21xp33_ASAP7_75t_L g975 ( 
.A1(n_784),
.A2(n_696),
.B(n_626),
.Y(n_975)
);

O2A1O1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_914),
.A2(n_3),
.B(n_6),
.C(n_13),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_L g977 ( 
.A1(n_861),
.A2(n_13),
.B1(n_15),
.B2(n_18),
.Y(n_977)
);

OAI21x1_ASAP7_75t_L g978 ( 
.A1(n_838),
.A2(n_393),
.B(n_146),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_772),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_877),
.B(n_787),
.Y(n_980)
);

INVx4_ASAP7_75t_L g981 ( 
.A(n_822),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_822),
.Y(n_982)
);

INVx4_ASAP7_75t_L g983 ( 
.A(n_822),
.Y(n_983)
);

O2A1O1Ixp5_ASAP7_75t_L g984 ( 
.A1(n_852),
.A2(n_111),
.B(n_143),
.C(n_136),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_921),
.B(n_130),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_918),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_926),
.A2(n_15),
.B(n_18),
.C(n_24),
.Y(n_987)
);

NAND2x1p5_ASAP7_75t_L g988 ( 
.A(n_805),
.B(n_115),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_SL g989 ( 
.A1(n_791),
.A2(n_102),
.B(n_101),
.C(n_89),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_871),
.Y(n_990)
);

AOI22xp5_ASAP7_75t_L g991 ( 
.A1(n_889),
.A2(n_393),
.B1(n_79),
.B2(n_60),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_787),
.B(n_25),
.Y(n_992)
);

BUFx10_ASAP7_75t_L g993 ( 
.A(n_829),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_942),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_774),
.B(n_25),
.Y(n_995)
);

AOI22xp33_ASAP7_75t_L g996 ( 
.A1(n_941),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_774),
.B(n_31),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_799),
.B(n_946),
.Y(n_998)
);

AOI22xp33_ASAP7_75t_L g999 ( 
.A1(n_941),
.A2(n_32),
.B1(n_34),
.B2(n_36),
.Y(n_999)
);

INVx1_ASAP7_75t_SL g1000 ( 
.A(n_946),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_824),
.A2(n_34),
.B1(n_41),
.B2(n_42),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_SL g1002 ( 
.A1(n_852),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_1002)
);

NOR2x1_ASAP7_75t_L g1003 ( 
.A(n_913),
.B(n_43),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_882),
.A2(n_48),
.B(n_820),
.C(n_796),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_882),
.B(n_796),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_780),
.A2(n_843),
.B(n_800),
.Y(n_1006)
);

AOI22x1_ASAP7_75t_L g1007 ( 
.A1(n_867),
.A2(n_809),
.B1(n_876),
.B2(n_905),
.Y(n_1007)
);

INVx4_ASAP7_75t_L g1008 ( 
.A(n_866),
.Y(n_1008)
);

AOI21x1_ASAP7_75t_L g1009 ( 
.A1(n_795),
.A2(n_872),
.B(n_848),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_866),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_820),
.B(n_792),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_880),
.B(n_886),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_816),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_840),
.B(n_802),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_909),
.B(n_921),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_866),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_936),
.A2(n_897),
.B(n_933),
.C(n_945),
.Y(n_1017)
);

INVx2_ASAP7_75t_SL g1018 ( 
.A(n_874),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_866),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_846),
.B(n_849),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_SL g1021 ( 
.A1(n_890),
.A2(n_878),
.B1(n_931),
.B2(n_881),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_799),
.B(n_930),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_798),
.A2(n_817),
.B(n_819),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_916),
.Y(n_1024)
);

INVx4_ASAP7_75t_L g1025 ( 
.A(n_928),
.Y(n_1025)
);

OAI21xp33_ASAP7_75t_SL g1026 ( 
.A1(n_835),
.A2(n_818),
.B(n_851),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_894),
.B(n_854),
.Y(n_1027)
);

INVxp67_ASAP7_75t_L g1028 ( 
.A(n_922),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_L g1029 ( 
.A1(n_943),
.A2(n_803),
.B1(n_827),
.B2(n_933),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_869),
.B(n_943),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_855),
.B(n_925),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_891),
.A2(n_865),
.B(n_910),
.C(n_934),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_859),
.B(n_829),
.Y(n_1033)
);

NOR2x1_ASAP7_75t_L g1034 ( 
.A(n_812),
.B(n_794),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_821),
.A2(n_823),
.B(n_826),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_928),
.Y(n_1036)
);

O2A1O1Ixp5_ASAP7_75t_L g1037 ( 
.A1(n_788),
.A2(n_789),
.B(n_947),
.C(n_771),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_891),
.B(n_927),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_927),
.B(n_923),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_818),
.B(n_801),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_797),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_801),
.B(n_815),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_917),
.B(n_931),
.Y(n_1043)
);

NOR2x1_ASAP7_75t_R g1044 ( 
.A(n_793),
.B(n_814),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_928),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_815),
.B(n_851),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_860),
.B(n_825),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_SL g1048 ( 
.A1(n_904),
.A2(n_939),
.B1(n_772),
.B2(n_937),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_803),
.A2(n_827),
.B(n_850),
.C(n_860),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_900),
.B(n_908),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_807),
.A2(n_808),
.B(n_786),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_899),
.A2(n_903),
.B(n_895),
.C(n_795),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_839),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_845),
.A2(n_804),
.B(n_832),
.Y(n_1054)
);

BUFx2_ASAP7_75t_L g1055 ( 
.A(n_904),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_841),
.B(n_928),
.Y(n_1056)
);

OR2x6_ASAP7_75t_L g1057 ( 
.A(n_881),
.B(n_794),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_810),
.A2(n_813),
.B(n_783),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_834),
.A2(n_841),
.B1(n_940),
.B2(n_935),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_858),
.B(n_884),
.Y(n_1060)
);

NOR3xp33_ASAP7_75t_SL g1061 ( 
.A(n_912),
.B(n_903),
.C(n_938),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_932),
.B(n_920),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_853),
.A2(n_844),
.B(n_864),
.C(n_924),
.Y(n_1063)
);

AOI221xp5_ASAP7_75t_L g1064 ( 
.A1(n_873),
.A2(n_885),
.B1(n_883),
.B2(n_875),
.C(n_778),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_879),
.A2(n_837),
.B(n_833),
.C(n_831),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_828),
.A2(n_888),
.B(n_893),
.C(n_915),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_932),
.Y(n_1067)
);

AOI21x1_ASAP7_75t_L g1068 ( 
.A1(n_912),
.A2(n_870),
.B(n_896),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_781),
.B(n_863),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_887),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_856),
.B(n_862),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_929),
.A2(n_919),
.B1(n_901),
.B2(n_902),
.Y(n_1072)
);

NAND2x1p5_ASAP7_75t_L g1073 ( 
.A(n_911),
.B(n_898),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_892),
.B(n_611),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_777),
.A2(n_806),
.B1(n_889),
.B2(n_811),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_944),
.B(n_785),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_857),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_857),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_777),
.A2(n_785),
.B1(n_641),
.B2(n_607),
.Y(n_1079)
);

INVx6_ASAP7_75t_L g1080 ( 
.A(n_782),
.Y(n_1080)
);

INVx4_ASAP7_75t_L g1081 ( 
.A(n_822),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_944),
.B(n_785),
.Y(n_1082)
);

BUFx12f_ASAP7_75t_L g1083 ( 
.A(n_881),
.Y(n_1083)
);

OR2x6_ASAP7_75t_L g1084 ( 
.A(n_881),
.B(n_658),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_944),
.B(n_619),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_847),
.A2(n_680),
.B(n_643),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_955),
.A2(n_1086),
.B(n_1006),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1085),
.B(n_980),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1069),
.A2(n_1082),
.B(n_1076),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1082),
.A2(n_1051),
.B(n_1020),
.Y(n_1090)
);

OA21x2_ASAP7_75t_L g1091 ( 
.A1(n_972),
.A2(n_1037),
.B(n_1049),
.Y(n_1091)
);

AOI21x1_ASAP7_75t_L g1092 ( 
.A1(n_1009),
.A2(n_962),
.B(n_956),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1020),
.A2(n_1023),
.B(n_1031),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_974),
.Y(n_1094)
);

NOR2xp67_ASAP7_75t_L g1095 ( 
.A(n_960),
.B(n_963),
.Y(n_1095)
);

AO32x2_ASAP7_75t_L g1096 ( 
.A1(n_1079),
.A2(n_977),
.A3(n_970),
.B1(n_1001),
.B2(n_1059),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_1054),
.A2(n_966),
.B(n_1035),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1012),
.B(n_1015),
.Y(n_1098)
);

OR2x6_ASAP7_75t_L g1099 ( 
.A(n_1084),
.B(n_1080),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_1022),
.B(n_1075),
.Y(n_1100)
);

NAND2x1p5_ASAP7_75t_L g1101 ( 
.A(n_1034),
.B(n_986),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_965),
.B(n_1027),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1005),
.B(n_950),
.Y(n_1103)
);

BUFx12f_ASAP7_75t_L g1104 ( 
.A(n_993),
.Y(n_1104)
);

O2A1O1Ixp5_ASAP7_75t_L g1105 ( 
.A1(n_1032),
.A2(n_992),
.B(n_1004),
.C(n_1062),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_1028),
.B(n_1039),
.Y(n_1106)
);

AO32x2_ASAP7_75t_L g1107 ( 
.A1(n_1079),
.A2(n_977),
.A3(n_1001),
.B1(n_1059),
.B2(n_1021),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_1007),
.A2(n_978),
.B(n_1058),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_1030),
.A2(n_1043),
.B1(n_996),
.B2(n_999),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_1017),
.A2(n_959),
.B(n_961),
.C(n_1029),
.Y(n_1110)
);

AO31x2_ASAP7_75t_L g1111 ( 
.A1(n_969),
.A2(n_1065),
.A3(n_1063),
.B(n_1072),
.Y(n_1111)
);

BUFx12f_ASAP7_75t_L g1112 ( 
.A(n_993),
.Y(n_1112)
);

BUFx10_ASAP7_75t_L g1113 ( 
.A(n_1080),
.Y(n_1113)
);

INVx3_ASAP7_75t_L g1114 ( 
.A(n_1057),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_949),
.Y(n_1115)
);

NAND3x1_ASAP7_75t_L g1116 ( 
.A(n_1003),
.B(n_1033),
.C(n_998),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_1057),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_1057),
.B(n_985),
.Y(n_1118)
);

INVxp67_ASAP7_75t_SL g1119 ( 
.A(n_990),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1071),
.A2(n_1011),
.B(n_973),
.Y(n_1120)
);

AO31x2_ASAP7_75t_L g1121 ( 
.A1(n_1072),
.A2(n_1066),
.A3(n_1074),
.B(n_995),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_1000),
.B(n_971),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1052),
.A2(n_1064),
.B(n_1026),
.Y(n_1123)
);

AO32x2_ASAP7_75t_L g1124 ( 
.A1(n_1002),
.A2(n_981),
.A3(n_1081),
.B1(n_1025),
.B2(n_983),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_967),
.A2(n_1038),
.B(n_1014),
.Y(n_1125)
);

AO31x2_ASAP7_75t_L g1126 ( 
.A1(n_995),
.A2(n_997),
.A3(n_1050),
.B(n_1040),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1068),
.A2(n_1073),
.B(n_953),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1013),
.B(n_951),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_1055),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_1018),
.B(n_964),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_948),
.A2(n_1073),
.B(n_1047),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_948),
.A2(n_1046),
.B(n_975),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1060),
.A2(n_1042),
.B(n_984),
.Y(n_1133)
);

AO31x2_ASAP7_75t_L g1134 ( 
.A1(n_997),
.A2(n_1024),
.A3(n_1060),
.B(n_1041),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1070),
.A2(n_988),
.B(n_989),
.Y(n_1135)
);

CKINVDCx8_ASAP7_75t_R g1136 ( 
.A(n_979),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_987),
.A2(n_976),
.B(n_954),
.C(n_1077),
.Y(n_1137)
);

AO31x2_ASAP7_75t_L g1138 ( 
.A1(n_968),
.A2(n_994),
.A3(n_1053),
.B(n_1067),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1078),
.B(n_1048),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_988),
.A2(n_1056),
.B(n_991),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_1010),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_952),
.Y(n_1142)
);

OAI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_957),
.A2(n_1019),
.B(n_982),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_957),
.B(n_1019),
.Y(n_1144)
);

AO32x2_ASAP7_75t_L g1145 ( 
.A1(n_981),
.A2(n_983),
.A3(n_1008),
.B1(n_1081),
.B2(n_1025),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1061),
.B(n_1084),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1010),
.A2(n_1016),
.B(n_1036),
.Y(n_1147)
);

A2O1A1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_1016),
.A2(n_1036),
.B(n_1045),
.C(n_1044),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1084),
.A2(n_1083),
.B(n_1036),
.C(n_1045),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1016),
.A2(n_955),
.B(n_847),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1045),
.A2(n_955),
.B(n_847),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_993),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_960),
.B(n_316),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_960),
.B(n_316),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1007),
.A2(n_966),
.B(n_1023),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_SL g1156 ( 
.A1(n_1079),
.A2(n_847),
.B(n_785),
.Y(n_1156)
);

AOI21x1_ASAP7_75t_L g1157 ( 
.A1(n_955),
.A2(n_1009),
.B(n_962),
.Y(n_1157)
);

AOI21x1_ASAP7_75t_L g1158 ( 
.A1(n_955),
.A2(n_1009),
.B(n_962),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_974),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1007),
.A2(n_966),
.B(n_1023),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_955),
.A2(n_847),
.B(n_1086),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_1057),
.B(n_985),
.Y(n_1162)
);

AO31x2_ASAP7_75t_L g1163 ( 
.A1(n_1049),
.A2(n_811),
.A3(n_969),
.B(n_1065),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_1057),
.B(n_985),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1007),
.A2(n_966),
.B(n_1023),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1007),
.A2(n_966),
.B(n_1023),
.Y(n_1166)
);

INVx5_ASAP7_75t_L g1167 ( 
.A(n_1010),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_955),
.A2(n_847),
.B(n_1086),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1012),
.B(n_880),
.Y(n_1169)
);

INVxp67_ASAP7_75t_L g1170 ( 
.A(n_974),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_958),
.Y(n_1171)
);

OAI21xp33_ASAP7_75t_L g1172 ( 
.A1(n_960),
.A2(n_700),
.B(n_784),
.Y(n_1172)
);

AO31x2_ASAP7_75t_L g1173 ( 
.A1(n_1049),
.A2(n_811),
.A3(n_969),
.B(n_1065),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_960),
.B(n_316),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_958),
.Y(n_1175)
);

A2O1A1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_960),
.A2(n_806),
.B(n_777),
.C(n_724),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_960),
.A2(n_806),
.B(n_777),
.C(n_724),
.Y(n_1177)
);

AO22x2_ASAP7_75t_L g1178 ( 
.A1(n_960),
.A2(n_777),
.B1(n_977),
.B2(n_1079),
.Y(n_1178)
);

AO31x2_ASAP7_75t_L g1179 ( 
.A1(n_1049),
.A2(n_811),
.A3(n_969),
.B(n_1065),
.Y(n_1179)
);

INVx2_ASAP7_75t_SL g1180 ( 
.A(n_993),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_958),
.Y(n_1181)
);

AOI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_960),
.A2(n_777),
.B1(n_316),
.B2(n_330),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_960),
.A2(n_777),
.B1(n_1082),
.B2(n_1076),
.Y(n_1183)
);

AO31x2_ASAP7_75t_L g1184 ( 
.A1(n_1049),
.A2(n_811),
.A3(n_969),
.B(n_1065),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_960),
.A2(n_806),
.B(n_777),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1085),
.B(n_980),
.Y(n_1186)
);

AO31x2_ASAP7_75t_L g1187 ( 
.A1(n_1049),
.A2(n_811),
.A3(n_969),
.B(n_1065),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1057),
.B(n_985),
.Y(n_1188)
);

AO31x2_ASAP7_75t_L g1189 ( 
.A1(n_1049),
.A2(n_811),
.A3(n_969),
.B(n_1065),
.Y(n_1189)
);

NOR2xp67_ASAP7_75t_L g1190 ( 
.A(n_960),
.B(n_963),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1057),
.B(n_985),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_958),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_955),
.A2(n_847),
.B(n_1086),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_960),
.A2(n_806),
.B(n_777),
.C(n_724),
.Y(n_1194)
);

BUFx10_ASAP7_75t_L g1195 ( 
.A(n_1080),
.Y(n_1195)
);

AO32x2_ASAP7_75t_L g1196 ( 
.A1(n_1079),
.A2(n_977),
.A3(n_970),
.B1(n_1001),
.B2(n_1059),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_955),
.A2(n_847),
.B(n_1086),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_960),
.B(n_777),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_958),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1085),
.B(n_980),
.Y(n_1200)
);

CKINVDCx6p67_ASAP7_75t_R g1201 ( 
.A(n_952),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1004),
.A2(n_806),
.B(n_777),
.C(n_395),
.Y(n_1202)
);

OAI21xp5_ASAP7_75t_SL g1203 ( 
.A1(n_960),
.A2(n_497),
.B(n_515),
.Y(n_1203)
);

O2A1O1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_1004),
.A2(n_806),
.B(n_777),
.C(n_395),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1007),
.A2(n_966),
.B(n_1023),
.Y(n_1205)
);

NOR2xp67_ASAP7_75t_L g1206 ( 
.A(n_960),
.B(n_963),
.Y(n_1206)
);

AOI211x1_ASAP7_75t_L g1207 ( 
.A1(n_960),
.A2(n_806),
.B(n_582),
.C(n_777),
.Y(n_1207)
);

A2O1A1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_960),
.A2(n_806),
.B(n_777),
.C(n_724),
.Y(n_1208)
);

A2O1A1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_960),
.A2(n_806),
.B(n_777),
.C(n_724),
.Y(n_1209)
);

AO31x2_ASAP7_75t_L g1210 ( 
.A1(n_1049),
.A2(n_811),
.A3(n_969),
.B(n_1065),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_1057),
.B(n_985),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_960),
.A2(n_806),
.B(n_777),
.Y(n_1212)
);

INVx8_ASAP7_75t_L g1213 ( 
.A(n_1057),
.Y(n_1213)
);

AOI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_960),
.A2(n_777),
.B1(n_316),
.B2(n_330),
.Y(n_1214)
);

INVx5_ASAP7_75t_L g1215 ( 
.A(n_1010),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_974),
.Y(n_1216)
);

OR2x6_ASAP7_75t_L g1217 ( 
.A(n_1084),
.B(n_1080),
.Y(n_1217)
);

AOI21x1_ASAP7_75t_SL g1218 ( 
.A1(n_992),
.A2(n_997),
.B(n_995),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1153),
.A2(n_1154),
.B1(n_1174),
.B2(n_1203),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_SL g1220 ( 
.A1(n_1178),
.A2(n_1212),
.B1(n_1185),
.B2(n_1139),
.Y(n_1220)
);

INVx5_ASAP7_75t_L g1221 ( 
.A(n_1167),
.Y(n_1221)
);

INVxp67_ASAP7_75t_L g1222 ( 
.A(n_1122),
.Y(n_1222)
);

OAI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1182),
.A2(n_1214),
.B1(n_1102),
.B2(n_1088),
.Y(n_1223)
);

AOI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1172),
.A2(n_1109),
.B1(n_1116),
.B2(n_1106),
.Y(n_1224)
);

CKINVDCx20_ASAP7_75t_R g1225 ( 
.A(n_1136),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1159),
.Y(n_1226)
);

CKINVDCx11_ASAP7_75t_R g1227 ( 
.A(n_1195),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1175),
.Y(n_1228)
);

CKINVDCx11_ASAP7_75t_R g1229 ( 
.A(n_1195),
.Y(n_1229)
);

INVx2_ASAP7_75t_SL g1230 ( 
.A(n_1113),
.Y(n_1230)
);

INVxp67_ASAP7_75t_SL g1231 ( 
.A(n_1115),
.Y(n_1231)
);

BUFx12f_ASAP7_75t_L g1232 ( 
.A(n_1142),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1186),
.A2(n_1200),
.B1(n_1110),
.B2(n_1103),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_SL g1234 ( 
.A1(n_1178),
.A2(n_1123),
.B1(n_1183),
.B2(n_1162),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1176),
.A2(n_1209),
.B1(n_1208),
.B2(n_1194),
.Y(n_1235)
);

OAI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1095),
.A2(n_1206),
.B1(n_1190),
.B2(n_1217),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_1129),
.Y(n_1237)
);

INVx6_ASAP7_75t_L g1238 ( 
.A(n_1167),
.Y(n_1238)
);

OAI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1099),
.A2(n_1217),
.B1(n_1100),
.B2(n_1125),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1094),
.Y(n_1240)
);

OAI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1099),
.A2(n_1198),
.B1(n_1114),
.B2(n_1117),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1098),
.A2(n_1169),
.B1(n_1130),
.B2(n_1146),
.Y(n_1242)
);

BUFx10_ASAP7_75t_L g1243 ( 
.A(n_1142),
.Y(n_1243)
);

BUFx4f_ASAP7_75t_SL g1244 ( 
.A(n_1104),
.Y(n_1244)
);

INVx6_ASAP7_75t_L g1245 ( 
.A(n_1215),
.Y(n_1245)
);

BUFx10_ASAP7_75t_L g1246 ( 
.A(n_1180),
.Y(n_1246)
);

CKINVDCx11_ASAP7_75t_R g1247 ( 
.A(n_1201),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1118),
.A2(n_1164),
.B1(n_1211),
.B2(n_1188),
.Y(n_1248)
);

CKINVDCx11_ASAP7_75t_R g1249 ( 
.A(n_1112),
.Y(n_1249)
);

CKINVDCx11_ASAP7_75t_R g1250 ( 
.A(n_1216),
.Y(n_1250)
);

BUFx12f_ASAP7_75t_L g1251 ( 
.A(n_1101),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_SL g1252 ( 
.A(n_1202),
.B(n_1204),
.Y(n_1252)
);

INVx6_ASAP7_75t_L g1253 ( 
.A(n_1215),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1118),
.A2(n_1211),
.B1(n_1162),
.B2(n_1188),
.Y(n_1254)
);

OAI22xp33_ASAP7_75t_R g1255 ( 
.A1(n_1119),
.A2(n_1181),
.B1(n_1192),
.B2(n_1199),
.Y(n_1255)
);

INVx6_ASAP7_75t_L g1256 ( 
.A(n_1215),
.Y(n_1256)
);

BUFx8_ASAP7_75t_SL g1257 ( 
.A(n_1152),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1177),
.A2(n_1191),
.B1(n_1164),
.B2(n_1089),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1120),
.B(n_1207),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1170),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_1141),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_1213),
.Y(n_1262)
);

BUFx8_ASAP7_75t_L g1263 ( 
.A(n_1145),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1128),
.A2(n_1137),
.B1(n_1090),
.B2(n_1156),
.Y(n_1264)
);

INVx1_ASAP7_75t_SL g1265 ( 
.A(n_1144),
.Y(n_1265)
);

CKINVDCx11_ASAP7_75t_R g1266 ( 
.A(n_1213),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1093),
.A2(n_1135),
.B1(n_1148),
.B2(n_1149),
.Y(n_1267)
);

NAND2x1p5_ASAP7_75t_L g1268 ( 
.A(n_1140),
.B(n_1127),
.Y(n_1268)
);

INVx1_ASAP7_75t_SL g1269 ( 
.A(n_1147),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_SL g1270 ( 
.A1(n_1107),
.A2(n_1091),
.B1(n_1196),
.B2(n_1096),
.Y(n_1270)
);

OR2x2_ASAP7_75t_L g1271 ( 
.A(n_1138),
.B(n_1126),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1133),
.A2(n_1132),
.B1(n_1131),
.B2(n_1143),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1138),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1150),
.A2(n_1151),
.B1(n_1161),
.B2(n_1168),
.Y(n_1274)
);

CKINVDCx16_ASAP7_75t_R g1275 ( 
.A(n_1218),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1134),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1126),
.B(n_1210),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_SL g1278 ( 
.A1(n_1107),
.A2(n_1196),
.B1(n_1096),
.B2(n_1163),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_SL g1279 ( 
.A1(n_1107),
.A2(n_1196),
.B1(n_1096),
.B2(n_1163),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1193),
.A2(n_1197),
.B1(n_1087),
.B2(n_1097),
.Y(n_1280)
);

CKINVDCx16_ASAP7_75t_R g1281 ( 
.A(n_1145),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1163),
.A2(n_1210),
.B1(n_1189),
.B2(n_1187),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1155),
.A2(n_1166),
.B1(n_1160),
.B2(n_1165),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_SL g1284 ( 
.A1(n_1173),
.A2(n_1187),
.B1(n_1184),
.B2(n_1179),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1092),
.B(n_1158),
.Y(n_1285)
);

CKINVDCx11_ASAP7_75t_R g1286 ( 
.A(n_1105),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1173),
.A2(n_1210),
.B1(n_1184),
.B2(n_1187),
.Y(n_1287)
);

INVx6_ASAP7_75t_L g1288 ( 
.A(n_1145),
.Y(n_1288)
);

NAND2x1p5_ASAP7_75t_L g1289 ( 
.A(n_1157),
.B(n_1108),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1205),
.A2(n_1189),
.B1(n_1184),
.B2(n_1179),
.Y(n_1290)
);

INVx6_ASAP7_75t_L g1291 ( 
.A(n_1124),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1179),
.A2(n_1189),
.B1(n_1111),
.B2(n_1121),
.Y(n_1292)
);

CKINVDCx6p67_ASAP7_75t_R g1293 ( 
.A(n_1124),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1111),
.A2(n_806),
.B1(n_960),
.B2(n_777),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1172),
.A2(n_806),
.B1(n_960),
.B2(n_777),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1172),
.A2(n_806),
.B1(n_960),
.B2(n_777),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1171),
.Y(n_1297)
);

INVxp67_ASAP7_75t_SL g1298 ( 
.A(n_1089),
.Y(n_1298)
);

BUFx12f_ASAP7_75t_L g1299 ( 
.A(n_1195),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1153),
.A2(n_398),
.B1(n_404),
.B2(n_389),
.Y(n_1300)
);

INVx6_ASAP7_75t_L g1301 ( 
.A(n_1195),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1172),
.A2(n_806),
.B1(n_960),
.B2(n_777),
.Y(n_1302)
);

OR2x2_ASAP7_75t_L g1303 ( 
.A(n_1102),
.B(n_1098),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_1094),
.Y(n_1304)
);

CKINVDCx11_ASAP7_75t_R g1305 ( 
.A(n_1136),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1172),
.A2(n_806),
.B1(n_960),
.B2(n_777),
.Y(n_1306)
);

CKINVDCx14_ASAP7_75t_R g1307 ( 
.A(n_1195),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1159),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_SL g1309 ( 
.A1(n_1153),
.A2(n_777),
.B1(n_960),
.B2(n_329),
.Y(n_1309)
);

INVx3_ASAP7_75t_SL g1310 ( 
.A(n_1201),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1172),
.A2(n_806),
.B1(n_960),
.B2(n_777),
.Y(n_1311)
);

CKINVDCx20_ASAP7_75t_R g1312 ( 
.A(n_1136),
.Y(n_1312)
);

INVx5_ASAP7_75t_L g1313 ( 
.A(n_1167),
.Y(n_1313)
);

CKINVDCx11_ASAP7_75t_R g1314 ( 
.A(n_1136),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1102),
.A2(n_777),
.B1(n_1109),
.B2(n_1088),
.Y(n_1315)
);

CKINVDCx11_ASAP7_75t_R g1316 ( 
.A(n_1136),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1171),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_1136),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1102),
.A2(n_777),
.B1(n_1109),
.B2(n_1088),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1195),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1172),
.A2(n_806),
.B1(n_960),
.B2(n_777),
.Y(n_1321)
);

CKINVDCx11_ASAP7_75t_R g1322 ( 
.A(n_1136),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1172),
.A2(n_806),
.B1(n_960),
.B2(n_777),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1102),
.A2(n_777),
.B1(n_1109),
.B2(n_1088),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1102),
.A2(n_777),
.B1(n_1109),
.B2(n_1088),
.Y(n_1325)
);

AOI22x1_ASAP7_75t_L g1326 ( 
.A1(n_1178),
.A2(n_1125),
.B1(n_1212),
.B2(n_1185),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1172),
.A2(n_806),
.B1(n_960),
.B2(n_777),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1273),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1276),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1263),
.Y(n_1330)
);

INVx2_ASAP7_75t_SL g1331 ( 
.A(n_1288),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1289),
.A2(n_1283),
.B(n_1268),
.Y(n_1332)
);

AOI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1252),
.A2(n_1264),
.B(n_1267),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1271),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1278),
.A2(n_1279),
.B1(n_1270),
.B2(n_1309),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1278),
.B(n_1279),
.Y(n_1336)
);

AO31x2_ASAP7_75t_L g1337 ( 
.A1(n_1282),
.A2(n_1287),
.A3(n_1264),
.B(n_1285),
.Y(n_1337)
);

INVx2_ASAP7_75t_SL g1338 ( 
.A(n_1238),
.Y(n_1338)
);

BUFx4f_ASAP7_75t_SL g1339 ( 
.A(n_1232),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_1305),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1277),
.Y(n_1341)
);

AO21x2_ASAP7_75t_L g1342 ( 
.A1(n_1259),
.A2(n_1298),
.B(n_1282),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1288),
.Y(n_1343)
);

AO21x2_ASAP7_75t_L g1344 ( 
.A1(n_1259),
.A2(n_1298),
.B(n_1287),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1263),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1288),
.Y(n_1346)
);

OR2x6_ASAP7_75t_L g1347 ( 
.A(n_1258),
.B(n_1291),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1222),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1326),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1284),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1284),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_1293),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1222),
.Y(n_1353)
);

INVx2_ASAP7_75t_SL g1354 ( 
.A(n_1221),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1274),
.A2(n_1280),
.B(n_1272),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1292),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1235),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1235),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1270),
.Y(n_1359)
);

AO21x2_ASAP7_75t_L g1360 ( 
.A1(n_1267),
.A2(n_1258),
.B(n_1239),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1290),
.Y(n_1361)
);

AO21x1_ASAP7_75t_SL g1362 ( 
.A1(n_1224),
.A2(n_1294),
.B(n_1327),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1233),
.B(n_1220),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1219),
.B(n_1303),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1228),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1233),
.A2(n_1325),
.B(n_1324),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1281),
.B(n_1220),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1234),
.B(n_1315),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1297),
.Y(n_1369)
);

AO21x2_ASAP7_75t_L g1370 ( 
.A1(n_1315),
.A2(n_1325),
.B(n_1324),
.Y(n_1370)
);

AO21x1_ASAP7_75t_SL g1371 ( 
.A1(n_1295),
.A2(n_1296),
.B(n_1321),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1300),
.B(n_1223),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1234),
.B(n_1317),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_1286),
.Y(n_1374)
);

INVx2_ASAP7_75t_SL g1375 ( 
.A(n_1238),
.Y(n_1375)
);

AO21x2_ASAP7_75t_L g1376 ( 
.A1(n_1319),
.A2(n_1241),
.B(n_1236),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1231),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1265),
.Y(n_1378)
);

OA21x2_ASAP7_75t_L g1379 ( 
.A1(n_1302),
.A2(n_1306),
.B(n_1311),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1269),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1255),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_1240),
.Y(n_1382)
);

AO21x2_ASAP7_75t_L g1383 ( 
.A1(n_1319),
.A2(n_1275),
.B(n_1323),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1221),
.A2(n_1313),
.B(n_1309),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1242),
.B(n_1304),
.Y(n_1385)
);

BUFx2_ASAP7_75t_L g1386 ( 
.A(n_1261),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1248),
.B(n_1254),
.Y(n_1387)
);

OA21x2_ASAP7_75t_L g1388 ( 
.A1(n_1260),
.A2(n_1226),
.B(n_1308),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1245),
.A2(n_1253),
.B(n_1256),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1237),
.B(n_1262),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1246),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1251),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1301),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1301),
.Y(n_1394)
);

O2A1O1Ixp33_ASAP7_75t_SL g1395 ( 
.A1(n_1363),
.A2(n_1230),
.B(n_1225),
.C(n_1318),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1377),
.B(n_1320),
.Y(n_1396)
);

A2O1A1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1366),
.A2(n_1307),
.B(n_1312),
.C(n_1266),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1330),
.B(n_1250),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1330),
.B(n_1243),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_1386),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1345),
.B(n_1243),
.Y(n_1401)
);

AO32x2_ASAP7_75t_L g1402 ( 
.A1(n_1335),
.A2(n_1257),
.A3(n_1301),
.B1(n_1229),
.B2(n_1227),
.Y(n_1402)
);

O2A1O1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1372),
.A2(n_1366),
.B(n_1363),
.C(n_1368),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1373),
.B(n_1322),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1367),
.B(n_1348),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1367),
.B(n_1316),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1353),
.B(n_1314),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1388),
.B(n_1310),
.Y(n_1408)
);

OA21x2_ASAP7_75t_L g1409 ( 
.A1(n_1355),
.A2(n_1244),
.B(n_1299),
.Y(n_1409)
);

AOI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1384),
.A2(n_1249),
.B(n_1247),
.Y(n_1410)
);

AOI221xp5_ASAP7_75t_L g1411 ( 
.A1(n_1335),
.A2(n_1368),
.B1(n_1364),
.B2(n_1357),
.C(n_1358),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1343),
.B(n_1346),
.Y(n_1412)
);

BUFx4f_ASAP7_75t_SL g1413 ( 
.A(n_1390),
.Y(n_1413)
);

INVx1_ASAP7_75t_SL g1414 ( 
.A(n_1378),
.Y(n_1414)
);

BUFx10_ASAP7_75t_L g1415 ( 
.A(n_1340),
.Y(n_1415)
);

A2O1A1Ixp33_ASAP7_75t_L g1416 ( 
.A1(n_1384),
.A2(n_1358),
.B(n_1357),
.C(n_1349),
.Y(n_1416)
);

AO21x2_ASAP7_75t_L g1417 ( 
.A1(n_1333),
.A2(n_1370),
.B(n_1332),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1339),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1374),
.A2(n_1381),
.B1(n_1385),
.B2(n_1387),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1371),
.A2(n_1370),
.B1(n_1362),
.B2(n_1379),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1333),
.A2(n_1379),
.B(n_1349),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1382),
.B(n_1386),
.Y(n_1422)
);

AND2x2_ASAP7_75t_SL g1423 ( 
.A(n_1374),
.B(n_1336),
.Y(n_1423)
);

OAI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1379),
.A2(n_1349),
.B(n_1355),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1379),
.A2(n_1355),
.B(n_1380),
.Y(n_1425)
);

AO32x2_ASAP7_75t_L g1426 ( 
.A1(n_1331),
.A2(n_1354),
.A3(n_1338),
.B1(n_1375),
.B2(n_1359),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1379),
.B(n_1383),
.Y(n_1427)
);

OAI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1380),
.A2(n_1387),
.B(n_1385),
.Y(n_1428)
);

AOI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1370),
.A2(n_1383),
.B1(n_1360),
.B2(n_1376),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_SL g1430 ( 
.A1(n_1370),
.A2(n_1374),
.B1(n_1360),
.B2(n_1383),
.Y(n_1430)
);

CKINVDCx20_ASAP7_75t_R g1431 ( 
.A(n_1374),
.Y(n_1431)
);

AO32x2_ASAP7_75t_L g1432 ( 
.A1(n_1331),
.A2(n_1354),
.A3(n_1338),
.B1(n_1375),
.B2(n_1359),
.Y(n_1432)
);

A2O1A1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1374),
.A2(n_1360),
.B(n_1350),
.C(n_1351),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1392),
.Y(n_1434)
);

OR2x6_ASAP7_75t_L g1435 ( 
.A(n_1347),
.B(n_1389),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1347),
.A2(n_1392),
.B1(n_1390),
.B2(n_1394),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1329),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1360),
.A2(n_1342),
.B(n_1344),
.Y(n_1438)
);

AO32x2_ASAP7_75t_L g1439 ( 
.A1(n_1354),
.A2(n_1350),
.A3(n_1351),
.B1(n_1334),
.B2(n_1337),
.Y(n_1439)
);

A2O1A1Ixp33_ASAP7_75t_L g1440 ( 
.A1(n_1362),
.A2(n_1371),
.B(n_1352),
.C(n_1383),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1439),
.B(n_1337),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1437),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1439),
.B(n_1337),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1439),
.B(n_1337),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1439),
.B(n_1337),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1435),
.B(n_1337),
.Y(n_1446)
);

OAI221xp5_ASAP7_75t_SL g1447 ( 
.A1(n_1403),
.A2(n_1347),
.B1(n_1352),
.B2(n_1356),
.C(n_1376),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1435),
.B(n_1344),
.Y(n_1448)
);

BUFx2_ASAP7_75t_L g1449 ( 
.A(n_1426),
.Y(n_1449)
);

INVx1_ASAP7_75t_SL g1450 ( 
.A(n_1408),
.Y(n_1450)
);

INVx1_ASAP7_75t_SL g1451 ( 
.A(n_1414),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1427),
.B(n_1341),
.Y(n_1452)
);

INVxp67_ASAP7_75t_SL g1453 ( 
.A(n_1421),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1411),
.A2(n_1376),
.B1(n_1347),
.B2(n_1361),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1426),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1432),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1417),
.B(n_1344),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1420),
.A2(n_1376),
.B1(n_1361),
.B2(n_1342),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1417),
.B(n_1342),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1432),
.Y(n_1460)
);

INVxp67_ASAP7_75t_SL g1461 ( 
.A(n_1425),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1433),
.A2(n_1391),
.B1(n_1394),
.B2(n_1393),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1446),
.B(n_1424),
.Y(n_1463)
);

INVx5_ASAP7_75t_L g1464 ( 
.A(n_1457),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1446),
.B(n_1430),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1462),
.B(n_1433),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1446),
.B(n_1430),
.Y(n_1467)
);

OAI221xp5_ASAP7_75t_L g1468 ( 
.A1(n_1447),
.A2(n_1420),
.B1(n_1397),
.B2(n_1440),
.C(n_1429),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1449),
.B(n_1412),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1452),
.B(n_1342),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1447),
.A2(n_1438),
.B(n_1440),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1451),
.B(n_1413),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1455),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1455),
.Y(n_1474)
);

OAI33xp33_ASAP7_75t_L g1475 ( 
.A1(n_1462),
.A2(n_1419),
.A3(n_1402),
.B1(n_1396),
.B2(n_1369),
.B3(n_1365),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1452),
.B(n_1405),
.Y(n_1476)
);

OAI211xp5_ASAP7_75t_L g1477 ( 
.A1(n_1454),
.A2(n_1397),
.B(n_1395),
.C(n_1428),
.Y(n_1477)
);

AOI33xp33_ASAP7_75t_L g1478 ( 
.A1(n_1454),
.A2(n_1395),
.A3(n_1406),
.B1(n_1404),
.B2(n_1402),
.B3(n_1422),
.Y(n_1478)
);

AOI33xp33_ASAP7_75t_L g1479 ( 
.A1(n_1458),
.A2(n_1441),
.A3(n_1443),
.B1(n_1444),
.B2(n_1445),
.B3(n_1457),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1442),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1453),
.A2(n_1416),
.B(n_1409),
.Y(n_1481)
);

AO21x2_ASAP7_75t_L g1482 ( 
.A1(n_1459),
.A2(n_1328),
.B(n_1416),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1442),
.Y(n_1483)
);

AOI33xp33_ASAP7_75t_L g1484 ( 
.A1(n_1458),
.A2(n_1445),
.A3(n_1444),
.B1(n_1443),
.B2(n_1441),
.B3(n_1459),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1473),
.B(n_1460),
.Y(n_1485)
);

NOR3xp33_ASAP7_75t_L g1486 ( 
.A(n_1477),
.B(n_1453),
.C(n_1461),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1480),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1480),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1473),
.B(n_1456),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1480),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1464),
.B(n_1448),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1483),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1469),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1473),
.B(n_1474),
.Y(n_1494)
);

AND2x4_ASAP7_75t_SL g1495 ( 
.A(n_1472),
.B(n_1431),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1464),
.B(n_1448),
.Y(n_1496)
);

BUFx3_ASAP7_75t_L g1497 ( 
.A(n_1472),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1473),
.B(n_1456),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1464),
.B(n_1461),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1483),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1483),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1464),
.B(n_1441),
.Y(n_1502)
);

INVxp67_ASAP7_75t_L g1503 ( 
.A(n_1466),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1464),
.B(n_1443),
.Y(n_1504)
);

INVx2_ASAP7_75t_SL g1505 ( 
.A(n_1464),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1464),
.B(n_1444),
.Y(n_1506)
);

CKINVDCx14_ASAP7_75t_R g1507 ( 
.A(n_1465),
.Y(n_1507)
);

OAI31xp33_ASAP7_75t_L g1508 ( 
.A1(n_1477),
.A2(n_1402),
.A3(n_1451),
.B(n_1436),
.Y(n_1508)
);

BUFx2_ASAP7_75t_L g1509 ( 
.A(n_1469),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1474),
.Y(n_1510)
);

INVx2_ASAP7_75t_SL g1511 ( 
.A(n_1464),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1476),
.B(n_1484),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1503),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1494),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1507),
.B(n_1509),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1509),
.B(n_1465),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1492),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1512),
.B(n_1503),
.Y(n_1518)
);

OR2x6_ASAP7_75t_L g1519 ( 
.A(n_1505),
.B(n_1481),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1491),
.B(n_1465),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1492),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1491),
.B(n_1467),
.Y(n_1522)
);

INVx1_ASAP7_75t_SL g1523 ( 
.A(n_1497),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1512),
.B(n_1479),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1487),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1493),
.B(n_1470),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1491),
.B(n_1467),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1486),
.B(n_1479),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1494),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1487),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1488),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1496),
.B(n_1467),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1496),
.B(n_1463),
.Y(n_1533)
);

NOR2x1_ASAP7_75t_L g1534 ( 
.A(n_1497),
.B(n_1466),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1488),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1496),
.B(n_1463),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1497),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1494),
.Y(n_1538)
);

NOR2xp67_ASAP7_75t_L g1539 ( 
.A(n_1505),
.B(n_1481),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1489),
.B(n_1470),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1490),
.Y(n_1541)
);

INVxp67_ASAP7_75t_SL g1542 ( 
.A(n_1486),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1485),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1489),
.B(n_1476),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1490),
.Y(n_1545)
);

INVxp33_ASAP7_75t_L g1546 ( 
.A(n_1508),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1500),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1508),
.B(n_1478),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1500),
.Y(n_1549)
);

INVx2_ASAP7_75t_SL g1550 ( 
.A(n_1495),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1501),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1501),
.Y(n_1552)
);

AND2x2_ASAP7_75t_SL g1553 ( 
.A(n_1495),
.B(n_1478),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1510),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1513),
.B(n_1489),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1515),
.B(n_1502),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1525),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1525),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1515),
.B(n_1502),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1516),
.B(n_1504),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1530),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1516),
.B(n_1504),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1523),
.Y(n_1563)
);

AND2x4_ASAP7_75t_SL g1564 ( 
.A(n_1537),
.B(n_1431),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1518),
.B(n_1463),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1543),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1518),
.B(n_1484),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1528),
.B(n_1498),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1528),
.B(n_1498),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1530),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1531),
.Y(n_1571)
);

NAND2x1p5_ASAP7_75t_L g1572 ( 
.A(n_1534),
.B(n_1523),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1520),
.B(n_1504),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1520),
.B(n_1506),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1543),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1542),
.B(n_1534),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1548),
.B(n_1495),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1531),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1524),
.B(n_1400),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1524),
.B(n_1450),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1550),
.Y(n_1581)
);

NAND2xp67_ASAP7_75t_L g1582 ( 
.A(n_1546),
.B(n_1398),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1543),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1522),
.B(n_1506),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1535),
.Y(n_1585)
);

NAND2x2_ASAP7_75t_L g1586 ( 
.A(n_1550),
.B(n_1410),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1535),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1522),
.B(n_1506),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1544),
.B(n_1498),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1553),
.B(n_1450),
.Y(n_1590)
);

AOI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1576),
.A2(n_1553),
.B(n_1519),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1572),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1567),
.B(n_1563),
.Y(n_1593)
);

OAI21xp33_ASAP7_75t_L g1594 ( 
.A1(n_1582),
.A2(n_1553),
.B(n_1471),
.Y(n_1594)
);

OAI21xp5_ASAP7_75t_SL g1595 ( 
.A1(n_1572),
.A2(n_1471),
.B(n_1468),
.Y(n_1595)
);

INVx2_ASAP7_75t_SL g1596 ( 
.A(n_1564),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1557),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1557),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1558),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1580),
.B(n_1544),
.Y(n_1600)
);

AOI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1564),
.A2(n_1468),
.B1(n_1475),
.B2(n_1482),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1558),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_L g1603 ( 
.A(n_1582),
.B(n_1418),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1561),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1556),
.B(n_1527),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1579),
.B(n_1526),
.Y(n_1606)
);

AOI21xp33_ASAP7_75t_L g1607 ( 
.A1(n_1572),
.A2(n_1519),
.B(n_1539),
.Y(n_1607)
);

O2A1O1Ixp5_ASAP7_75t_L g1608 ( 
.A1(n_1590),
.A2(n_1577),
.B(n_1565),
.C(n_1475),
.Y(n_1608)
);

OAI221xp5_ASAP7_75t_L g1609 ( 
.A1(n_1586),
.A2(n_1539),
.B1(n_1519),
.B2(n_1505),
.C(n_1511),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1581),
.B(n_1418),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1568),
.B(n_1526),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1556),
.Y(n_1612)
);

AOI221xp5_ASAP7_75t_L g1613 ( 
.A1(n_1581),
.A2(n_1532),
.B1(n_1527),
.B2(n_1517),
.C(n_1521),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1559),
.B(n_1560),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1561),
.Y(n_1615)
);

NOR3xp33_ASAP7_75t_L g1616 ( 
.A(n_1595),
.B(n_1594),
.C(n_1593),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1596),
.B(n_1559),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1593),
.B(n_1560),
.Y(n_1618)
);

AOI211xp5_ASAP7_75t_SL g1619 ( 
.A1(n_1591),
.A2(n_1568),
.B(n_1569),
.C(n_1555),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1610),
.B(n_1562),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1597),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1601),
.B(n_1555),
.Y(n_1622)
);

OAI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1608),
.A2(n_1569),
.B(n_1519),
.Y(n_1623)
);

AOI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1603),
.A2(n_1586),
.B1(n_1562),
.B2(n_1532),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1605),
.B(n_1573),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1613),
.B(n_1573),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1612),
.B(n_1574),
.Y(n_1627)
);

INVx3_ASAP7_75t_L g1628 ( 
.A(n_1592),
.Y(n_1628)
);

OAI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1592),
.A2(n_1519),
.B1(n_1588),
.B2(n_1584),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1614),
.B(n_1574),
.Y(n_1630)
);

NOR2x1_ASAP7_75t_L g1631 ( 
.A(n_1598),
.B(n_1570),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1599),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1602),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1611),
.Y(n_1634)
);

AOI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1616),
.A2(n_1609),
.B1(n_1606),
.B2(n_1600),
.Y(n_1635)
);

OAI21xp33_ASAP7_75t_L g1636 ( 
.A1(n_1626),
.A2(n_1607),
.B(n_1604),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1631),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1634),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1634),
.Y(n_1639)
);

OAI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1619),
.A2(n_1607),
.B(n_1615),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1628),
.Y(n_1641)
);

OAI221xp5_ASAP7_75t_L g1642 ( 
.A1(n_1616),
.A2(n_1623),
.B1(n_1622),
.B2(n_1624),
.C(n_1617),
.Y(n_1642)
);

INVxp33_ASAP7_75t_L g1643 ( 
.A(n_1620),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1628),
.Y(n_1644)
);

AO21x1_ASAP7_75t_L g1645 ( 
.A1(n_1622),
.A2(n_1571),
.B(n_1570),
.Y(n_1645)
);

INVxp67_ASAP7_75t_SL g1646 ( 
.A(n_1645),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1641),
.B(n_1618),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1643),
.B(n_1625),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1644),
.B(n_1629),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1638),
.B(n_1630),
.Y(n_1650)
);

NOR3xp33_ASAP7_75t_L g1651 ( 
.A(n_1642),
.B(n_1632),
.C(n_1621),
.Y(n_1651)
);

OAI21xp5_ASAP7_75t_SL g1652 ( 
.A1(n_1640),
.A2(n_1627),
.B(n_1633),
.Y(n_1652)
);

O2A1O1Ixp33_ASAP7_75t_L g1653 ( 
.A1(n_1640),
.A2(n_1637),
.B(n_1636),
.C(n_1639),
.Y(n_1653)
);

OAI21xp33_ASAP7_75t_L g1654 ( 
.A1(n_1635),
.A2(n_1588),
.B(n_1584),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1641),
.B(n_1585),
.Y(n_1655)
);

AOI221xp5_ASAP7_75t_L g1656 ( 
.A1(n_1653),
.A2(n_1566),
.B1(n_1575),
.B2(n_1583),
.C(n_1578),
.Y(n_1656)
);

OAI211xp5_ASAP7_75t_SL g1657 ( 
.A1(n_1652),
.A2(n_1649),
.B(n_1651),
.C(n_1646),
.Y(n_1657)
);

AOI222xp33_ASAP7_75t_L g1658 ( 
.A1(n_1654),
.A2(n_1571),
.B1(n_1587),
.B2(n_1578),
.C1(n_1583),
.C2(n_1575),
.Y(n_1658)
);

OAI21xp33_ASAP7_75t_SL g1659 ( 
.A1(n_1648),
.A2(n_1566),
.B(n_1587),
.Y(n_1659)
);

AOI211xp5_ASAP7_75t_L g1660 ( 
.A1(n_1647),
.A2(n_1589),
.B(n_1499),
.C(n_1511),
.Y(n_1660)
);

OAI21xp33_ASAP7_75t_SL g1661 ( 
.A1(n_1650),
.A2(n_1589),
.B(n_1536),
.Y(n_1661)
);

AOI221xp5_ASAP7_75t_L g1662 ( 
.A1(n_1655),
.A2(n_1521),
.B1(n_1517),
.B2(n_1554),
.C(n_1499),
.Y(n_1662)
);

A2O1A1Ixp33_ASAP7_75t_L g1663 ( 
.A1(n_1657),
.A2(n_1511),
.B(n_1499),
.C(n_1554),
.Y(n_1663)
);

NOR3xp33_ASAP7_75t_SL g1664 ( 
.A(n_1659),
.B(n_1434),
.C(n_1415),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_SL g1665 ( 
.A(n_1661),
.B(n_1415),
.Y(n_1665)
);

AOI221x1_ASAP7_75t_SL g1666 ( 
.A1(n_1660),
.A2(n_1529),
.B1(n_1538),
.B2(n_1514),
.C(n_1547),
.Y(n_1666)
);

OAI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1662),
.A2(n_1656),
.B1(n_1533),
.B2(n_1536),
.Y(n_1667)
);

NOR3xp33_ASAP7_75t_L g1668 ( 
.A(n_1658),
.B(n_1392),
.C(n_1407),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1667),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1668),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1666),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1664),
.B(n_1415),
.Y(n_1672)
);

XOR2x2_ASAP7_75t_L g1673 ( 
.A(n_1665),
.B(n_1423),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1669),
.B(n_1663),
.Y(n_1674)
);

NOR3xp33_ASAP7_75t_L g1675 ( 
.A(n_1669),
.B(n_1670),
.C(n_1671),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1672),
.A2(n_1529),
.B(n_1514),
.Y(n_1676)
);

AOI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1676),
.A2(n_1673),
.B(n_1529),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1677),
.A2(n_1674),
.B1(n_1675),
.B2(n_1673),
.Y(n_1678)
);

OR2x6_ASAP7_75t_L g1679 ( 
.A(n_1678),
.B(n_1391),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_SL g1680 ( 
.A1(n_1678),
.A2(n_1434),
.B1(n_1413),
.B2(n_1391),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1679),
.Y(n_1681)
);

AOI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1680),
.A2(n_1538),
.B(n_1514),
.Y(n_1682)
);

AOI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1681),
.A2(n_1538),
.B(n_1541),
.Y(n_1683)
);

OAI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1682),
.A2(n_1540),
.B1(n_1551),
.B2(n_1549),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1683),
.B(n_1541),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1685),
.B(n_1684),
.Y(n_1686)
);

OAI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1686),
.A2(n_1552),
.B1(n_1551),
.B2(n_1549),
.Y(n_1687)
);

OAI221xp5_ASAP7_75t_R g1688 ( 
.A1(n_1687),
.A2(n_1552),
.B1(n_1547),
.B2(n_1545),
.C(n_1540),
.Y(n_1688)
);

AOI211xp5_ASAP7_75t_L g1689 ( 
.A1(n_1688),
.A2(n_1545),
.B(n_1401),
.C(n_1399),
.Y(n_1689)
);


endmodule