module fake_netlist_6_3873_n_1481 (n_52, n_1, n_91, n_256, n_209, n_63, n_223, n_278, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_56, n_119, n_235, n_147, n_191, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_53, n_44, n_232, n_16, n_163, n_46, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_152, n_92, n_321, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_231, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_215, n_178, n_247, n_225, n_308, n_309, n_317, n_149, n_90, n_24, n_54, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_315, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1481);

input n_52;
input n_1;
input n_91;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_152;
input n_92;
input n_321;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_231;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_317;
input n_149;
input n_90;
input n_24;
input n_54;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1481;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1415;
wire n_1370;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1393;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_1094;
wire n_953;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1339;
wire n_537;
wire n_1427;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_1429;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1443;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_942;
wire n_543;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1416;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_1311;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_339;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_241),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_268),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g325 ( 
.A(n_39),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_3),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_123),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_78),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_174),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_216),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_195),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_307),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_310),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_210),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_263),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_90),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_204),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_181),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_217),
.Y(n_339)
);

BUFx10_ASAP7_75t_L g340 ( 
.A(n_37),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_265),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_186),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_88),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_59),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_243),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_130),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_175),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_211),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_169),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_272),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_190),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_31),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_27),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_258),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_237),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_144),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_320),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_203),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_12),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_126),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_72),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_231),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_139),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_40),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_318),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_201),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_22),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_260),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_35),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_207),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_114),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_58),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_254),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_242),
.Y(n_374)
);

BUFx10_ASAP7_75t_L g375 ( 
.A(n_69),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_47),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_109),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_63),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_113),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_256),
.Y(n_380)
);

CKINVDCx14_ASAP7_75t_R g381 ( 
.A(n_51),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_167),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_292),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_249),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_51),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_37),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_25),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_108),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_12),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_42),
.Y(n_390)
);

BUFx8_ASAP7_75t_SL g391 ( 
.A(n_236),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_194),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_166),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_208),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_116),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_84),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_252),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_285),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_81),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_189),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_255),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_184),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_304),
.Y(n_403)
);

INVx2_ASAP7_75t_SL g404 ( 
.A(n_27),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_9),
.Y(n_405)
);

INVx2_ASAP7_75t_SL g406 ( 
.A(n_15),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_38),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_110),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_302),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_74),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_111),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_240),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_104),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_250),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_176),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_192),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_38),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_212),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_30),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_209),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_287),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_1),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_178),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_278),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_151),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_129),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_264),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_245),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_145),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_96),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_157),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_49),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_44),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_134),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_213),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_165),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_317),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_3),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_259),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_149),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_308),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_170),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_58),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_262),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_202),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_271),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_215),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_125),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_183),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_182),
.Y(n_450)
);

BUFx10_ASAP7_75t_L g451 ( 
.A(n_11),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_261),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_312),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_257),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_293),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_180),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_36),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_280),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_275),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_16),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_74),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_0),
.Y(n_462)
);

BUFx5_ASAP7_75t_L g463 ( 
.A(n_34),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_300),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_187),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_54),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_6),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_72),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_253),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_296),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_112),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_117),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_311),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_159),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_173),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_127),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_172),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_4),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_306),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_188),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_197),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_20),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_267),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_160),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_246),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_150),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_57),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_21),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_14),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_122),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_193),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_20),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_238),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_131),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_40),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_309),
.Y(n_496)
);

INVx1_ASAP7_75t_SL g497 ( 
.A(n_200),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_305),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_219),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_313),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_297),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_282),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_239),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_128),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_94),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_298),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_191),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_44),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_42),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_303),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_99),
.Y(n_511)
);

BUFx2_ASAP7_75t_SL g512 ( 
.A(n_315),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_9),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_66),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_79),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_322),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_266),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_269),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_98),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_155),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_137),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_163),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_156),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_224),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_223),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_161),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_286),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_140),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_23),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_52),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_87),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_26),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_281),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_85),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_34),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g536 ( 
.A(n_214),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_277),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_43),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_55),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_115),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_319),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_92),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_14),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_248),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_321),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_45),
.Y(n_546)
);

BUFx10_ASAP7_75t_L g547 ( 
.A(n_230),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_118),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_143),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_102),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_185),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_331),
.B(n_1),
.Y(n_552)
);

INVx5_ASAP7_75t_L g553 ( 
.A(n_338),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_381),
.B(n_2),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_338),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_463),
.Y(n_556)
);

BUFx8_ASAP7_75t_L g557 ( 
.A(n_430),
.Y(n_557)
);

INVx5_ASAP7_75t_L g558 ( 
.A(n_338),
.Y(n_558)
);

BUFx12f_ASAP7_75t_L g559 ( 
.A(n_340),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_381),
.B(n_2),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_463),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_353),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_338),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_331),
.B(n_4),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_536),
.B(n_5),
.Y(n_565)
);

INVx5_ASAP7_75t_L g566 ( 
.A(n_476),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_463),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_344),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_323),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_333),
.B(n_5),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_333),
.B(n_6),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_463),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_463),
.B(n_7),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_355),
.B(n_7),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_524),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_447),
.B(n_516),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_SL g577 ( 
.A(n_324),
.B(n_8),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_355),
.B(n_8),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_463),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_358),
.B(n_10),
.Y(n_580)
);

INVx5_ASAP7_75t_L g581 ( 
.A(n_476),
.Y(n_581)
);

INVx5_ASAP7_75t_L g582 ( 
.A(n_476),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_463),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_397),
.B(n_10),
.Y(n_584)
);

BUFx8_ASAP7_75t_SL g585 ( 
.A(n_391),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_476),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_344),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_344),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_420),
.B(n_11),
.Y(n_589)
);

BUFx8_ASAP7_75t_SL g590 ( 
.A(n_391),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_549),
.B(n_327),
.Y(n_591)
);

BUFx8_ASAP7_75t_SL g592 ( 
.A(n_457),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_344),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_352),
.Y(n_594)
);

INVx5_ASAP7_75t_L g595 ( 
.A(n_352),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_327),
.B(n_13),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_341),
.B(n_13),
.Y(n_597)
);

BUFx12f_ASAP7_75t_L g598 ( 
.A(n_340),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_401),
.B(n_16),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_341),
.B(n_17),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_352),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_401),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_352),
.Y(n_603)
);

BUFx12f_ASAP7_75t_L g604 ( 
.A(n_375),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_SL g605 ( 
.A(n_490),
.B(n_17),
.Y(n_605)
);

INVx5_ASAP7_75t_L g606 ( 
.A(n_547),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_359),
.Y(n_607)
);

INVx5_ASAP7_75t_L g608 ( 
.A(n_547),
.Y(n_608)
);

BUFx12f_ASAP7_75t_L g609 ( 
.A(n_375),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_393),
.B(n_18),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_415),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_393),
.B(n_18),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_494),
.B(n_496),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_494),
.B(n_19),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_415),
.B(n_21),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_483),
.B(n_22),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_483),
.B(n_23),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_496),
.B(n_24),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_520),
.B(n_334),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_328),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_326),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_520),
.B(n_24),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_335),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_422),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_372),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_342),
.B(n_25),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_547),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_329),
.Y(n_628)
);

INVx5_ASAP7_75t_L g629 ( 
.A(n_375),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_325),
.B(n_26),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_416),
.B(n_28),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_451),
.B(n_28),
.Y(n_632)
);

INVx5_ASAP7_75t_L g633 ( 
.A(n_451),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_497),
.B(n_29),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_343),
.B(n_347),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_378),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_348),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_330),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_404),
.B(n_29),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_356),
.B(n_30),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_357),
.B(n_31),
.Y(n_641)
);

INVx5_ASAP7_75t_L g642 ( 
.A(n_451),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_386),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_384),
.B(n_32),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_332),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_336),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_399),
.Y(n_647)
);

BUFx12f_ASAP7_75t_L g648 ( 
.A(n_361),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_408),
.B(n_409),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_414),
.B(n_32),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_418),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_422),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_424),
.B(n_33),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_487),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_431),
.B(n_33),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_435),
.B(n_35),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_440),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_445),
.B(n_39),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_465),
.B(n_41),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_471),
.B(n_41),
.Y(n_660)
);

INVx5_ASAP7_75t_L g661 ( 
.A(n_406),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_337),
.Y(n_662)
);

INVx5_ASAP7_75t_L g663 ( 
.A(n_487),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_509),
.B(n_43),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_514),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_475),
.Y(n_666)
);

INVx5_ASAP7_75t_L g667 ( 
.A(n_514),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_477),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_480),
.B(n_481),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_387),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_530),
.B(n_45),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_405),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_407),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_467),
.B(n_46),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_491),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_493),
.B(n_46),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_498),
.B(n_47),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_503),
.B(n_48),
.Y(n_678)
);

INVx4_ASAP7_75t_L g679 ( 
.A(n_339),
.Y(n_679)
);

INVx4_ASAP7_75t_L g680 ( 
.A(n_345),
.Y(n_680)
);

INVx5_ASAP7_75t_L g681 ( 
.A(n_535),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_535),
.B(n_48),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_504),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_433),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_505),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_438),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_510),
.B(n_49),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_443),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_460),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_521),
.B(n_50),
.Y(n_690)
);

INVx5_ASAP7_75t_L g691 ( 
.A(n_512),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_466),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_364),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_522),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_523),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_528),
.B(n_50),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_544),
.B(n_52),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_550),
.B(n_53),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_551),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_346),
.B(n_53),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_478),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_489),
.B(n_54),
.Y(n_702)
);

CKINVDCx6p67_ASAP7_75t_R g703 ( 
.A(n_380),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_349),
.B(n_56),
.Y(n_704)
);

INVx5_ASAP7_75t_L g705 ( 
.A(n_367),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_508),
.Y(n_706)
);

INVx5_ASAP7_75t_L g707 ( 
.A(n_369),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_376),
.B(n_56),
.Y(n_708)
);

OAI22xp33_ASAP7_75t_L g709 ( 
.A1(n_577),
.A2(n_385),
.B1(n_390),
.B2(n_389),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_SL g710 ( 
.A(n_605),
.B(n_380),
.Y(n_710)
);

OAI22xp33_ASAP7_75t_L g711 ( 
.A1(n_560),
.A2(n_419),
.B1(n_432),
.B2(n_410),
.Y(n_711)
);

OAI22xp33_ASAP7_75t_SL g712 ( 
.A1(n_576),
.A2(n_462),
.B1(n_468),
.B2(n_461),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_562),
.B(n_350),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_588),
.Y(n_714)
);

OAI22xp33_ASAP7_75t_L g715 ( 
.A1(n_606),
.A2(n_482),
.B1(n_495),
.B2(n_488),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_619),
.B(n_351),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_607),
.B(n_354),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_587),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_629),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_693),
.B(n_360),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_565),
.A2(n_400),
.B1(n_458),
.B2(n_392),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_587),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_593),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_606),
.B(n_362),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_601),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_608),
.B(n_363),
.Y(n_726)
);

INVx4_ASAP7_75t_L g727 ( 
.A(n_569),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_568),
.Y(n_728)
);

OAI22xp33_ASAP7_75t_SL g729 ( 
.A1(n_632),
.A2(n_589),
.B1(n_704),
.B2(n_591),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_627),
.B(n_532),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_568),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_608),
.B(n_365),
.Y(n_732)
);

AO22x2_ASAP7_75t_L g733 ( 
.A1(n_552),
.A2(n_529),
.B1(n_539),
.B2(n_513),
.Y(n_733)
);

OAI22xp33_ASAP7_75t_SL g734 ( 
.A1(n_552),
.A2(n_538),
.B1(n_546),
.B2(n_543),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_628),
.B(n_366),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_594),
.Y(n_736)
);

OAI22xp33_ASAP7_75t_L g737 ( 
.A1(n_596),
.A2(n_492),
.B1(n_417),
.B2(n_400),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_554),
.A2(n_458),
.B1(n_479),
.B2(n_392),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_631),
.A2(n_485),
.B1(n_479),
.B2(n_492),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_601),
.Y(n_740)
);

AO22x2_ASAP7_75t_L g741 ( 
.A1(n_564),
.A2(n_60),
.B1(n_57),
.B2(n_59),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_634),
.A2(n_485),
.B1(n_370),
.B2(n_371),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_638),
.B(n_368),
.Y(n_743)
);

OAI22xp33_ASAP7_75t_SL g744 ( 
.A1(n_564),
.A2(n_571),
.B1(n_578),
.B2(n_570),
.Y(n_744)
);

AO22x2_ASAP7_75t_L g745 ( 
.A1(n_570),
.A2(n_578),
.B1(n_599),
.B2(n_571),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_645),
.B(n_373),
.Y(n_746)
);

OA22x2_ASAP7_75t_L g747 ( 
.A1(n_688),
.A2(n_377),
.B1(n_379),
.B2(n_374),
.Y(n_747)
);

AO22x2_ASAP7_75t_L g748 ( 
.A1(n_599),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_662),
.B(n_382),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_648),
.A2(n_388),
.B1(n_394),
.B2(n_383),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_603),
.Y(n_751)
);

OAI22xp33_ASAP7_75t_L g752 ( 
.A1(n_597),
.A2(n_396),
.B1(n_398),
.B2(n_395),
.Y(n_752)
);

AO22x2_ASAP7_75t_L g753 ( 
.A1(n_615),
.A2(n_64),
.B1(n_61),
.B2(n_62),
.Y(n_753)
);

BUFx10_ASAP7_75t_L g754 ( 
.A(n_620),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_674),
.A2(n_584),
.B1(n_580),
.B2(n_708),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_559),
.A2(n_403),
.B1(n_411),
.B2(n_402),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_594),
.Y(n_757)
);

OAI22xp33_ASAP7_75t_SL g758 ( 
.A1(n_615),
.A2(n_413),
.B1(n_421),
.B2(n_412),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_629),
.B(n_423),
.Y(n_759)
);

NAND2xp33_ASAP7_75t_SL g760 ( 
.A(n_574),
.B(n_425),
.Y(n_760)
);

AO22x2_ASAP7_75t_L g761 ( 
.A1(n_616),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_555),
.Y(n_762)
);

OAI22xp33_ASAP7_75t_SL g763 ( 
.A1(n_573),
.A2(n_548),
.B1(n_545),
.B2(n_542),
.Y(n_763)
);

INVx8_ASAP7_75t_L g764 ( 
.A(n_585),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_617),
.B(n_426),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_691),
.B(n_427),
.Y(n_766)
);

OR2x2_ASAP7_75t_L g767 ( 
.A(n_602),
.B(n_65),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_629),
.B(n_428),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_555),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_633),
.B(n_429),
.Y(n_770)
);

AO22x2_ASAP7_75t_L g771 ( 
.A1(n_626),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_603),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_555),
.Y(n_773)
);

BUFx10_ASAP7_75t_L g774 ( 
.A(n_635),
.Y(n_774)
);

BUFx6f_ASAP7_75t_SL g775 ( 
.A(n_702),
.Y(n_775)
);

OAI22xp33_ASAP7_75t_L g776 ( 
.A1(n_600),
.A2(n_541),
.B1(n_540),
.B2(n_537),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_633),
.B(n_434),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_633),
.B(n_436),
.Y(n_778)
);

OAI22xp33_ASAP7_75t_SL g779 ( 
.A1(n_614),
.A2(n_534),
.B1(n_533),
.B2(n_531),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_642),
.B(n_437),
.Y(n_780)
);

OA22x2_ASAP7_75t_L g781 ( 
.A1(n_621),
.A2(n_527),
.B1(n_526),
.B2(n_525),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_642),
.B(n_439),
.Y(n_782)
);

OAI22xp33_ASAP7_75t_SL g783 ( 
.A1(n_622),
.A2(n_519),
.B1(n_518),
.B2(n_517),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_642),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_563),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_602),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_598),
.A2(n_515),
.B1(n_511),
.B2(n_507),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_586),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_705),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_602),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_646),
.B(n_441),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_646),
.B(n_442),
.Y(n_792)
);

AO22x2_ASAP7_75t_L g793 ( 
.A1(n_626),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_793)
);

AO22x2_ASAP7_75t_L g794 ( 
.A1(n_655),
.A2(n_696),
.B1(n_698),
.B2(n_690),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_604),
.A2(n_464),
.B1(n_502),
.B2(n_501),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_679),
.B(n_680),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_SL g797 ( 
.A1(n_575),
.A2(n_506),
.B1(n_500),
.B2(n_499),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_586),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_SL g799 ( 
.A1(n_641),
.A2(n_486),
.B1(n_484),
.B2(n_474),
.Y(n_799)
);

OAI22xp33_ASAP7_75t_L g800 ( 
.A1(n_640),
.A2(n_473),
.B1(n_472),
.B2(n_470),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_609),
.A2(n_452),
.B1(n_459),
.B2(n_456),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_700),
.A2(n_469),
.B1(n_455),
.B2(n_454),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_679),
.B(n_444),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_664),
.A2(n_453),
.B1(n_450),
.B2(n_449),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_680),
.B(n_446),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_561),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_561),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_806),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_806),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_744),
.A2(n_669),
.B(n_649),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_807),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_716),
.B(n_691),
.Y(n_812)
);

NAND2xp33_ASAP7_75t_R g813 ( 
.A(n_730),
.B(n_702),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_786),
.B(n_655),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_807),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_762),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_774),
.B(n_755),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_762),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_773),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_774),
.B(n_661),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_718),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_713),
.B(n_661),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_717),
.B(n_661),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_729),
.B(n_690),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_718),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_769),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_722),
.Y(n_827)
);

INVxp33_ASAP7_75t_L g828 ( 
.A(n_710),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_754),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_709),
.B(n_727),
.Y(n_830)
);

BUFx6f_ASAP7_75t_SL g831 ( 
.A(n_754),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_720),
.B(n_705),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_785),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_788),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_798),
.Y(n_835)
);

NAND2xp33_ASAP7_75t_R g836 ( 
.A(n_743),
.B(n_696),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_728),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_790),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_728),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_751),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_731),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_736),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_757),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_714),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_723),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_766),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_722),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_745),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_725),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_727),
.B(n_691),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_725),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_759),
.B(n_705),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_740),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_742),
.B(n_613),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_SL g855 ( 
.A(n_737),
.B(n_590),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_740),
.Y(n_856)
);

XOR2xp5_ASAP7_75t_L g857 ( 
.A(n_738),
.B(n_448),
.Y(n_857)
);

OR2x6_ASAP7_75t_L g858 ( 
.A(n_764),
.B(n_658),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_770),
.B(n_707),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_772),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_711),
.B(n_611),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_766),
.Y(n_862)
);

XOR2xp5_ASAP7_75t_L g863 ( 
.A(n_721),
.B(n_703),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_777),
.B(n_707),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_772),
.Y(n_865)
);

XOR2xp5_ASAP7_75t_L g866 ( 
.A(n_739),
.B(n_592),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_767),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_778),
.B(n_707),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_745),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_734),
.B(n_611),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_800),
.B(n_611),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_752),
.B(n_630),
.Y(n_872)
);

INVx1_ASAP7_75t_SL g873 ( 
.A(n_784),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_794),
.Y(n_874)
);

CKINVDCx20_ASAP7_75t_R g875 ( 
.A(n_797),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_794),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_780),
.B(n_671),
.Y(n_877)
);

NOR2xp67_ASAP7_75t_L g878 ( 
.A(n_802),
.B(n_553),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_733),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_735),
.Y(n_880)
);

AOI21x1_ASAP7_75t_L g881 ( 
.A1(n_796),
.A2(n_583),
.B(n_567),
.Y(n_881)
);

CKINVDCx16_ASAP7_75t_R g882 ( 
.A(n_775),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_743),
.B(n_698),
.Y(n_883)
);

XNOR2xp5_ASAP7_75t_L g884 ( 
.A(n_750),
.B(n_756),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_746),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_775),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_749),
.B(n_625),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_781),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_765),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_765),
.Y(n_890)
);

NOR2xp67_ASAP7_75t_L g891 ( 
.A(n_719),
.B(n_553),
.Y(n_891)
);

INVxp67_ASAP7_75t_SL g892 ( 
.A(n_741),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_749),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_747),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_815),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_848),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_839),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_844),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_893),
.B(n_763),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_845),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_820),
.B(n_828),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_877),
.B(n_791),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_849),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_851),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_828),
.B(n_782),
.Y(n_905)
);

INVx1_ASAP7_75t_SL g906 ( 
.A(n_873),
.Y(n_906)
);

AND2x2_ASAP7_75t_SL g907 ( 
.A(n_830),
.B(n_682),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_830),
.A2(n_760),
.B1(n_804),
.B2(n_776),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_822),
.B(n_792),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_823),
.B(n_803),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_854),
.B(n_758),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_810),
.B(n_805),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_854),
.B(n_712),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_831),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_808),
.B(n_724),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_893),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_815),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_821),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_809),
.B(n_726),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_872),
.A2(n_783),
.B(n_779),
.Y(n_920)
);

BUFx3_ASAP7_75t_L g921 ( 
.A(n_893),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_887),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_853),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_817),
.B(n_732),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_811),
.B(n_639),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_817),
.B(n_787),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_887),
.B(n_795),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_869),
.B(n_670),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_856),
.Y(n_929)
);

INVxp67_ASAP7_75t_SL g930 ( 
.A(n_821),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_867),
.B(n_801),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_832),
.B(n_789),
.Y(n_932)
);

INVxp67_ASAP7_75t_L g933 ( 
.A(n_813),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_825),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_860),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_883),
.B(n_741),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_865),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_848),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_893),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_814),
.B(n_636),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_825),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_827),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_872),
.B(n_799),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_847),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_847),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_883),
.B(n_748),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_814),
.B(n_643),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_846),
.B(n_672),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_824),
.B(n_583),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_846),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_874),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_841),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_824),
.B(n_768),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_876),
.B(n_861),
.Y(n_954)
);

INVxp67_ASAP7_75t_L g955 ( 
.A(n_813),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_862),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_862),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_836),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_840),
.Y(n_959)
);

INVx2_ASAP7_75t_SL g960 ( 
.A(n_837),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_837),
.B(n_812),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_894),
.Y(n_962)
);

AND2x4_ASAP7_75t_SL g963 ( 
.A(n_829),
.B(n_673),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_842),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_880),
.B(n_885),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_871),
.B(n_623),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_889),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_881),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_843),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_826),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_889),
.B(n_753),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_871),
.B(n_623),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_833),
.Y(n_973)
);

NAND2x1p5_ASAP7_75t_L g974 ( 
.A(n_890),
.B(n_556),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_852),
.B(n_623),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_859),
.B(n_637),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_864),
.B(n_637),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_834),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_870),
.B(n_753),
.Y(n_979)
);

INVxp67_ASAP7_75t_L g980 ( 
.A(n_836),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_879),
.B(n_686),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_835),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_888),
.A2(n_676),
.B(n_659),
.Y(n_983)
);

AND2x6_ASAP7_75t_L g984 ( 
.A(n_861),
.B(n_610),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_868),
.B(n_637),
.Y(n_985)
);

NAND2x1p5_ASAP7_75t_L g986 ( 
.A(n_916),
.B(n_838),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_981),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_895),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_948),
.B(n_886),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_906),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_901),
.B(n_882),
.Y(n_991)
);

INVx5_ASAP7_75t_L g992 ( 
.A(n_916),
.Y(n_992)
);

INVx5_ASAP7_75t_L g993 ( 
.A(n_916),
.Y(n_993)
);

OR2x2_ASAP7_75t_L g994 ( 
.A(n_943),
.B(n_857),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_965),
.B(n_892),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_895),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_917),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_916),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_930),
.B(n_892),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_896),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_930),
.B(n_850),
.Y(n_1001)
);

NAND2x1p5_ASAP7_75t_L g1002 ( 
.A(n_939),
.B(n_816),
.Y(n_1002)
);

AND2x6_ASAP7_75t_L g1003 ( 
.A(n_912),
.B(n_761),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_917),
.Y(n_1004)
);

AND2x4_ASAP7_75t_SL g1005 ( 
.A(n_939),
.B(n_858),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_958),
.B(n_980),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_896),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_918),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_939),
.Y(n_1009)
);

OR2x2_ASAP7_75t_L g1010 ( 
.A(n_938),
.B(n_863),
.Y(n_1010)
);

BUFx2_ASAP7_75t_L g1011 ( 
.A(n_938),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_924),
.B(n_905),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_907),
.B(n_850),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_939),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_918),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_907),
.B(n_878),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_954),
.B(n_884),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_933),
.B(n_955),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_934),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_933),
.B(n_858),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_934),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_948),
.B(n_858),
.Y(n_1022)
);

NAND2x1p5_ASAP7_75t_L g1023 ( 
.A(n_921),
.B(n_818),
.Y(n_1023)
);

BUFx12f_ASAP7_75t_L g1024 ( 
.A(n_914),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_954),
.B(n_771),
.Y(n_1025)
);

OR2x2_ASAP7_75t_L g1026 ( 
.A(n_926),
.B(n_866),
.Y(n_1026)
);

HB1xp67_ASAP7_75t_L g1027 ( 
.A(n_951),
.Y(n_1027)
);

INVx4_ASAP7_75t_L g1028 ( 
.A(n_950),
.Y(n_1028)
);

INVx6_ASAP7_75t_L g1029 ( 
.A(n_981),
.Y(n_1029)
);

INVx1_ASAP7_75t_SL g1030 ( 
.A(n_963),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_955),
.B(n_855),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_984),
.B(n_771),
.Y(n_1032)
);

NAND2x1p5_ASAP7_75t_L g1033 ( 
.A(n_921),
.B(n_819),
.Y(n_1033)
);

OR2x6_ASAP7_75t_L g1034 ( 
.A(n_936),
.B(n_793),
.Y(n_1034)
);

INVx4_ASAP7_75t_L g1035 ( 
.A(n_950),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_984),
.B(n_793),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_942),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_967),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_950),
.B(n_875),
.Y(n_1039)
);

NAND2x1p5_ASAP7_75t_L g1040 ( 
.A(n_950),
.B(n_572),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_956),
.Y(n_1041)
);

INVx3_ASAP7_75t_L g1042 ( 
.A(n_967),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_956),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_956),
.B(n_875),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_984),
.B(n_579),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_984),
.B(n_612),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_967),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_984),
.B(n_618),
.Y(n_1048)
);

CKINVDCx16_ASAP7_75t_R g1049 ( 
.A(n_946),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_956),
.B(n_684),
.Y(n_1050)
);

INVx6_ASAP7_75t_L g1051 ( 
.A(n_928),
.Y(n_1051)
);

NAND2x1p5_ASAP7_75t_L g1052 ( 
.A(n_957),
.B(n_891),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_909),
.B(n_701),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_944),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_944),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_949),
.B(n_677),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_910),
.B(n_701),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_941),
.Y(n_1058)
);

BUFx12f_ASAP7_75t_L g1059 ( 
.A(n_914),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_966),
.B(n_697),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_959),
.Y(n_1061)
);

OR2x6_ASAP7_75t_L g1062 ( 
.A(n_957),
.B(n_958),
.Y(n_1062)
);

INVx2_ASAP7_75t_SL g1063 ( 
.A(n_962),
.Y(n_1063)
);

OR2x2_ASAP7_75t_L g1064 ( 
.A(n_913),
.B(n_715),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_932),
.B(n_706),
.Y(n_1065)
);

INVx4_ASAP7_75t_L g1066 ( 
.A(n_992),
.Y(n_1066)
);

INVx6_ASAP7_75t_L g1067 ( 
.A(n_1041),
.Y(n_1067)
);

BUFx4_ASAP7_75t_SL g1068 ( 
.A(n_1034),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_990),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_1009),
.Y(n_1070)
);

INVx1_ASAP7_75t_SL g1071 ( 
.A(n_1000),
.Y(n_1071)
);

BUFx12f_ASAP7_75t_L g1072 ( 
.A(n_1024),
.Y(n_1072)
);

INVx5_ASAP7_75t_L g1073 ( 
.A(n_1009),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1006),
.B(n_980),
.Y(n_1074)
);

BUFx12f_ASAP7_75t_L g1075 ( 
.A(n_1059),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_996),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1015),
.Y(n_1077)
);

INVx2_ASAP7_75t_SL g1078 ( 
.A(n_1011),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1054),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_1039),
.Y(n_1080)
);

CKINVDCx16_ASAP7_75t_R g1081 ( 
.A(n_1049),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_1009),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_1012),
.Y(n_1083)
);

INVx8_ASAP7_75t_L g1084 ( 
.A(n_992),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_1039),
.Y(n_1085)
);

NAND2x1p5_ASAP7_75t_L g1086 ( 
.A(n_993),
.B(n_967),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_1014),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_1044),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_1041),
.Y(n_1089)
);

BUFx8_ASAP7_75t_SL g1090 ( 
.A(n_1044),
.Y(n_1090)
);

BUFx3_ASAP7_75t_L g1091 ( 
.A(n_989),
.Y(n_1091)
);

BUFx12f_ASAP7_75t_L g1092 ( 
.A(n_989),
.Y(n_1092)
);

INVx8_ASAP7_75t_L g1093 ( 
.A(n_993),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_1007),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_987),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_988),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1055),
.Y(n_1097)
);

INVx5_ASAP7_75t_SL g1098 ( 
.A(n_1022),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_1041),
.Y(n_1099)
);

BUFx12f_ASAP7_75t_L g1100 ( 
.A(n_1022),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_997),
.Y(n_1101)
);

BUFx12f_ASAP7_75t_L g1102 ( 
.A(n_1063),
.Y(n_1102)
);

OR2x2_ASAP7_75t_L g1103 ( 
.A(n_1017),
.B(n_902),
.Y(n_1103)
);

INVx4_ASAP7_75t_L g1104 ( 
.A(n_993),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_1043),
.Y(n_1105)
);

INVx4_ASAP7_75t_L g1106 ( 
.A(n_993),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_1050),
.B(n_922),
.Y(n_1107)
);

BUFx12f_ASAP7_75t_L g1108 ( 
.A(n_1010),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_1014),
.Y(n_1109)
);

NAND2x1p5_ASAP7_75t_L g1110 ( 
.A(n_1028),
.B(n_960),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_1014),
.Y(n_1111)
);

INVx5_ASAP7_75t_L g1112 ( 
.A(n_1043),
.Y(n_1112)
);

CKINVDCx16_ASAP7_75t_R g1113 ( 
.A(n_991),
.Y(n_1113)
);

INVx4_ASAP7_75t_L g1114 ( 
.A(n_1043),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_995),
.Y(n_1115)
);

INVx4_ASAP7_75t_L g1116 ( 
.A(n_1028),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_1062),
.Y(n_1117)
);

NAND2x1p5_ASAP7_75t_L g1118 ( 
.A(n_1035),
.B(n_982),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1004),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_1029),
.Y(n_1120)
);

INVx2_ASAP7_75t_SL g1121 ( 
.A(n_1029),
.Y(n_1121)
);

BUFx4f_ASAP7_75t_L g1122 ( 
.A(n_1018),
.Y(n_1122)
);

INVx4_ASAP7_75t_L g1123 ( 
.A(n_1035),
.Y(n_1123)
);

CKINVDCx16_ASAP7_75t_R g1124 ( 
.A(n_1026),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1008),
.Y(n_1125)
);

INVx6_ASAP7_75t_L g1126 ( 
.A(n_1051),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_1031),
.Y(n_1127)
);

BUFx12f_ASAP7_75t_L g1128 ( 
.A(n_1034),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1019),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1021),
.Y(n_1130)
);

INVx1_ASAP7_75t_SL g1131 ( 
.A(n_1027),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_1070),
.Y(n_1132)
);

OAI21xp33_ASAP7_75t_L g1133 ( 
.A1(n_1103),
.A2(n_1017),
.B(n_911),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1074),
.B(n_1006),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1074),
.B(n_999),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1076),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1096),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_1127),
.A2(n_911),
.B1(n_994),
.B2(n_1064),
.Y(n_1138)
);

INVx2_ASAP7_75t_SL g1139 ( 
.A(n_1069),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1066),
.A2(n_1001),
.B(n_1045),
.Y(n_1140)
);

AOI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1083),
.A2(n_1013),
.B1(n_908),
.B2(n_1003),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1077),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1079),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_1083),
.B(n_1053),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1096),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1097),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_L g1147 ( 
.A1(n_1122),
.A2(n_1003),
.B1(n_1013),
.B2(n_920),
.Y(n_1147)
);

CKINVDCx11_ASAP7_75t_R g1148 ( 
.A(n_1072),
.Y(n_1148)
);

BUFx10_ASAP7_75t_L g1149 ( 
.A(n_1078),
.Y(n_1149)
);

AOI22xp33_ASAP7_75t_SL g1150 ( 
.A1(n_1113),
.A2(n_557),
.B1(n_1003),
.B2(n_1025),
.Y(n_1150)
);

BUFx3_ASAP7_75t_L g1151 ( 
.A(n_1069),
.Y(n_1151)
);

AOI22xp33_ASAP7_75t_SL g1152 ( 
.A1(n_1080),
.A2(n_1085),
.B1(n_1088),
.B2(n_1124),
.Y(n_1152)
);

CKINVDCx20_ASAP7_75t_R g1153 ( 
.A(n_1081),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1101),
.Y(n_1154)
);

BUFx8_ASAP7_75t_L g1155 ( 
.A(n_1075),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_1108),
.Y(n_1156)
);

INVx6_ASAP7_75t_L g1157 ( 
.A(n_1102),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1115),
.B(n_999),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1119),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1129),
.Y(n_1160)
);

INVx5_ASAP7_75t_L g1161 ( 
.A(n_1084),
.Y(n_1161)
);

AOI22xp33_ASAP7_75t_L g1162 ( 
.A1(n_1107),
.A2(n_1020),
.B1(n_1016),
.B2(n_931),
.Y(n_1162)
);

CKINVDCx11_ASAP7_75t_R g1163 ( 
.A(n_1092),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_SL g1164 ( 
.A1(n_1107),
.A2(n_979),
.B1(n_1036),
.B2(n_1032),
.Y(n_1164)
);

INVx3_ASAP7_75t_SL g1165 ( 
.A(n_1071),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1117),
.A2(n_1016),
.B1(n_1036),
.B2(n_1032),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1117),
.A2(n_1051),
.B1(n_927),
.B2(n_962),
.Y(n_1167)
);

CKINVDCx6p67_ASAP7_75t_R g1168 ( 
.A(n_1100),
.Y(n_1168)
);

CKINVDCx14_ASAP7_75t_R g1169 ( 
.A(n_1095),
.Y(n_1169)
);

INVx4_ASAP7_75t_L g1170 ( 
.A(n_1084),
.Y(n_1170)
);

INVx4_ASAP7_75t_L g1171 ( 
.A(n_1084),
.Y(n_1171)
);

INVx2_ASAP7_75t_SL g1172 ( 
.A(n_1094),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1125),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_1095),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1130),
.Y(n_1175)
);

OAI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1131),
.A2(n_1030),
.B1(n_1062),
.B2(n_953),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_SL g1177 ( 
.A1(n_1131),
.A2(n_1005),
.B1(n_963),
.B2(n_1057),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1070),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1117),
.Y(n_1179)
);

BUFx2_ASAP7_75t_L g1180 ( 
.A(n_1090),
.Y(n_1180)
);

NAND2x1p5_ASAP7_75t_L g1181 ( 
.A(n_1112),
.B(n_998),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1089),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_L g1183 ( 
.A1(n_1091),
.A2(n_1050),
.B1(n_1048),
.B2(n_1046),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1126),
.A2(n_971),
.B1(n_1048),
.B2(n_1046),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1091),
.B(n_1065),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1098),
.A2(n_940),
.B1(n_947),
.B2(n_899),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_1070),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1098),
.A2(n_940),
.B1(n_947),
.B2(n_899),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1086),
.A2(n_1056),
.B1(n_1060),
.B2(n_972),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1099),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1098),
.A2(n_928),
.B1(n_1061),
.B2(n_959),
.Y(n_1191)
);

AO22x1_ASAP7_75t_L g1192 ( 
.A1(n_1120),
.A2(n_928),
.B1(n_983),
.B2(n_1058),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1086),
.A2(n_1056),
.B1(n_1060),
.B2(n_903),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1099),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1126),
.B(n_951),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_SL g1196 ( 
.A1(n_1144),
.A2(n_1128),
.B1(n_1126),
.B2(n_644),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_1132),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1138),
.B(n_1121),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1173),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_1132),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1133),
.A2(n_653),
.B1(n_656),
.B2(n_650),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1133),
.A2(n_678),
.B1(n_687),
.B2(n_660),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1185),
.B(n_904),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1134),
.A2(n_1090),
.B1(n_929),
.B2(n_935),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_1134),
.B(n_915),
.Y(n_1205)
);

INVx6_ASAP7_75t_L g1206 ( 
.A(n_1161),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1158),
.B(n_919),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1136),
.Y(n_1208)
);

BUFx4f_ASAP7_75t_SL g1209 ( 
.A(n_1155),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1141),
.B(n_923),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1142),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1143),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1164),
.B(n_937),
.Y(n_1213)
);

INVx3_ASAP7_75t_L g1214 ( 
.A(n_1170),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1175),
.Y(n_1215)
);

OAI21xp33_ASAP7_75t_L g1216 ( 
.A1(n_1162),
.A2(n_900),
.B(n_898),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_1146),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1141),
.B(n_897),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1150),
.A2(n_952),
.B1(n_969),
.B2(n_964),
.Y(n_1219)
);

OAI21xp33_ASAP7_75t_L g1220 ( 
.A1(n_1167),
.A2(n_925),
.B(n_973),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1154),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_1132),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1152),
.B(n_970),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1147),
.A2(n_1118),
.B1(n_1110),
.B2(n_986),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1160),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_SL g1226 ( 
.A1(n_1177),
.A2(n_1052),
.B(n_961),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1193),
.A2(n_689),
.B1(n_692),
.B2(n_684),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1165),
.B(n_1105),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_SL g1229 ( 
.A1(n_1153),
.A2(n_1093),
.B1(n_1118),
.B2(n_1110),
.Y(n_1229)
);

BUFx2_ASAP7_75t_L g1230 ( 
.A(n_1151),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1159),
.Y(n_1231)
);

AOI21xp33_ASAP7_75t_L g1232 ( 
.A1(n_1193),
.A2(n_1045),
.B(n_976),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1166),
.A2(n_986),
.B1(n_1052),
.B2(n_1042),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1135),
.A2(n_692),
.B1(n_978),
.B2(n_945),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_SL g1235 ( 
.A1(n_1169),
.A2(n_1093),
.B1(n_1112),
.B2(n_1073),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_1172),
.Y(n_1236)
);

OAI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1184),
.A2(n_1037),
.B1(n_1112),
.B2(n_1042),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_SL g1238 ( 
.A1(n_1180),
.A2(n_1093),
.B1(n_1112),
.B2(n_1073),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1195),
.B(n_1105),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_1174),
.Y(n_1240)
);

OAI21xp33_ASAP7_75t_L g1241 ( 
.A1(n_1186),
.A2(n_977),
.B(n_975),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1137),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1189),
.A2(n_706),
.B1(n_647),
.B2(n_651),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1145),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1182),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_1179),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_1192),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1176),
.B(n_985),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1188),
.A2(n_1038),
.B1(n_1047),
.B2(n_1073),
.Y(n_1249)
);

BUFx8_ASAP7_75t_SL g1250 ( 
.A(n_1156),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1190),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1189),
.A2(n_683),
.B1(n_647),
.B2(n_651),
.Y(n_1252)
);

INVx4_ASAP7_75t_L g1253 ( 
.A(n_1161),
.Y(n_1253)
);

NAND3xp33_ASAP7_75t_L g1254 ( 
.A(n_1183),
.B(n_651),
.C(n_647),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1139),
.B(n_1194),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1203),
.B(n_1149),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1210),
.A2(n_1191),
.B1(n_1157),
.B2(n_1168),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1198),
.A2(n_1163),
.B1(n_1148),
.B2(n_1155),
.Y(n_1258)
);

OAI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1219),
.A2(n_1140),
.B1(n_1171),
.B2(n_1123),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1205),
.B(n_1187),
.Y(n_1260)
);

AOI221xp5_ASAP7_75t_L g1261 ( 
.A1(n_1201),
.A2(n_665),
.B1(n_654),
.B2(n_694),
.C(n_657),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1204),
.A2(n_1171),
.B1(n_1033),
.B2(n_1023),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1217),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1210),
.A2(n_974),
.B1(n_1040),
.B2(n_1047),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1239),
.B(n_1178),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1216),
.A2(n_974),
.B1(n_1040),
.B2(n_1038),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1204),
.A2(n_1023),
.B1(n_1033),
.B2(n_1181),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1217),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1223),
.B(n_1178),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1201),
.A2(n_1067),
.B1(n_1178),
.B2(n_1187),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1208),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1202),
.A2(n_1067),
.B1(n_1187),
.B2(n_998),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1202),
.A2(n_1116),
.B1(n_683),
.B2(n_699),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1220),
.A2(n_683),
.B1(n_657),
.B2(n_666),
.Y(n_1274)
);

OAI221xp5_ASAP7_75t_L g1275 ( 
.A1(n_1196),
.A2(n_654),
.B1(n_665),
.B2(n_1002),
.C(n_652),
.Y(n_1275)
);

AOI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1248),
.A2(n_968),
.B(n_1002),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_SL g1277 ( 
.A1(n_1247),
.A2(n_1114),
.B1(n_685),
.B2(n_699),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1218),
.A2(n_685),
.B1(n_657),
.B2(n_666),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1228),
.B(n_1082),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1205),
.B(n_1082),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1207),
.B(n_1082),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1213),
.A2(n_685),
.B1(n_699),
.B2(n_695),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1199),
.B(n_1087),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1247),
.A2(n_668),
.B1(n_675),
.B2(n_694),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1255),
.B(n_1087),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1241),
.A2(n_668),
.B1(n_675),
.B2(n_694),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1254),
.A2(n_675),
.B1(n_695),
.B2(n_1111),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1215),
.Y(n_1288)
);

OAI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1209),
.A2(n_1111),
.B1(n_1109),
.B2(n_1087),
.Y(n_1289)
);

OAI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1209),
.A2(n_1212),
.B1(n_1211),
.B2(n_1221),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1225),
.B(n_1109),
.Y(n_1291)
);

AOI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1226),
.A2(n_695),
.B1(n_624),
.B2(n_1111),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1236),
.B(n_1109),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1236),
.A2(n_968),
.B1(n_1104),
.B2(n_1066),
.Y(n_1294)
);

OAI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1231),
.A2(n_1068),
.B1(n_1104),
.B2(n_1106),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1242),
.B(n_70),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1245),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1227),
.A2(n_681),
.B1(n_667),
.B2(n_663),
.Y(n_1298)
);

OA21x2_ASAP7_75t_L g1299 ( 
.A1(n_1232),
.A2(n_71),
.B(n_73),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1237),
.A2(n_681),
.B1(n_667),
.B2(n_663),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_SL g1301 ( 
.A1(n_1224),
.A2(n_581),
.B1(n_558),
.B2(n_566),
.Y(n_1301)
);

AOI221xp5_ASAP7_75t_L g1302 ( 
.A1(n_1243),
.A2(n_71),
.B1(n_75),
.B2(n_76),
.C(n_595),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1237),
.A2(n_595),
.B1(n_582),
.B2(n_581),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1229),
.A2(n_582),
.B1(n_581),
.B2(n_566),
.Y(n_1304)
);

OAI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1230),
.A2(n_75),
.B1(n_582),
.B2(n_566),
.Y(n_1305)
);

OAI21xp33_ASAP7_75t_SL g1306 ( 
.A1(n_1252),
.A2(n_77),
.B(n_80),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1234),
.A2(n_595),
.B1(n_558),
.B2(n_553),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_SL g1308 ( 
.A1(n_1233),
.A2(n_1206),
.B1(n_1240),
.B2(n_1249),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1234),
.A2(n_1243),
.B1(n_1240),
.B2(n_1246),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1246),
.A2(n_558),
.B1(n_83),
.B2(n_86),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1244),
.A2(n_82),
.B1(n_89),
.B2(n_91),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_SL g1312 ( 
.A1(n_1206),
.A2(n_93),
.B1(n_95),
.B2(n_97),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_SL g1313 ( 
.A1(n_1206),
.A2(n_100),
.B1(n_101),
.B2(n_103),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1238),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1271),
.B(n_1251),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1280),
.B(n_1197),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1290),
.B(n_1235),
.Y(n_1317)
);

AND2x2_ASAP7_75t_SL g1318 ( 
.A(n_1299),
.B(n_1253),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1260),
.B(n_1197),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1297),
.B(n_1197),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1268),
.B(n_1197),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1263),
.B(n_1200),
.Y(n_1322)
);

OR2x2_ASAP7_75t_L g1323 ( 
.A(n_1263),
.B(n_1200),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1281),
.B(n_1200),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_SL g1325 ( 
.A(n_1290),
.B(n_1214),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1288),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1269),
.B(n_1200),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1265),
.B(n_1222),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1276),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1299),
.B(n_1222),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1256),
.B(n_1222),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1299),
.B(n_119),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_SL g1333 ( 
.A(n_1257),
.B(n_1250),
.Y(n_1333)
);

NAND4xp25_ASAP7_75t_L g1334 ( 
.A(n_1302),
.B(n_120),
.C(n_121),
.D(n_124),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1309),
.A2(n_132),
.B1(n_133),
.B2(n_135),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1285),
.B(n_1293),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1296),
.B(n_136),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1279),
.B(n_138),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1283),
.B(n_141),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1305),
.A2(n_142),
.B1(n_146),
.B2(n_147),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1308),
.B(n_148),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1291),
.B(n_152),
.Y(n_1342)
);

NAND3xp33_ASAP7_75t_L g1343 ( 
.A(n_1305),
.B(n_153),
.C(n_154),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1292),
.B(n_158),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1275),
.A2(n_162),
.B1(n_164),
.B2(n_168),
.Y(n_1345)
);

NAND4xp25_ASAP7_75t_SL g1346 ( 
.A(n_1258),
.B(n_171),
.C(n_177),
.D(n_179),
.Y(n_1346)
);

AOI221xp5_ASAP7_75t_L g1347 ( 
.A1(n_1261),
.A2(n_1282),
.B1(n_1295),
.B2(n_1304),
.C(n_1311),
.Y(n_1347)
);

AOI211xp5_ASAP7_75t_L g1348 ( 
.A1(n_1314),
.A2(n_196),
.B(n_198),
.C(n_199),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1311),
.B(n_205),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1301),
.B(n_206),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1300),
.B(n_218),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1303),
.B(n_220),
.Y(n_1352)
);

OAI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1306),
.A2(n_221),
.B(n_222),
.Y(n_1353)
);

NAND3xp33_ASAP7_75t_L g1354 ( 
.A(n_1273),
.B(n_225),
.C(n_226),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1259),
.B(n_1270),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1321),
.B(n_1286),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1323),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1323),
.B(n_1262),
.Y(n_1358)
);

AO21x2_ASAP7_75t_L g1359 ( 
.A1(n_1329),
.A2(n_1289),
.B(n_1267),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1321),
.B(n_1274),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1315),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1326),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1330),
.B(n_1264),
.Y(n_1363)
);

AND2x4_ASAP7_75t_L g1364 ( 
.A(n_1322),
.B(n_1272),
.Y(n_1364)
);

NOR3xp33_ASAP7_75t_L g1365 ( 
.A(n_1343),
.B(n_1313),
.C(n_1312),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1330),
.B(n_1322),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1336),
.B(n_1310),
.Y(n_1367)
);

NOR2x1_ASAP7_75t_L g1368 ( 
.A(n_1331),
.B(n_1289),
.Y(n_1368)
);

NAND4xp75_ASAP7_75t_L g1369 ( 
.A(n_1317),
.B(n_1277),
.C(n_1287),
.D(n_1284),
.Y(n_1369)
);

OR2x2_ASAP7_75t_L g1370 ( 
.A(n_1329),
.B(n_1278),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1326),
.B(n_1316),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1336),
.B(n_1294),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1324),
.B(n_1266),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1334),
.A2(n_1349),
.B1(n_1346),
.B2(n_1347),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1319),
.B(n_1307),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1320),
.Y(n_1376)
);

NOR3xp33_ASAP7_75t_L g1377 ( 
.A(n_1334),
.B(n_1298),
.C(n_227),
.Y(n_1377)
);

AO22x1_ASAP7_75t_L g1378 ( 
.A1(n_1332),
.A2(n_228),
.B1(n_229),
.B2(n_232),
.Y(n_1378)
);

NAND3xp33_ASAP7_75t_L g1379 ( 
.A(n_1348),
.B(n_1340),
.C(n_1341),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1327),
.B(n_1328),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1318),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1332),
.Y(n_1382)
);

AO21x2_ASAP7_75t_L g1383 ( 
.A1(n_1355),
.A2(n_233),
.B(n_234),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1318),
.B(n_235),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1362),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1362),
.Y(n_1386)
);

XOR2xp5_ASAP7_75t_L g1387 ( 
.A(n_1374),
.B(n_1333),
.Y(n_1387)
);

INVx2_ASAP7_75t_SL g1388 ( 
.A(n_1366),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1361),
.Y(n_1389)
);

INVxp67_ASAP7_75t_SL g1390 ( 
.A(n_1357),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1382),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1371),
.Y(n_1392)
);

INVx2_ASAP7_75t_SL g1393 ( 
.A(n_1376),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1381),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1380),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1358),
.Y(n_1396)
);

NAND4xp75_ASAP7_75t_L g1397 ( 
.A(n_1384),
.B(n_1353),
.C(n_1325),
.D(n_1350),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1363),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1363),
.B(n_1328),
.Y(n_1399)
);

INVxp67_ASAP7_75t_SL g1400 ( 
.A(n_1368),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1384),
.B(n_1338),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1359),
.Y(n_1402)
);

INVx1_ASAP7_75t_SL g1403 ( 
.A(n_1372),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1370),
.Y(n_1404)
);

XNOR2xp5_ASAP7_75t_L g1405 ( 
.A(n_1374),
.B(n_1338),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1359),
.Y(n_1406)
);

XNOR2xp5_ASAP7_75t_L g1407 ( 
.A(n_1387),
.B(n_1367),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_1404),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1390),
.Y(n_1409)
);

INVxp67_ASAP7_75t_L g1410 ( 
.A(n_1400),
.Y(n_1410)
);

XOR2x2_ASAP7_75t_L g1411 ( 
.A(n_1387),
.B(n_1379),
.Y(n_1411)
);

AO22x2_ASAP7_75t_L g1412 ( 
.A1(n_1406),
.A2(n_1369),
.B1(n_1365),
.B2(n_1377),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1393),
.Y(n_1413)
);

INVx1_ASAP7_75t_SL g1414 ( 
.A(n_1403),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1393),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1405),
.B(n_1401),
.Y(n_1416)
);

AO22x2_ASAP7_75t_L g1417 ( 
.A1(n_1397),
.A2(n_1373),
.B1(n_1364),
.B2(n_1354),
.Y(n_1417)
);

INVx1_ASAP7_75t_SL g1418 ( 
.A(n_1398),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1391),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1389),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1385),
.Y(n_1421)
);

INVxp67_ASAP7_75t_L g1422 ( 
.A(n_1398),
.Y(n_1422)
);

XOR2x2_ASAP7_75t_L g1423 ( 
.A(n_1405),
.B(n_1367),
.Y(n_1423)
);

XNOR2xp5_ASAP7_75t_L g1424 ( 
.A(n_1401),
.B(n_1372),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1386),
.Y(n_1425)
);

INVx1_ASAP7_75t_SL g1426 ( 
.A(n_1414),
.Y(n_1426)
);

INVxp67_ASAP7_75t_L g1427 ( 
.A(n_1416),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1422),
.Y(n_1428)
);

AOI22x1_ASAP7_75t_SL g1429 ( 
.A1(n_1411),
.A2(n_1396),
.B1(n_1402),
.B2(n_1391),
.Y(n_1429)
);

OA22x2_ASAP7_75t_L g1430 ( 
.A1(n_1407),
.A2(n_1424),
.B1(n_1410),
.B2(n_1422),
.Y(n_1430)
);

AO22x2_ASAP7_75t_L g1431 ( 
.A1(n_1410),
.A2(n_1418),
.B1(n_1415),
.B2(n_1413),
.Y(n_1431)
);

OA22x2_ASAP7_75t_L g1432 ( 
.A1(n_1409),
.A2(n_1388),
.B1(n_1394),
.B2(n_1399),
.Y(n_1432)
);

OA22x2_ASAP7_75t_L g1433 ( 
.A1(n_1423),
.A2(n_1388),
.B1(n_1399),
.B2(n_1395),
.Y(n_1433)
);

INVx2_ASAP7_75t_SL g1434 ( 
.A(n_1408),
.Y(n_1434)
);

XNOR2x1_ASAP7_75t_L g1435 ( 
.A(n_1412),
.B(n_1378),
.Y(n_1435)
);

AOI22x1_ASAP7_75t_L g1436 ( 
.A1(n_1412),
.A2(n_1350),
.B1(n_1402),
.B2(n_1352),
.Y(n_1436)
);

AOI22x1_ASAP7_75t_L g1437 ( 
.A1(n_1412),
.A2(n_1352),
.B1(n_1351),
.B2(n_1392),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1413),
.B(n_1364),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1421),
.Y(n_1439)
);

INVx1_ASAP7_75t_SL g1440 ( 
.A(n_1435),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1438),
.Y(n_1441)
);

OA22x2_ASAP7_75t_L g1442 ( 
.A1(n_1427),
.A2(n_1417),
.B1(n_1415),
.B2(n_1419),
.Y(n_1442)
);

OAI322xp33_ASAP7_75t_L g1443 ( 
.A1(n_1430),
.A2(n_1419),
.A3(n_1420),
.B1(n_1425),
.B2(n_1417),
.C1(n_1375),
.C2(n_1337),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1428),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1439),
.Y(n_1445)
);

INVx1_ASAP7_75t_SL g1446 ( 
.A(n_1426),
.Y(n_1446)
);

INVx1_ASAP7_75t_SL g1447 ( 
.A(n_1429),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1431),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1431),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1445),
.Y(n_1450)
);

NAND4xp75_ASAP7_75t_L g1451 ( 
.A(n_1448),
.B(n_1429),
.C(n_1434),
.D(n_1436),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1447),
.A2(n_1437),
.B1(n_1436),
.B2(n_1417),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1444),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1449),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1453),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1454),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1450),
.Y(n_1457)
);

O2A1O1Ixp33_ASAP7_75t_L g1458 ( 
.A1(n_1452),
.A2(n_1447),
.B(n_1440),
.C(n_1443),
.Y(n_1458)
);

OA22x2_ASAP7_75t_L g1459 ( 
.A1(n_1451),
.A2(n_1440),
.B1(n_1446),
.B2(n_1441),
.Y(n_1459)
);

NAND4xp25_ASAP7_75t_SL g1460 ( 
.A(n_1458),
.B(n_1456),
.C(n_1442),
.D(n_1455),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1457),
.B(n_1433),
.Y(n_1461)
);

AOI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1459),
.A2(n_1432),
.B1(n_1383),
.B2(n_1360),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1461),
.Y(n_1463)
);

AOI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1460),
.A2(n_1383),
.B1(n_1356),
.B2(n_1359),
.Y(n_1464)
);

OR3x2_ASAP7_75t_L g1465 ( 
.A(n_1463),
.B(n_1462),
.C(n_1335),
.Y(n_1465)
);

NOR4xp25_ASAP7_75t_L g1466 ( 
.A(n_1464),
.B(n_1354),
.C(n_1339),
.D(n_1342),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1465),
.Y(n_1467)
);

INVx3_ASAP7_75t_L g1468 ( 
.A(n_1466),
.Y(n_1468)
);

AOI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1467),
.A2(n_1351),
.B1(n_1344),
.B2(n_1345),
.Y(n_1469)
);

AOI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1468),
.A2(n_244),
.B1(n_247),
.B2(n_251),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1469),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1470),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1472),
.A2(n_270),
.B1(n_273),
.B2(n_274),
.Y(n_1473)
);

OAI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1471),
.A2(n_276),
.B1(n_279),
.B2(n_283),
.Y(n_1474)
);

INVxp67_ASAP7_75t_SL g1475 ( 
.A(n_1474),
.Y(n_1475)
);

OAI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1475),
.A2(n_1473),
.B1(n_288),
.B2(n_289),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1475),
.A2(n_284),
.B1(n_290),
.B2(n_291),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1477),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1476),
.Y(n_1479)
);

AOI221xp5_ASAP7_75t_L g1480 ( 
.A1(n_1479),
.A2(n_294),
.B1(n_295),
.B2(n_299),
.C(n_301),
.Y(n_1480)
);

AOI211xp5_ASAP7_75t_L g1481 ( 
.A1(n_1480),
.A2(n_1478),
.B(n_314),
.C(n_316),
.Y(n_1481)
);


endmodule