module fake_netlist_5_1294_n_1863 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1863);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1863;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_770;
wire n_458;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1835;
wire n_1726;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_190),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_75),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_39),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_164),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_62),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_5),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_154),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_161),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_121),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_10),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_5),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_76),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_12),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_38),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_98),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_141),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_136),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_104),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_173),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_122),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_149),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g214 ( 
.A(n_42),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_54),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_94),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_115),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_14),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_81),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_116),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_67),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_177),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_157),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_78),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_156),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_107),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_179),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_38),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_112),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_146),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_43),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_2),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_117),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_150),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_137),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_96),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_108),
.Y(n_237)
);

BUFx5_ASAP7_75t_L g238 ( 
.A(n_25),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_41),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_138),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_12),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_165),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_34),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_131),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_144),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_135),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_24),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_180),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_176),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_1),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_129),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_39),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_14),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_128),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_44),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_124),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_63),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_7),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_85),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_97),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_52),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_53),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_101),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_152),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_184),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_187),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_16),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_43),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_174),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_182),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_110),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_132),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_123),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_130),
.Y(n_274)
);

BUFx10_ASAP7_75t_L g275 ( 
.A(n_27),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_84),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_58),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_178),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_189),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_28),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_69),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_83),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_3),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_18),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_181),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_44),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_10),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_92),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_171),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_72),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_0),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_51),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_118),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_162),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_183),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_61),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_11),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_66),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_59),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_11),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_175),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_56),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_17),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_170),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_6),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_160),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_86),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_147),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_37),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_155),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_169),
.Y(n_311)
);

BUFx10_ASAP7_75t_L g312 ( 
.A(n_172),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_139),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_99),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_163),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_53),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_168),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_79),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_8),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_191),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_17),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_34),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_113),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_26),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_19),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_102),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_80),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_145),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_40),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_73),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_143),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_100),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_114),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_185),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_33),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_28),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_186),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_59),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_8),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_13),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_49),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_32),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_18),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_49),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_127),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_27),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_30),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_167),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_54),
.Y(n_349)
);

BUFx10_ASAP7_75t_L g350 ( 
.A(n_52),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_6),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_41),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_45),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_90),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_64),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_48),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_9),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_51),
.Y(n_358)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_23),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_22),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_46),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_31),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_140),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_1),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_88),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_23),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_134),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_7),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_31),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_4),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_40),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_56),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_77),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_13),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_89),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_87),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_21),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_70),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_103),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_133),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_48),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_26),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_71),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_153),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_238),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_238),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_243),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g388 ( 
.A(n_294),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_192),
.Y(n_389)
);

INVxp33_ASAP7_75t_L g390 ( 
.A(n_302),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_238),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_238),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_238),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_198),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_225),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_238),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_238),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_201),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_259),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_226),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_238),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_227),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_202),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_202),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_202),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_202),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_202),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_325),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_325),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_229),
.Y(n_410)
);

BUFx10_ASAP7_75t_L g411 ( 
.A(n_375),
.Y(n_411)
);

INVxp67_ASAP7_75t_SL g412 ( 
.A(n_219),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_267),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_359),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_325),
.Y(n_415)
);

INVxp33_ASAP7_75t_SL g416 ( 
.A(n_372),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_260),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_230),
.Y(n_418)
);

INVxp33_ASAP7_75t_SL g419 ( 
.A(n_194),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_325),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_194),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_234),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_325),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_357),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_235),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_300),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_214),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_278),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_357),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_300),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_203),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_217),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_222),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_357),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g435 ( 
.A(n_217),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_357),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_357),
.Y(n_437)
);

INVxp33_ASAP7_75t_SL g438 ( 
.A(n_203),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_240),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_358),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_358),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_358),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_358),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_358),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_288),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_205),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_364),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_364),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_364),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_245),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_318),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_364),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_364),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_370),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_370),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_293),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_246),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_370),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_248),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_254),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_330),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_370),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_370),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_214),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_284),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_284),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_205),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_263),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_264),
.Y(n_469)
);

CKINVDCx14_ASAP7_75t_R g470 ( 
.A(n_335),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_299),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_299),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_324),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_324),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_244),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_378),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_266),
.Y(n_477)
);

BUFx2_ASAP7_75t_SL g478 ( 
.A(n_236),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_214),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_398),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_403),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_424),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_451),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_451),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_424),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_416),
.A2(n_239),
.B1(n_277),
.B2(n_218),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_434),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_403),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_404),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_404),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_451),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_434),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_478),
.B(n_236),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_440),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_405),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_405),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_406),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_389),
.B(n_244),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_406),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_451),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_395),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_399),
.Y(n_502)
);

INVx6_ASAP7_75t_L g503 ( 
.A(n_451),
.Y(n_503)
);

NAND2x1p5_ASAP7_75t_L g504 ( 
.A(n_385),
.B(n_310),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_432),
.B(n_261),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_400),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_440),
.B(n_249),
.Y(n_507)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_386),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_442),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_417),
.Y(n_510)
);

OA21x2_ASAP7_75t_L g511 ( 
.A1(n_385),
.A2(n_392),
.B(n_391),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_442),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_407),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_428),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_449),
.B(n_249),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_426),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_402),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_410),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_407),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_413),
.A2(n_309),
.B1(n_319),
.B2(n_286),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_418),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_394),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_408),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_449),
.B(n_272),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_422),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_425),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_408),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_412),
.A2(n_360),
.B1(n_342),
.B2(n_382),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_430),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_435),
.B(n_261),
.Y(n_530)
);

BUFx8_ASAP7_75t_L g531 ( 
.A(n_446),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_386),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_409),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_439),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_409),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_415),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_415),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_470),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_420),
.B(n_272),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_420),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_423),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_423),
.B(n_281),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_429),
.B(n_310),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_478),
.B(n_450),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_457),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_429),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_436),
.Y(n_547)
);

NAND2xp33_ASAP7_75t_R g548 ( 
.A(n_419),
.B(n_193),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_R g549 ( 
.A(n_477),
.B(n_269),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_436),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_459),
.B(n_308),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_437),
.Y(n_552)
);

NOR2x1_ASAP7_75t_L g553 ( 
.A(n_437),
.B(n_310),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_441),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_441),
.B(n_308),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_443),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_460),
.B(n_213),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_445),
.A2(n_280),
.B1(n_283),
.B2(n_366),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g559 ( 
.A(n_522),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_482),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_544),
.B(n_433),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_508),
.Y(n_562)
);

BUFx4f_ASAP7_75t_L g563 ( 
.A(n_511),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_482),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_508),
.Y(n_565)
);

AND2x6_ASAP7_75t_L g566 ( 
.A(n_505),
.B(n_213),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_505),
.B(n_475),
.Y(n_567)
);

AND2x6_ASAP7_75t_L g568 ( 
.A(n_530),
.B(n_223),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_531),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_485),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_491),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_531),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_485),
.Y(n_573)
);

BUFx10_ASAP7_75t_L g574 ( 
.A(n_501),
.Y(n_574)
);

AND3x1_ASAP7_75t_L g575 ( 
.A(n_493),
.B(n_431),
.C(n_421),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_508),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_491),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_508),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_487),
.Y(n_579)
);

AO21x2_ASAP7_75t_L g580 ( 
.A1(n_557),
.A2(n_199),
.B(n_197),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_487),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_481),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_481),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_506),
.B(n_461),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_551),
.B(n_468),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_488),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_491),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_498),
.B(n_469),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_492),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_492),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_494),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_488),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_489),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_494),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_533),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_489),
.Y(n_596)
);

INVx5_ASAP7_75t_L g597 ( 
.A(n_491),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g598 ( 
.A(n_531),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g599 ( 
.A(n_480),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_491),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_533),
.Y(n_601)
);

AOI21x1_ASAP7_75t_L g602 ( 
.A1(n_553),
.A2(n_392),
.B(n_391),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_490),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_490),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_491),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_484),
.Y(n_606)
);

INVx5_ASAP7_75t_L g607 ( 
.A(n_532),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_495),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_484),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_530),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_517),
.B(n_479),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_L g612 ( 
.A(n_504),
.B(n_318),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_555),
.B(n_388),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_495),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_539),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_531),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_496),
.Y(n_617)
);

INVx8_ASAP7_75t_L g618 ( 
.A(n_518),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_496),
.Y(n_619)
);

CKINVDCx16_ASAP7_75t_R g620 ( 
.A(n_548),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_521),
.B(n_438),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_525),
.B(n_411),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_526),
.B(n_387),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_555),
.B(n_465),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_497),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_534),
.B(n_411),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_497),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_545),
.B(n_414),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_511),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_535),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_535),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_539),
.B(n_444),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_555),
.B(n_507),
.Y(n_633)
);

CKINVDCx16_ASAP7_75t_R g634 ( 
.A(n_549),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_499),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_555),
.B(n_465),
.Y(n_636)
);

NAND3xp33_ASAP7_75t_L g637 ( 
.A(n_511),
.B(n_396),
.C(n_393),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_484),
.Y(n_638)
);

AND2x6_ASAP7_75t_L g639 ( 
.A(n_553),
.B(n_223),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_499),
.Y(n_640)
);

INVx4_ASAP7_75t_L g641 ( 
.A(n_511),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_513),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_513),
.Y(n_643)
);

OAI22xp33_ASAP7_75t_L g644 ( 
.A1(n_528),
.A2(n_390),
.B1(n_351),
.B2(n_338),
.Y(n_644)
);

OAI21xp33_ASAP7_75t_SL g645 ( 
.A1(n_519),
.A2(n_396),
.B(n_393),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_540),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_540),
.Y(n_647)
);

INVx8_ASAP7_75t_L g648 ( 
.A(n_543),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_484),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_538),
.B(n_411),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_484),
.Y(n_651)
);

OR2x6_ASAP7_75t_L g652 ( 
.A(n_504),
.B(n_242),
.Y(n_652)
);

INVxp33_ASAP7_75t_L g653 ( 
.A(n_520),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_519),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_541),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_504),
.A2(n_349),
.B1(n_341),
.B2(n_446),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_538),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_509),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_516),
.B(n_427),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_523),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_523),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_541),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_509),
.Y(n_663)
);

OAI22xp33_ASAP7_75t_L g664 ( 
.A1(n_516),
.A2(n_231),
.B1(n_247),
.B2(n_228),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_547),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_507),
.B(n_466),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_547),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_556),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_507),
.B(n_466),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_527),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_527),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_539),
.B(n_444),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_556),
.Y(n_673)
);

INVx4_ASAP7_75t_L g674 ( 
.A(n_509),
.Y(n_674)
);

INVxp33_ASAP7_75t_L g675 ( 
.A(n_520),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_539),
.B(n_447),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_536),
.Y(n_677)
);

INVx1_ASAP7_75t_SL g678 ( 
.A(n_502),
.Y(n_678)
);

AND3x2_ASAP7_75t_L g679 ( 
.A(n_542),
.B(n_282),
.C(n_242),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_532),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_536),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_542),
.B(n_447),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_537),
.Y(n_683)
);

NAND2xp33_ASAP7_75t_L g684 ( 
.A(n_509),
.B(n_318),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_529),
.B(n_467),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_SL g686 ( 
.A(n_486),
.B(n_368),
.Y(n_686)
);

AO22x2_ASAP7_75t_L g687 ( 
.A1(n_543),
.A2(n_349),
.B1(n_341),
.B2(n_346),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_532),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_542),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_510),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_529),
.B(n_464),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_507),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_537),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_532),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_542),
.B(n_456),
.Y(n_695)
);

INVxp67_ASAP7_75t_SL g696 ( 
.A(n_483),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_514),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_546),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_515),
.B(n_312),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_546),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_515),
.B(n_312),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_515),
.B(n_312),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_550),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_550),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_552),
.B(n_476),
.Y(n_705)
);

BUFx4f_ASAP7_75t_L g706 ( 
.A(n_509),
.Y(n_706)
);

AND3x2_ASAP7_75t_L g707 ( 
.A(n_515),
.B(n_282),
.C(n_210),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_552),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_554),
.Y(n_709)
);

INVx1_ASAP7_75t_SL g710 ( 
.A(n_558),
.Y(n_710)
);

A2O1A1Ixp33_ASAP7_75t_L g711 ( 
.A1(n_645),
.A2(n_322),
.B(n_316),
.C(n_287),
.Y(n_711)
);

NAND2xp33_ASAP7_75t_L g712 ( 
.A(n_566),
.B(n_270),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_563),
.B(n_318),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_666),
.B(n_524),
.Y(n_714)
);

BUFx8_ASAP7_75t_L g715 ( 
.A(n_657),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_559),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_588),
.B(n_524),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_610),
.B(n_524),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_610),
.B(n_193),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_700),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_680),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_680),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_567),
.A2(n_306),
.B1(n_334),
.B2(n_298),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_562),
.B(n_543),
.Y(n_724)
);

INVx4_ASAP7_75t_L g725 ( 
.A(n_648),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_562),
.B(n_554),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_563),
.B(n_629),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_565),
.B(n_483),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_685),
.B(n_585),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_613),
.A2(n_333),
.B1(n_331),
.B2(n_326),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_692),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_688),
.Y(n_732)
);

INVxp67_ASAP7_75t_L g733 ( 
.A(n_691),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_666),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_565),
.B(n_483),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_576),
.B(n_483),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_669),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_576),
.B(n_500),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_563),
.B(n_318),
.Y(n_739)
);

NAND2xp33_ASAP7_75t_L g740 ( 
.A(n_566),
.B(n_304),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_669),
.Y(n_741)
);

NAND2xp33_ASAP7_75t_L g742 ( 
.A(n_566),
.B(n_311),
.Y(n_742)
);

A2O1A1Ixp33_ASAP7_75t_L g743 ( 
.A1(n_645),
.A2(n_268),
.B(n_262),
.C(n_258),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_578),
.B(n_500),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_578),
.B(n_500),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_641),
.B(n_195),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_629),
.B(n_363),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_633),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_700),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_688),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_633),
.B(n_500),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_629),
.B(n_363),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_615),
.B(n_509),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_615),
.B(n_512),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_694),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_689),
.B(n_512),
.Y(n_756)
);

INVx8_ASAP7_75t_L g757 ( 
.A(n_618),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_632),
.Y(n_758)
);

HB1xp67_ASAP7_75t_L g759 ( 
.A(n_613),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_689),
.B(n_512),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_695),
.A2(n_314),
.B1(n_315),
.B2(n_317),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_641),
.B(n_195),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_641),
.B(n_363),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_641),
.B(n_200),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_561),
.B(n_200),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_694),
.Y(n_766)
);

OR2x2_ASAP7_75t_L g767 ( 
.A(n_620),
.B(n_558),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_582),
.B(n_512),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_672),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_637),
.B(n_363),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_637),
.B(n_363),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_676),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_560),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_682),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_582),
.B(n_512),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_559),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_648),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_620),
.B(n_275),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_652),
.A2(n_257),
.B1(n_295),
.B2(n_289),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_583),
.B(n_512),
.Y(n_780)
);

OAI22x1_ASAP7_75t_SL g781 ( 
.A1(n_710),
.A2(n_352),
.B1(n_342),
.B2(n_344),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_583),
.B(n_209),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_564),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_705),
.B(n_204),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_703),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_564),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_586),
.B(n_212),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_703),
.B(n_380),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_570),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_570),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_653),
.B(n_204),
.Y(n_791)
);

NAND2xp33_ASAP7_75t_SL g792 ( 
.A(n_675),
.B(n_657),
.Y(n_792)
);

INVxp67_ASAP7_75t_SL g793 ( 
.A(n_606),
.Y(n_793)
);

INVxp33_ASAP7_75t_L g794 ( 
.A(n_623),
.Y(n_794)
);

NOR2xp67_ASAP7_75t_L g795 ( 
.A(n_628),
.B(n_313),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_592),
.B(n_221),
.Y(n_796)
);

OAI22xp33_ASAP7_75t_L g797 ( 
.A1(n_686),
.A2(n_339),
.B1(n_362),
.B2(n_369),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_566),
.A2(n_323),
.B1(n_216),
.B2(n_211),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_566),
.A2(n_216),
.B1(n_276),
.B2(n_290),
.Y(n_799)
);

NOR2xp67_ASAP7_75t_L g800 ( 
.A(n_622),
.B(n_207),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_704),
.B(n_380),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_593),
.B(n_224),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_573),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_624),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_593),
.B(n_233),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_704),
.B(n_380),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_596),
.B(n_603),
.Y(n_807)
);

INVxp67_ASAP7_75t_L g808 ( 
.A(n_575),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_596),
.B(n_237),
.Y(n_809)
);

INVxp67_ASAP7_75t_L g810 ( 
.A(n_575),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_603),
.B(n_251),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_604),
.B(n_256),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_618),
.Y(n_813)
);

OAI22xp33_ASAP7_75t_L g814 ( 
.A1(n_686),
.A2(n_371),
.B1(n_255),
.B2(n_241),
.Y(n_814)
);

NAND2xp33_ASAP7_75t_L g815 ( 
.A(n_566),
.B(n_380),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_604),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_624),
.B(n_471),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_659),
.B(n_207),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_664),
.B(n_208),
.Y(n_819)
);

NOR3xp33_ASAP7_75t_L g820 ( 
.A(n_644),
.B(n_486),
.C(n_252),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_SL g821 ( 
.A(n_634),
.B(n_208),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_708),
.B(n_380),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_573),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_608),
.B(n_614),
.Y(n_824)
);

A2O1A1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_636),
.A2(n_340),
.B(n_343),
.C(n_353),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_708),
.B(n_265),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_SL g827 ( 
.A(n_634),
.B(n_569),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_608),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_579),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_614),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_579),
.Y(n_831)
);

AO22x2_ASAP7_75t_L g832 ( 
.A1(n_687),
.A2(n_196),
.B1(n_206),
.B2(n_215),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_617),
.B(n_271),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_636),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_648),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_617),
.B(n_273),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_619),
.B(n_625),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_619),
.B(n_274),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_625),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_581),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_627),
.B(n_279),
.Y(n_841)
);

INVx4_ASAP7_75t_L g842 ( 
.A(n_648),
.Y(n_842)
);

A2O1A1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_656),
.A2(n_232),
.B(n_397),
.C(n_401),
.Y(n_843)
);

BUFx6f_ASAP7_75t_SL g844 ( 
.A(n_574),
.Y(n_844)
);

HB1xp67_ASAP7_75t_L g845 ( 
.A(n_687),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_574),
.B(n_275),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_581),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_627),
.B(n_635),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_589),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_L g850 ( 
.A(n_566),
.B(n_211),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_568),
.A2(n_345),
.B1(n_276),
.B2(n_290),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_590),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_687),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_635),
.B(n_285),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_R g855 ( 
.A(n_697),
.B(n_618),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_696),
.A2(n_397),
.B(n_401),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_640),
.B(n_301),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_574),
.B(n_621),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_640),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_699),
.B(n_220),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_652),
.A2(n_354),
.B1(n_355),
.B2(n_365),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_642),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_642),
.A2(n_328),
.B(n_373),
.C(n_307),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_643),
.B(n_320),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_643),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_590),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_654),
.B(n_327),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_654),
.B(n_332),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_660),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_591),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_648),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_661),
.B(n_384),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_661),
.B(n_448),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_748),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_855),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_727),
.B(n_670),
.Y(n_876)
);

INVx3_ASAP7_75t_L g877 ( 
.A(n_714),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_777),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_794),
.B(n_584),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_720),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_720),
.Y(n_881)
);

NAND3xp33_ASAP7_75t_SL g882 ( 
.A(n_784),
.B(n_626),
.C(n_701),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_749),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_727),
.B(n_709),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_749),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_829),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_845),
.A2(n_687),
.B1(n_568),
.B2(n_580),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_785),
.Y(n_888)
);

BUFx8_ASAP7_75t_L g889 ( 
.A(n_844),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_785),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_714),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_729),
.B(n_580),
.Y(n_892)
);

NAND2x1p5_ASAP7_75t_L g893 ( 
.A(n_777),
.B(n_670),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_717),
.A2(n_652),
.B(n_706),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_729),
.A2(n_652),
.B1(n_618),
.B2(n_709),
.Y(n_895)
);

OR2x2_ASAP7_75t_L g896 ( 
.A(n_716),
.B(n_599),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_733),
.B(n_759),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_784),
.A2(n_568),
.B1(n_652),
.B2(n_580),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_870),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_816),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_758),
.B(n_568),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_763),
.A2(n_568),
.B(n_602),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_759),
.B(n_791),
.Y(n_903)
);

AO21x1_ASAP7_75t_L g904 ( 
.A1(n_713),
.A2(n_612),
.B(n_671),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_828),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_830),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_831),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_769),
.B(n_568),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_813),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_791),
.B(n_611),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_831),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_772),
.B(n_677),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_840),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_804),
.A2(n_702),
.B1(n_693),
.B2(n_681),
.Y(n_914)
);

BUFx12f_ASAP7_75t_L g915 ( 
.A(n_715),
.Y(n_915)
);

AOI22xp33_ASAP7_75t_L g916 ( 
.A1(n_845),
.A2(n_639),
.B1(n_698),
.B2(n_693),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_774),
.B(n_677),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_839),
.B(n_681),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_808),
.B(n_810),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_853),
.A2(n_639),
.B1(n_698),
.B2(n_683),
.Y(n_920)
);

AND2x6_ASAP7_75t_SL g921 ( 
.A(n_819),
.B(n_697),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_859),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_815),
.A2(n_706),
.B(n_674),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_862),
.B(n_683),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_840),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_777),
.B(n_618),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_865),
.B(n_649),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_819),
.A2(n_598),
.B(n_572),
.C(n_616),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_869),
.B(n_649),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_773),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_778),
.B(n_569),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_777),
.B(n_572),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_846),
.B(n_598),
.Y(n_933)
);

INVx4_ASAP7_75t_L g934 ( 
.A(n_757),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_L g935 ( 
.A1(n_853),
.A2(n_639),
.B1(n_630),
.B2(n_673),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_807),
.B(n_651),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_824),
.B(n_651),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_731),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_835),
.B(n_871),
.Y(n_939)
);

NOR2xp67_ASAP7_75t_L g940 ( 
.A(n_761),
.B(n_650),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_776),
.B(n_616),
.Y(n_941)
);

OR2x6_ASAP7_75t_L g942 ( 
.A(n_757),
.B(n_678),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_837),
.B(n_848),
.Y(n_943)
);

OR2x6_ASAP7_75t_L g944 ( 
.A(n_757),
.B(n_690),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_834),
.B(n_651),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_835),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_718),
.B(n_571),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_719),
.B(n_571),
.Y(n_948)
);

INVx2_ASAP7_75t_SL g949 ( 
.A(n_817),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_734),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_783),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_813),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_737),
.A2(n_639),
.B1(n_658),
.B2(n_663),
.Y(n_953)
);

INVx2_ASAP7_75t_SL g954 ( 
.A(n_817),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_786),
.Y(n_955)
);

NOR2xp67_ASAP7_75t_L g956 ( 
.A(n_719),
.B(n_595),
.Y(n_956)
);

BUFx2_ASAP7_75t_L g957 ( 
.A(n_715),
.Y(n_957)
);

NOR3xp33_ASAP7_75t_SL g958 ( 
.A(n_797),
.B(n_814),
.C(n_792),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_767),
.Y(n_959)
);

AOI22xp5_ASAP7_75t_L g960 ( 
.A1(n_741),
.A2(n_639),
.B1(n_658),
.B2(n_663),
.Y(n_960)
);

BUFx12f_ASAP7_75t_L g961 ( 
.A(n_858),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_835),
.B(n_658),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_855),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_751),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_835),
.B(n_663),
.Y(n_965)
);

AND2x4_ASAP7_75t_SL g966 ( 
.A(n_871),
.B(n_350),
.Y(n_966)
);

BUFx10_ASAP7_75t_L g967 ( 
.A(n_844),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_789),
.Y(n_968)
);

BUFx2_ASAP7_75t_L g969 ( 
.A(n_832),
.Y(n_969)
);

AOI221xp5_ASAP7_75t_SL g970 ( 
.A1(n_797),
.A2(n_474),
.B1(n_473),
.B2(n_472),
.C(n_471),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_790),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_746),
.B(n_762),
.Y(n_972)
);

NOR2x1_ASAP7_75t_R g973 ( 
.A(n_841),
.B(n_344),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_821),
.B(n_250),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_803),
.Y(n_975)
);

INVx2_ASAP7_75t_SL g976 ( 
.A(n_841),
.Y(n_976)
);

OR2x2_ASAP7_75t_L g977 ( 
.A(n_765),
.B(n_347),
.Y(n_977)
);

BUFx2_ASAP7_75t_L g978 ( 
.A(n_832),
.Y(n_978)
);

AOI21x1_ASAP7_75t_L g979 ( 
.A1(n_713),
.A2(n_667),
.B(n_646),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_871),
.B(n_707),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_823),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_847),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_L g983 ( 
.A1(n_832),
.A2(n_639),
.B1(n_662),
.B2(n_655),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_871),
.B(n_706),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_781),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_764),
.B(n_577),
.Y(n_986)
);

CKINVDCx6p67_ASAP7_75t_R g987 ( 
.A(n_864),
.Y(n_987)
);

INVx2_ASAP7_75t_SL g988 ( 
.A(n_782),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_849),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_725),
.B(n_606),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_725),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_764),
.A2(n_639),
.B1(n_647),
.B2(n_646),
.Y(n_992)
);

AOI22xp33_ASAP7_75t_L g993 ( 
.A1(n_814),
.A2(n_630),
.B1(n_601),
.B2(n_595),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_795),
.B(n_587),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_852),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_866),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_747),
.B(n_587),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_842),
.B(n_606),
.Y(n_998)
);

BUFx3_ASAP7_75t_L g999 ( 
.A(n_873),
.Y(n_999)
);

AOI22xp33_ASAP7_75t_SL g1000 ( 
.A1(n_765),
.A2(n_350),
.B1(n_347),
.B2(n_352),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_721),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_768),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_775),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_780),
.Y(n_1004)
);

OR2x6_ASAP7_75t_L g1005 ( 
.A(n_825),
.B(n_472),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_747),
.A2(n_655),
.B(n_601),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_722),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_732),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_750),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_752),
.B(n_587),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_860),
.B(n_253),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_842),
.B(n_606),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_755),
.Y(n_1013)
);

NAND3xp33_ASAP7_75t_L g1014 ( 
.A(n_820),
.B(n_291),
.C(n_292),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_766),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_818),
.B(n_350),
.Y(n_1016)
);

NAND2x1_ASAP7_75t_L g1017 ( 
.A(n_753),
.B(n_674),
.Y(n_1017)
);

BUFx12f_ASAP7_75t_L g1018 ( 
.A(n_827),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_724),
.A2(n_674),
.B(n_606),
.Y(n_1019)
);

INVx5_ASAP7_75t_L g1020 ( 
.A(n_739),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_787),
.B(n_600),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_796),
.B(n_600),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_802),
.B(n_605),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_860),
.A2(n_668),
.B1(n_631),
.B2(n_662),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_711),
.A2(n_360),
.B(n_361),
.C(n_356),
.Y(n_1025)
);

INVx2_ASAP7_75t_SL g1026 ( 
.A(n_805),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_799),
.B(n_609),
.Y(n_1027)
);

AND3x1_ASAP7_75t_L g1028 ( 
.A(n_818),
.B(n_825),
.C(n_743),
.Y(n_1028)
);

NAND2xp33_ASAP7_75t_SL g1029 ( 
.A(n_739),
.B(n_220),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_770),
.A2(n_376),
.B1(n_379),
.B2(n_337),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_728),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_735),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_736),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_851),
.B(n_609),
.Y(n_1034)
);

OR2x2_ASAP7_75t_L g1035 ( 
.A(n_723),
.B(n_356),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_730),
.B(n_296),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_800),
.B(n_843),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_809),
.B(n_605),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_798),
.B(n_609),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_811),
.B(n_605),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_738),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_770),
.A2(n_379),
.B1(n_383),
.B2(n_337),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_754),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_744),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_812),
.B(n_361),
.Y(n_1045)
);

INVx1_ASAP7_75t_SL g1046 ( 
.A(n_833),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_843),
.B(n_836),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_711),
.B(n_679),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_745),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_838),
.B(n_631),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_943),
.A2(n_740),
.B(n_742),
.Y(n_1051)
);

OR2x6_ASAP7_75t_L g1052 ( 
.A(n_942),
.B(n_743),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_R g1053 ( 
.A(n_875),
.B(n_850),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_SL g1054 ( 
.A1(n_1011),
.A2(n_712),
.B(n_868),
.C(n_867),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_923),
.A2(n_793),
.B(n_756),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_903),
.B(n_854),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_910),
.B(n_771),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_910),
.B(n_903),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_1011),
.A2(n_857),
.B(n_872),
.C(n_861),
.Y(n_1059)
);

O2A1O1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_958),
.A2(n_972),
.B(n_977),
.C(n_882),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_961),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_964),
.B(n_726),
.Y(n_1062)
);

BUFx2_ASAP7_75t_L g1063 ( 
.A(n_896),
.Y(n_1063)
);

O2A1O1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_958),
.A2(n_826),
.B(n_863),
.C(n_779),
.Y(n_1064)
);

NAND2xp33_ASAP7_75t_SL g1065 ( 
.A(n_991),
.B(n_771),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_892),
.B(n_856),
.Y(n_1066)
);

INVx5_ASAP7_75t_L g1067 ( 
.A(n_878),
.Y(n_1067)
);

O2A1O1Ixp33_ASAP7_75t_SL g1068 ( 
.A1(n_876),
.A2(n_863),
.B(n_822),
.C(n_806),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_1036),
.A2(n_826),
.B1(n_760),
.B2(n_806),
.Y(n_1069)
);

BUFx12f_ASAP7_75t_L g1070 ( 
.A(n_967),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_912),
.B(n_647),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_886),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_SL g1073 ( 
.A(n_934),
.B(n_345),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_882),
.A2(n_822),
.B(n_801),
.C(n_788),
.Y(n_1074)
);

INVx2_ASAP7_75t_SL g1075 ( 
.A(n_959),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_917),
.B(n_665),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_1036),
.A2(n_801),
.B(n_788),
.C(n_665),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_1018),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1002),
.B(n_667),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_899),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_900),
.Y(n_1081)
);

NOR2xp67_ASAP7_75t_SL g1082 ( 
.A(n_991),
.B(n_348),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_905),
.Y(n_1083)
);

AOI22x1_ASAP7_75t_L g1084 ( 
.A1(n_894),
.A2(n_673),
.B1(n_668),
.B2(n_591),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_916),
.A2(n_374),
.B1(n_381),
.B2(n_382),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_1001),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_878),
.Y(n_1087)
);

BUFx3_ASAP7_75t_L g1088 ( 
.A(n_915),
.Y(n_1088)
);

O2A1O1Ixp5_ASAP7_75t_L g1089 ( 
.A1(n_904),
.A2(n_594),
.B(n_448),
.C(n_452),
.Y(n_1089)
);

AOI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_940),
.A2(n_367),
.B1(n_376),
.B2(n_383),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_906),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_1046),
.B(n_348),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_922),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_1000),
.A2(n_367),
.B1(n_594),
.B2(n_452),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_880),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_879),
.B(n_297),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_879),
.B(n_303),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_901),
.A2(n_638),
.B(n_609),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1001),
.Y(n_1099)
);

AOI21x1_ASAP7_75t_L g1100 ( 
.A1(n_876),
.A2(n_453),
.B(n_454),
.Y(n_1100)
);

OAI21xp33_ASAP7_75t_L g1101 ( 
.A1(n_1000),
.A2(n_381),
.B(n_377),
.Y(n_1101)
);

NOR3xp33_ASAP7_75t_L g1102 ( 
.A(n_931),
.B(n_305),
.C(n_336),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_908),
.A2(n_638),
.B(n_684),
.Y(n_1103)
);

NOR3xp33_ASAP7_75t_SL g1104 ( 
.A(n_985),
.B(n_374),
.C(n_377),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_SL g1105 ( 
.A1(n_919),
.A2(n_974),
.B(n_895),
.C(n_902),
.Y(n_1105)
);

A2O1A1Ixp33_ASAP7_75t_SL g1106 ( 
.A1(n_919),
.A2(n_463),
.B(n_454),
.C(n_455),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1019),
.A2(n_638),
.B(n_597),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_974),
.A2(n_321),
.B(n_329),
.C(n_474),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_897),
.B(n_607),
.Y(n_1109)
);

OR2x6_ASAP7_75t_SL g1110 ( 
.A(n_963),
.B(n_473),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_907),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_969),
.A2(n_462),
.B1(n_455),
.B2(n_458),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_949),
.B(n_126),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_988),
.B(n_0),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_986),
.A2(n_607),
.B(n_597),
.Y(n_1115)
);

OR2x6_ASAP7_75t_SL g1116 ( 
.A(n_1014),
.B(n_463),
.Y(n_1116)
);

CKINVDCx8_ASAP7_75t_R g1117 ( 
.A(n_921),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_878),
.Y(n_1118)
);

NOR3xp33_ASAP7_75t_SL g1119 ( 
.A(n_928),
.B(n_2),
.C(n_3),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_954),
.B(n_119),
.Y(n_1120)
);

AOI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_877),
.A2(n_607),
.B1(n_503),
.B2(n_597),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_1026),
.B(n_4),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_933),
.B(n_607),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1039),
.A2(n_597),
.B(n_503),
.Y(n_1124)
);

NAND2x1p5_ASAP7_75t_L g1125 ( 
.A(n_991),
.B(n_111),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_889),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1016),
.B(n_9),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_881),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1039),
.A2(n_503),
.B(n_188),
.Y(n_1129)
);

CKINVDCx20_ASAP7_75t_R g1130 ( 
.A(n_889),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_1035),
.B(n_15),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_941),
.B(n_15),
.Y(n_1132)
);

OAI21xp33_ASAP7_75t_L g1133 ( 
.A1(n_1045),
.A2(n_16),
.B(n_19),
.Y(n_1133)
);

CKINVDCx14_ASAP7_75t_R g1134 ( 
.A(n_957),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_948),
.A2(n_503),
.B(n_166),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_987),
.B(n_20),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_907),
.Y(n_1137)
);

INVx6_ASAP7_75t_L g1138 ( 
.A(n_967),
.Y(n_1138)
);

A2O1A1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_976),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_1139)
);

CKINVDCx20_ASAP7_75t_R g1140 ( 
.A(n_942),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_883),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_916),
.A2(n_920),
.B1(n_935),
.B2(n_1020),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_950),
.B(n_24),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_874),
.B(n_25),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_891),
.B(n_106),
.Y(n_1145)
);

AOI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_1037),
.A2(n_158),
.B1(n_151),
.B2(n_148),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1027),
.A2(n_95),
.B(n_142),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1003),
.B(n_1004),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_942),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_980),
.B(n_93),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_885),
.Y(n_1151)
);

O2A1O1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1025),
.A2(n_29),
.B(n_30),
.C(n_32),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_888),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1027),
.A2(n_1034),
.B(n_937),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_890),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1031),
.B(n_125),
.Y(n_1156)
);

OA22x2_ASAP7_75t_L g1157 ( 
.A1(n_978),
.A2(n_29),
.B1(n_33),
.B2(n_35),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_SL g1158 ( 
.A1(n_945),
.A2(n_898),
.B(n_1043),
.C(n_1006),
.Y(n_1158)
);

AO32x2_ASAP7_75t_L g1159 ( 
.A1(n_1030),
.A2(n_35),
.A3(n_36),
.B1(n_37),
.B2(n_42),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_SL g1160 ( 
.A1(n_1028),
.A2(n_36),
.B1(n_45),
.B2(n_46),
.Y(n_1160)
);

OR2x2_ASAP7_75t_L g1161 ( 
.A(n_944),
.B(n_47),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1032),
.B(n_65),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_878),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_981),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1034),
.A2(n_109),
.B(n_105),
.Y(n_1165)
);

NAND3xp33_ASAP7_75t_L g1166 ( 
.A(n_914),
.B(n_47),
.C(n_50),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_973),
.B(n_50),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1033),
.B(n_120),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1037),
.B(n_91),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_984),
.A2(n_82),
.B(n_74),
.Y(n_1170)
);

OAI22x1_ASAP7_75t_L g1171 ( 
.A1(n_1048),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_1171)
);

AND2x2_ASAP7_75t_SL g1172 ( 
.A(n_966),
.B(n_55),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_991),
.B(n_918),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_920),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_981),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_911),
.Y(n_1176)
);

INVx4_ASAP7_75t_L g1177 ( 
.A(n_946),
.Y(n_1177)
);

NOR2x1p5_ASAP7_75t_L g1178 ( 
.A(n_909),
.B(n_68),
.Y(n_1178)
);

AND2x2_ASAP7_75t_SL g1179 ( 
.A(n_966),
.B(n_60),
.Y(n_1179)
);

AOI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1029),
.A2(n_62),
.B1(n_956),
.B2(n_932),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_924),
.B(n_946),
.Y(n_1181)
);

INVx4_ASAP7_75t_L g1182 ( 
.A(n_946),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_984),
.A2(n_947),
.B(n_994),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_999),
.B(n_938),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_946),
.B(n_1020),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_944),
.Y(n_1186)
);

NOR2x1_ASAP7_75t_R g1187 ( 
.A(n_980),
.B(n_909),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_999),
.B(n_928),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_944),
.Y(n_1189)
);

OR2x2_ASAP7_75t_L g1190 ( 
.A(n_968),
.B(n_971),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1047),
.A2(n_1049),
.B(n_1044),
.C(n_1041),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_982),
.Y(n_1192)
);

NAND3xp33_ASAP7_75t_SL g1193 ( 
.A(n_1025),
.B(n_932),
.C(n_1042),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_913),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_989),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_1048),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_936),
.A2(n_884),
.B(n_1020),
.Y(n_1197)
);

AND2x6_ASAP7_75t_SL g1198 ( 
.A(n_1005),
.B(n_945),
.Y(n_1198)
);

INVx2_ASAP7_75t_SL g1199 ( 
.A(n_930),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1051),
.A2(n_1020),
.B(n_1012),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1058),
.B(n_1043),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1057),
.B(n_1050),
.Y(n_1202)
);

O2A1O1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1131),
.A2(n_884),
.B(n_926),
.C(n_1005),
.Y(n_1203)
);

OA21x2_ASAP7_75t_L g1204 ( 
.A1(n_1154),
.A2(n_970),
.B(n_992),
.Y(n_1204)
);

NAND3xp33_ASAP7_75t_SL g1205 ( 
.A(n_1096),
.B(n_887),
.C(n_1024),
.Y(n_1205)
);

AOI21xp33_ASAP7_75t_L g1206 ( 
.A1(n_1060),
.A2(n_887),
.B(n_1040),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1066),
.A2(n_990),
.B(n_1012),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1062),
.B(n_975),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1142),
.A2(n_1148),
.B1(n_1160),
.B2(n_1062),
.Y(n_1209)
);

O2A1O1Ixp5_ASAP7_75t_L g1210 ( 
.A1(n_1065),
.A2(n_990),
.B(n_998),
.C(n_939),
.Y(n_1210)
);

NAND3xp33_ASAP7_75t_L g1211 ( 
.A(n_1097),
.B(n_983),
.C(n_1005),
.Y(n_1211)
);

AO22x2_ASAP7_75t_L g1212 ( 
.A1(n_1174),
.A2(n_926),
.B1(n_939),
.B2(n_998),
.Y(n_1212)
);

NOR2xp67_ASAP7_75t_L g1213 ( 
.A(n_1075),
.B(n_996),
.Y(n_1213)
);

AOI221x1_ASAP7_75t_L g1214 ( 
.A1(n_1166),
.A2(n_1038),
.B1(n_1022),
.B2(n_1023),
.C(n_1021),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_SL g1215 ( 
.A1(n_1142),
.A2(n_934),
.B(n_952),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1056),
.B(n_935),
.Y(n_1216)
);

BUFx10_ASAP7_75t_L g1217 ( 
.A(n_1138),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1055),
.A2(n_893),
.B(n_1017),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_1063),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1098),
.A2(n_962),
.B(n_965),
.Y(n_1220)
);

AOI21x1_ASAP7_75t_SL g1221 ( 
.A1(n_1127),
.A2(n_997),
.B(n_1010),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1183),
.A2(n_927),
.B(n_929),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1184),
.B(n_995),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1066),
.A2(n_960),
.B(n_953),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1107),
.A2(n_1124),
.B(n_1154),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1196),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1087),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1188),
.B(n_955),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1064),
.A2(n_983),
.B(n_1015),
.C(n_1008),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1103),
.A2(n_1100),
.B(n_1115),
.Y(n_1230)
);

INVx2_ASAP7_75t_SL g1231 ( 
.A(n_1138),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1081),
.B(n_1083),
.Y(n_1232)
);

AO31x2_ASAP7_75t_L g1233 ( 
.A1(n_1191),
.A2(n_1007),
.A3(n_1009),
.B(n_1013),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1089),
.A2(n_993),
.B(n_951),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1092),
.B(n_925),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1091),
.B(n_1093),
.Y(n_1236)
);

OAI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1059),
.A2(n_993),
.B(n_952),
.Y(n_1237)
);

BUFx2_ASAP7_75t_R g1238 ( 
.A(n_1088),
.Y(n_1238)
);

OA21x2_ASAP7_75t_L g1239 ( 
.A1(n_1197),
.A2(n_1135),
.B(n_1077),
.Y(n_1239)
);

AOI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1133),
.A2(n_1174),
.B1(n_1167),
.B2(n_1114),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1071),
.B(n_1076),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1197),
.A2(n_1129),
.B(n_1147),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1071),
.B(n_1076),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1079),
.B(n_1095),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1079),
.B(n_1128),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1054),
.A2(n_1158),
.B(n_1105),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1173),
.A2(n_1156),
.B(n_1162),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1156),
.A2(n_1162),
.B(n_1168),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1151),
.B(n_1155),
.Y(n_1249)
);

A2O1A1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1180),
.A2(n_1165),
.B(n_1147),
.C(n_1193),
.Y(n_1250)
);

INVx2_ASAP7_75t_SL g1251 ( 
.A(n_1186),
.Y(n_1251)
);

INVx6_ASAP7_75t_SL g1252 ( 
.A(n_1150),
.Y(n_1252)
);

AO21x1_ASAP7_75t_L g1253 ( 
.A1(n_1165),
.A2(n_1135),
.B(n_1168),
.Y(n_1253)
);

INVx4_ASAP7_75t_L g1254 ( 
.A(n_1067),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1069),
.A2(n_1185),
.B(n_1074),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1181),
.A2(n_1170),
.B(n_1109),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_R g1257 ( 
.A(n_1134),
.B(n_1140),
.Y(n_1257)
);

AND2x2_ASAP7_75t_SL g1258 ( 
.A(n_1172),
.B(n_1179),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_1130),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1068),
.A2(n_1067),
.B(n_1169),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1122),
.A2(n_1102),
.B1(n_1132),
.B2(n_1101),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1143),
.B(n_1144),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1199),
.B(n_1192),
.Y(n_1263)
);

INVx6_ASAP7_75t_L g1264 ( 
.A(n_1070),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1111),
.A2(n_1137),
.B(n_1141),
.Y(n_1265)
);

NOR2xp67_ASAP7_75t_SL g1266 ( 
.A(n_1067),
.B(n_1117),
.Y(n_1266)
);

OA21x2_ASAP7_75t_L g1267 ( 
.A1(n_1123),
.A2(n_1153),
.B(n_1086),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1099),
.A2(n_1125),
.B(n_1080),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1150),
.B(n_1189),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1190),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1108),
.A2(n_1152),
.B(n_1094),
.Y(n_1271)
);

O2A1O1Ixp5_ASAP7_75t_L g1272 ( 
.A1(n_1082),
.A2(n_1106),
.B(n_1139),
.C(n_1195),
.Y(n_1272)
);

BUFx8_ASAP7_75t_L g1273 ( 
.A(n_1078),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1145),
.B(n_1116),
.Y(n_1274)
);

OR2x2_ASAP7_75t_L g1275 ( 
.A(n_1164),
.B(n_1175),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1145),
.B(n_1120),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_1090),
.B(n_1113),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_SL g1278 ( 
.A(n_1187),
.B(n_1073),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1113),
.B(n_1120),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1125),
.A2(n_1072),
.B(n_1121),
.Y(n_1280)
);

AO31x2_ASAP7_75t_L g1281 ( 
.A1(n_1171),
.A2(n_1176),
.A3(n_1194),
.B(n_1085),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1157),
.Y(n_1282)
);

INVx2_ASAP7_75t_SL g1283 ( 
.A(n_1061),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1104),
.B(n_1136),
.Y(n_1284)
);

INVx2_ASAP7_75t_SL g1285 ( 
.A(n_1149),
.Y(n_1285)
);

AO21x2_ASAP7_75t_L g1286 ( 
.A1(n_1146),
.A2(n_1119),
.B(n_1053),
.Y(n_1286)
);

OAI21xp5_ASAP7_75t_SL g1287 ( 
.A1(n_1085),
.A2(n_1161),
.B(n_1112),
.Y(n_1287)
);

OA21x2_ASAP7_75t_L g1288 ( 
.A1(n_1159),
.A2(n_1052),
.B(n_1198),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1052),
.B(n_1178),
.Y(n_1289)
);

OAI21xp33_ASAP7_75t_SL g1290 ( 
.A1(n_1157),
.A2(n_1052),
.B(n_1182),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1177),
.A2(n_1182),
.B(n_1159),
.Y(n_1291)
);

OR2x6_ASAP7_75t_L g1292 ( 
.A(n_1177),
.B(n_1087),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1087),
.A2(n_1163),
.B(n_1118),
.Y(n_1293)
);

CKINVDCx6p67_ASAP7_75t_R g1294 ( 
.A(n_1110),
.Y(n_1294)
);

OA21x2_ASAP7_75t_L g1295 ( 
.A1(n_1159),
.A2(n_1118),
.B(n_1163),
.Y(n_1295)
);

OR2x2_ASAP7_75t_L g1296 ( 
.A(n_1063),
.B(n_599),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1084),
.A2(n_1055),
.B(n_979),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1058),
.A2(n_1142),
.B1(n_1057),
.B2(n_958),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1058),
.B(n_903),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1084),
.A2(n_1055),
.B(n_979),
.Y(n_1300)
);

AOI221x1_ASAP7_75t_L g1301 ( 
.A1(n_1058),
.A2(n_972),
.B1(n_1011),
.B2(n_1057),
.C(n_1160),
.Y(n_1301)
);

NOR2x1_ASAP7_75t_L g1302 ( 
.A(n_1177),
.B(n_813),
.Y(n_1302)
);

A2O1A1Ixp33_ASAP7_75t_L g1303 ( 
.A1(n_1057),
.A2(n_1060),
.B(n_910),
.C(n_1058),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1063),
.B(n_599),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1058),
.B(n_903),
.Y(n_1305)
);

NOR2xp67_ASAP7_75t_L g1306 ( 
.A(n_1075),
.B(n_716),
.Y(n_1306)
);

AOI211x1_ASAP7_75t_L g1307 ( 
.A1(n_1174),
.A2(n_797),
.B(n_814),
.C(n_1101),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1058),
.B(n_903),
.Y(n_1308)
);

BUFx3_ASAP7_75t_L g1309 ( 
.A(n_1138),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_SL g1310 ( 
.A1(n_1142),
.A2(n_991),
.B(n_842),
.Y(n_1310)
);

OAI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1057),
.A2(n_972),
.B(n_1154),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1058),
.B(n_903),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1058),
.B(n_903),
.Y(n_1313)
);

INVx5_ASAP7_75t_L g1314 ( 
.A(n_1087),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1063),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1084),
.A2(n_1055),
.B(n_979),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1051),
.A2(n_1066),
.B(n_972),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1051),
.A2(n_1066),
.B(n_972),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1051),
.A2(n_1066),
.B(n_972),
.Y(n_1319)
);

AOI21xp33_ASAP7_75t_L g1320 ( 
.A1(n_1060),
.A2(n_1058),
.B(n_1057),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1063),
.B(n_599),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1051),
.A2(n_1066),
.B(n_972),
.Y(n_1322)
);

O2A1O1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1058),
.A2(n_1011),
.B(n_910),
.C(n_784),
.Y(n_1323)
);

OAI22x1_ASAP7_75t_L g1324 ( 
.A1(n_1058),
.A2(n_1131),
.B1(n_910),
.B2(n_1180),
.Y(n_1324)
);

INVx1_ASAP7_75t_SL g1325 ( 
.A(n_1063),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1051),
.A2(n_1066),
.B(n_972),
.Y(n_1326)
);

AO31x2_ASAP7_75t_L g1327 ( 
.A1(n_1154),
.A2(n_904),
.A3(n_1191),
.B(n_972),
.Y(n_1327)
);

BUFx2_ASAP7_75t_R g1328 ( 
.A(n_1126),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_SL g1329 ( 
.A(n_1058),
.B(n_620),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_1063),
.Y(n_1330)
);

BUFx10_ASAP7_75t_L g1331 ( 
.A(n_1138),
.Y(n_1331)
);

INVx1_ASAP7_75t_SL g1332 ( 
.A(n_1063),
.Y(n_1332)
);

AO21x2_ASAP7_75t_L g1333 ( 
.A1(n_1154),
.A2(n_972),
.B(n_1051),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1196),
.B(n_1150),
.Y(n_1334)
);

NAND2xp33_ASAP7_75t_L g1335 ( 
.A(n_1053),
.B(n_757),
.Y(n_1335)
);

INVx2_ASAP7_75t_SL g1336 ( 
.A(n_1063),
.Y(n_1336)
);

INVx4_ASAP7_75t_L g1337 ( 
.A(n_1067),
.Y(n_1337)
);

OAI22x1_ASAP7_75t_L g1338 ( 
.A1(n_1058),
.A2(n_1131),
.B1(n_910),
.B2(n_1180),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1058),
.B(n_903),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1058),
.B(n_903),
.Y(n_1340)
);

BUFx6f_ASAP7_75t_L g1341 ( 
.A(n_1087),
.Y(n_1341)
);

AND2x6_ASAP7_75t_L g1342 ( 
.A(n_1150),
.B(n_1145),
.Y(n_1342)
);

BUFx2_ASAP7_75t_SL g1343 ( 
.A(n_1061),
.Y(n_1343)
);

A2O1A1Ixp33_ASAP7_75t_L g1344 ( 
.A1(n_1057),
.A2(n_1060),
.B(n_910),
.C(n_1058),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1058),
.B(n_903),
.Y(n_1345)
);

OAI22x1_ASAP7_75t_L g1346 ( 
.A1(n_1058),
.A2(n_1131),
.B1(n_910),
.B2(n_1180),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_1314),
.Y(n_1347)
);

NAND3xp33_ASAP7_75t_L g1348 ( 
.A(n_1323),
.B(n_1301),
.C(n_1303),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1324),
.A2(n_1338),
.B1(n_1346),
.B2(n_1298),
.Y(n_1349)
);

A2O1A1Ixp33_ASAP7_75t_L g1350 ( 
.A1(n_1344),
.A2(n_1237),
.B(n_1298),
.C(n_1211),
.Y(n_1350)
);

AO21x2_ASAP7_75t_L g1351 ( 
.A1(n_1246),
.A2(n_1242),
.B(n_1255),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_1315),
.Y(n_1352)
);

BUFx8_ASAP7_75t_L g1353 ( 
.A(n_1226),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1334),
.B(n_1342),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1299),
.A2(n_1308),
.B1(n_1313),
.B2(n_1339),
.Y(n_1355)
);

AO31x2_ASAP7_75t_L g1356 ( 
.A1(n_1253),
.A2(n_1250),
.A3(n_1317),
.B(n_1322),
.Y(n_1356)
);

INVx3_ASAP7_75t_L g1357 ( 
.A(n_1254),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1305),
.A2(n_1312),
.B1(n_1340),
.B2(n_1345),
.Y(n_1358)
);

INVx6_ASAP7_75t_L g1359 ( 
.A(n_1217),
.Y(n_1359)
);

INVx3_ASAP7_75t_L g1360 ( 
.A(n_1254),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1320),
.A2(n_1240),
.B1(n_1205),
.B2(n_1209),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1232),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1236),
.Y(n_1363)
);

NOR4xp25_ASAP7_75t_L g1364 ( 
.A(n_1320),
.B(n_1271),
.C(n_1287),
.D(n_1209),
.Y(n_1364)
);

AOI222xp33_ASAP7_75t_L g1365 ( 
.A1(n_1258),
.A2(n_1287),
.B1(n_1271),
.B2(n_1277),
.C1(n_1290),
.C2(n_1329),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1309),
.Y(n_1366)
);

OAI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1240),
.A2(n_1278),
.B1(n_1261),
.B2(n_1211),
.Y(n_1367)
);

BUFx3_ASAP7_75t_L g1368 ( 
.A(n_1217),
.Y(n_1368)
);

OA21x2_ASAP7_75t_L g1369 ( 
.A1(n_1318),
.A2(n_1319),
.B(n_1326),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1261),
.A2(n_1276),
.B1(n_1279),
.B2(n_1334),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1218),
.A2(n_1230),
.B(n_1225),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1248),
.A2(n_1311),
.B(n_1202),
.Y(n_1372)
);

BUFx2_ASAP7_75t_L g1373 ( 
.A(n_1219),
.Y(n_1373)
);

NAND2x1p5_ASAP7_75t_L g1374 ( 
.A(n_1337),
.B(n_1266),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1342),
.B(n_1269),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1262),
.B(n_1269),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1222),
.A2(n_1220),
.B(n_1200),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1311),
.A2(n_1286),
.B1(n_1206),
.B2(n_1288),
.Y(n_1378)
);

INVx4_ASAP7_75t_SL g1379 ( 
.A(n_1342),
.Y(n_1379)
);

O2A1O1Ixp33_ASAP7_75t_SL g1380 ( 
.A1(n_1237),
.A2(n_1229),
.B(n_1289),
.C(n_1206),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1201),
.B(n_1208),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1247),
.A2(n_1272),
.B(n_1224),
.Y(n_1382)
);

INVx6_ASAP7_75t_L g1383 ( 
.A(n_1331),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1256),
.A2(n_1207),
.B(n_1260),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1280),
.A2(n_1210),
.B(n_1221),
.Y(n_1385)
);

CKINVDCx20_ASAP7_75t_R g1386 ( 
.A(n_1259),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1265),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1268),
.A2(n_1239),
.B(n_1234),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1203),
.A2(n_1228),
.B(n_1243),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1286),
.A2(n_1288),
.B1(n_1282),
.B2(n_1278),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1239),
.A2(n_1234),
.B(n_1204),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_1331),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1204),
.A2(n_1291),
.B(n_1310),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1325),
.A2(n_1332),
.B1(n_1274),
.B2(n_1321),
.Y(n_1394)
);

BUFx3_ASAP7_75t_L g1395 ( 
.A(n_1231),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1325),
.B(n_1332),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1296),
.A2(n_1304),
.B1(n_1223),
.B2(n_1336),
.Y(n_1397)
);

AO21x2_ASAP7_75t_L g1398 ( 
.A1(n_1333),
.A2(n_1241),
.B(n_1215),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1212),
.A2(n_1284),
.B1(n_1294),
.B2(n_1290),
.Y(n_1399)
);

AO31x2_ASAP7_75t_L g1400 ( 
.A1(n_1214),
.A2(n_1216),
.A3(n_1245),
.B(n_1244),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1330),
.B(n_1285),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1267),
.A2(n_1293),
.B(n_1302),
.Y(n_1402)
);

AOI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1235),
.A2(n_1306),
.B1(n_1213),
.B2(n_1283),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1275),
.B(n_1249),
.Y(n_1404)
);

BUFx3_ASAP7_75t_L g1405 ( 
.A(n_1314),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1267),
.A2(n_1245),
.B(n_1249),
.Y(n_1406)
);

INVx3_ASAP7_75t_L g1407 ( 
.A(n_1337),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1263),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1233),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1212),
.A2(n_1307),
.B1(n_1295),
.B2(n_1252),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1252),
.B(n_1251),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1233),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1327),
.A2(n_1281),
.B(n_1335),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1343),
.A2(n_1292),
.B1(n_1314),
.B2(n_1238),
.Y(n_1414)
);

A2O1A1Ixp33_ASAP7_75t_L g1415 ( 
.A1(n_1327),
.A2(n_1227),
.B(n_1341),
.C(n_1292),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_SL g1416 ( 
.A(n_1341),
.B(n_1257),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1327),
.A2(n_1341),
.B(n_1264),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1264),
.A2(n_1273),
.B(n_1328),
.Y(n_1418)
);

OAI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1301),
.A2(n_1240),
.B1(n_1058),
.B2(n_1339),
.Y(n_1419)
);

OR2x6_ASAP7_75t_L g1420 ( 
.A(n_1310),
.B(n_1215),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1324),
.A2(n_1058),
.B1(n_1346),
.B2(n_1338),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1299),
.B(n_1058),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1324),
.A2(n_1058),
.B1(n_1346),
.B2(n_1338),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1323),
.B(n_1058),
.Y(n_1424)
);

CKINVDCx8_ASAP7_75t_R g1425 ( 
.A(n_1343),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1262),
.B(n_1334),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_SL g1427 ( 
.A1(n_1258),
.A2(n_1000),
.B1(n_1160),
.B2(n_1058),
.Y(n_1427)
);

AO21x1_ASAP7_75t_L g1428 ( 
.A1(n_1323),
.A2(n_1298),
.B(n_1320),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1265),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1299),
.B(n_1058),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1270),
.B(n_1325),
.Y(n_1431)
);

INVx3_ASAP7_75t_L g1432 ( 
.A(n_1254),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1297),
.A2(n_1316),
.B(n_1300),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1297),
.A2(n_1316),
.B(n_1300),
.Y(n_1434)
);

BUFx3_ASAP7_75t_L g1435 ( 
.A(n_1309),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1297),
.A2(n_1316),
.B(n_1300),
.Y(n_1436)
);

AO31x2_ASAP7_75t_L g1437 ( 
.A1(n_1253),
.A2(n_1246),
.A3(n_1250),
.B(n_1255),
.Y(n_1437)
);

AOI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1324),
.A2(n_1011),
.B1(n_910),
.B2(n_1058),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1254),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1291),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1323),
.A2(n_1011),
.B(n_1303),
.Y(n_1441)
);

INVx3_ASAP7_75t_L g1442 ( 
.A(n_1254),
.Y(n_1442)
);

O2A1O1Ixp33_ASAP7_75t_L g1443 ( 
.A1(n_1323),
.A2(n_1344),
.B(n_1303),
.C(n_1011),
.Y(n_1443)
);

CKINVDCx16_ASAP7_75t_R g1444 ( 
.A(n_1257),
.Y(n_1444)
);

OAI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1323),
.A2(n_1011),
.B(n_1303),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1324),
.A2(n_1058),
.B1(n_1346),
.B2(n_1338),
.Y(n_1446)
);

OAI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1323),
.A2(n_1011),
.B(n_1303),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1265),
.Y(n_1448)
);

NOR2xp67_ASAP7_75t_L g1449 ( 
.A(n_1296),
.B(n_716),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1317),
.A2(n_1319),
.B(n_1318),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1317),
.A2(n_1319),
.B(n_1318),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_1217),
.Y(n_1452)
);

NOR2xp67_ASAP7_75t_SL g1453 ( 
.A(n_1343),
.B(n_634),
.Y(n_1453)
);

OR2x6_ASAP7_75t_L g1454 ( 
.A(n_1310),
.B(n_1215),
.Y(n_1454)
);

BUFx2_ASAP7_75t_L g1455 ( 
.A(n_1315),
.Y(n_1455)
);

INVxp67_ASAP7_75t_SL g1456 ( 
.A(n_1237),
.Y(n_1456)
);

AO21x2_ASAP7_75t_L g1457 ( 
.A1(n_1246),
.A2(n_1242),
.B(n_1255),
.Y(n_1457)
);

NAND3xp33_ASAP7_75t_L g1458 ( 
.A(n_1323),
.B(n_1011),
.C(n_784),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1323),
.A2(n_1011),
.B(n_1303),
.Y(n_1459)
);

A2O1A1Ixp33_ASAP7_75t_L g1460 ( 
.A1(n_1323),
.A2(n_1058),
.B(n_1057),
.C(n_1303),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1265),
.Y(n_1461)
);

A2O1A1Ixp33_ASAP7_75t_L g1462 ( 
.A1(n_1323),
.A2(n_1058),
.B(n_1057),
.C(n_1303),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1232),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1262),
.B(n_1334),
.Y(n_1464)
);

AOI211xp5_ASAP7_75t_L g1465 ( 
.A1(n_1427),
.A2(n_1367),
.B(n_1458),
.C(n_1447),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1376),
.B(n_1426),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_SL g1467 ( 
.A1(n_1443),
.A2(n_1445),
.B(n_1441),
.Y(n_1467)
);

A2O1A1Ixp33_ASAP7_75t_L g1468 ( 
.A1(n_1459),
.A2(n_1438),
.B(n_1424),
.C(n_1348),
.Y(n_1468)
);

O2A1O1Ixp5_ASAP7_75t_L g1469 ( 
.A1(n_1428),
.A2(n_1382),
.B(n_1460),
.C(n_1462),
.Y(n_1469)
);

O2A1O1Ixp33_ASAP7_75t_L g1470 ( 
.A1(n_1460),
.A2(n_1462),
.B(n_1424),
.C(n_1419),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1355),
.B(n_1358),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1422),
.B(n_1430),
.Y(n_1472)
);

NOR2xp67_ASAP7_75t_L g1473 ( 
.A(n_1452),
.B(n_1397),
.Y(n_1473)
);

AOI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1450),
.A2(n_1451),
.B(n_1372),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1381),
.B(n_1408),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1379),
.B(n_1354),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1379),
.B(n_1354),
.Y(n_1477)
);

A2O1A1Ixp33_ASAP7_75t_SL g1478 ( 
.A1(n_1421),
.A2(n_1446),
.B(n_1423),
.C(n_1389),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1464),
.B(n_1421),
.Y(n_1479)
);

OAI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1361),
.A2(n_1446),
.B1(n_1423),
.B2(n_1399),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1396),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1362),
.B(n_1363),
.Y(n_1482)
);

NOR2xp67_ASAP7_75t_L g1483 ( 
.A(n_1403),
.B(n_1411),
.Y(n_1483)
);

OA21x2_ASAP7_75t_L g1484 ( 
.A1(n_1388),
.A2(n_1391),
.B(n_1433),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1404),
.B(n_1349),
.Y(n_1485)
);

AOI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1369),
.A2(n_1456),
.B(n_1420),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1366),
.Y(n_1487)
);

OA21x2_ASAP7_75t_L g1488 ( 
.A1(n_1388),
.A2(n_1391),
.B(n_1434),
.Y(n_1488)
);

OR2x6_ASAP7_75t_L g1489 ( 
.A(n_1420),
.B(n_1454),
.Y(n_1489)
);

NOR2xp67_ASAP7_75t_L g1490 ( 
.A(n_1411),
.B(n_1449),
.Y(n_1490)
);

O2A1O1Ixp33_ASAP7_75t_L g1491 ( 
.A1(n_1419),
.A2(n_1367),
.B(n_1350),
.C(n_1364),
.Y(n_1491)
);

AOI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1456),
.A2(n_1454),
.B(n_1420),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1349),
.B(n_1431),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1361),
.A2(n_1399),
.B1(n_1350),
.B2(n_1390),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1463),
.B(n_1373),
.Y(n_1495)
);

INVx2_ASAP7_75t_SL g1496 ( 
.A(n_1359),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1365),
.B(n_1370),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1352),
.B(n_1455),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1375),
.B(n_1394),
.Y(n_1499)
);

O2A1O1Ixp5_ASAP7_75t_L g1500 ( 
.A1(n_1409),
.A2(n_1412),
.B(n_1415),
.C(n_1429),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1390),
.A2(n_1378),
.B1(n_1425),
.B2(n_1410),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1401),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1378),
.A2(n_1410),
.B1(n_1414),
.B2(n_1416),
.Y(n_1503)
);

AOI211xp5_ASAP7_75t_L g1504 ( 
.A1(n_1380),
.A2(n_1453),
.B(n_1416),
.C(n_1418),
.Y(n_1504)
);

BUFx6f_ASAP7_75t_L g1505 ( 
.A(n_1366),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1406),
.Y(n_1506)
);

CKINVDCx20_ASAP7_75t_R g1507 ( 
.A(n_1386),
.Y(n_1507)
);

A2O1A1Ixp33_ASAP7_75t_L g1508 ( 
.A1(n_1393),
.A2(n_1417),
.B(n_1413),
.C(n_1440),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1374),
.B(n_1444),
.Y(n_1509)
);

AOI21xp5_ASAP7_75t_SL g1510 ( 
.A1(n_1347),
.A2(n_1405),
.B(n_1374),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1400),
.B(n_1457),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1437),
.Y(n_1512)
);

AOI21xp5_ASAP7_75t_SL g1513 ( 
.A1(n_1347),
.A2(n_1405),
.B(n_1392),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1437),
.B(n_1351),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_R g1515 ( 
.A(n_1386),
.B(n_1383),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1437),
.B(n_1351),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1353),
.B(n_1395),
.Y(n_1517)
);

O2A1O1Ixp33_ASAP7_75t_L g1518 ( 
.A1(n_1398),
.A2(n_1395),
.B(n_1461),
.C(n_1387),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1402),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1353),
.B(n_1398),
.Y(n_1520)
);

AOI221xp5_ASAP7_75t_L g1521 ( 
.A1(n_1435),
.A2(n_1392),
.B1(n_1368),
.B2(n_1448),
.C(n_1360),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1353),
.B(n_1356),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1357),
.B(n_1360),
.Y(n_1523)
);

O2A1O1Ixp5_ASAP7_75t_L g1524 ( 
.A1(n_1357),
.A2(n_1442),
.B(n_1439),
.C(n_1432),
.Y(n_1524)
);

O2A1O1Ixp5_ASAP7_75t_L g1525 ( 
.A1(n_1407),
.A2(n_1442),
.B(n_1432),
.C(n_1356),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1356),
.B(n_1435),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1359),
.B(n_1383),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1359),
.B(n_1383),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1385),
.B(n_1384),
.Y(n_1529)
);

NOR2xp67_ASAP7_75t_L g1530 ( 
.A(n_1377),
.B(n_1371),
.Y(n_1530)
);

BUFx2_ASAP7_75t_L g1531 ( 
.A(n_1377),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1436),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1396),
.Y(n_1533)
);

NOR2x1_ASAP7_75t_SL g1534 ( 
.A(n_1420),
.B(n_1454),
.Y(n_1534)
);

AOI21xp5_ASAP7_75t_SL g1535 ( 
.A1(n_1443),
.A2(n_813),
.B(n_1323),
.Y(n_1535)
);

O2A1O1Ixp5_ASAP7_75t_L g1536 ( 
.A1(n_1441),
.A2(n_1445),
.B(n_1459),
.C(n_1447),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1431),
.B(n_1396),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1355),
.B(n_1358),
.Y(n_1538)
);

AOI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1450),
.A2(n_1451),
.B(n_1372),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1355),
.B(n_1358),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1427),
.A2(n_1438),
.B1(n_1058),
.B2(n_1240),
.Y(n_1541)
);

O2A1O1Ixp33_ASAP7_75t_L g1542 ( 
.A1(n_1441),
.A2(n_1323),
.B(n_1447),
.C(n_1445),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1427),
.A2(n_1438),
.B1(n_1058),
.B2(n_1240),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1422),
.B(n_794),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1379),
.B(n_1354),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1427),
.A2(n_1438),
.B1(n_1058),
.B2(n_1240),
.Y(n_1546)
);

A2O1A1Ixp33_ASAP7_75t_L g1547 ( 
.A1(n_1443),
.A2(n_1323),
.B(n_910),
.C(n_1458),
.Y(n_1547)
);

BUFx3_ASAP7_75t_L g1548 ( 
.A(n_1366),
.Y(n_1548)
);

AOI221x1_ASAP7_75t_SL g1549 ( 
.A1(n_1367),
.A2(n_814),
.B1(n_797),
.B2(n_1101),
.C(n_1419),
.Y(n_1549)
);

AOI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1450),
.A2(n_1451),
.B(n_1372),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1355),
.B(n_1358),
.Y(n_1551)
);

OA21x2_ASAP7_75t_L g1552 ( 
.A1(n_1382),
.A2(n_1246),
.B(n_1388),
.Y(n_1552)
);

O2A1O1Ixp33_ASAP7_75t_L g1553 ( 
.A1(n_1441),
.A2(n_1323),
.B(n_1447),
.C(n_1445),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1355),
.B(n_1358),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1376),
.B(n_1426),
.Y(n_1555)
);

INVx3_ASAP7_75t_L g1556 ( 
.A(n_1375),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1355),
.B(n_1358),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1376),
.B(n_1426),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1514),
.B(n_1516),
.Y(n_1559)
);

INVx3_ASAP7_75t_L g1560 ( 
.A(n_1484),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1506),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1471),
.B(n_1538),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1512),
.B(n_1552),
.Y(n_1563)
);

INVxp67_ASAP7_75t_L g1564 ( 
.A(n_1526),
.Y(n_1564)
);

AO21x2_ASAP7_75t_L g1565 ( 
.A1(n_1474),
.A2(n_1550),
.B(n_1539),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1552),
.B(n_1511),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1540),
.B(n_1551),
.Y(n_1567)
);

AO21x2_ASAP7_75t_L g1568 ( 
.A1(n_1486),
.A2(n_1518),
.B(n_1467),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1500),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1519),
.B(n_1529),
.Y(n_1570)
);

INVx4_ASAP7_75t_L g1571 ( 
.A(n_1489),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1554),
.B(n_1557),
.Y(n_1572)
);

BUFx6f_ASAP7_75t_L g1573 ( 
.A(n_1488),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1500),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1531),
.B(n_1508),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1532),
.B(n_1493),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1485),
.B(n_1522),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1536),
.B(n_1469),
.Y(n_1578)
);

AO21x2_ASAP7_75t_L g1579 ( 
.A1(n_1518),
.A2(n_1542),
.B(n_1553),
.Y(n_1579)
);

INVxp67_ASAP7_75t_SL g1580 ( 
.A(n_1542),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1520),
.Y(n_1581)
);

AO21x2_ASAP7_75t_L g1582 ( 
.A1(n_1553),
.A2(n_1468),
.B(n_1530),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1541),
.A2(n_1546),
.B1(n_1543),
.B2(n_1480),
.Y(n_1583)
);

BUFx2_ASAP7_75t_SL g1584 ( 
.A(n_1473),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1525),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1525),
.Y(n_1586)
);

AOI21xp5_ASAP7_75t_L g1587 ( 
.A1(n_1469),
.A2(n_1547),
.B(n_1492),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_SL g1588 ( 
.A(n_1491),
.B(n_1470),
.Y(n_1588)
);

OR2x6_ASAP7_75t_L g1589 ( 
.A(n_1489),
.B(n_1492),
.Y(n_1589)
);

INVx3_ASAP7_75t_L g1590 ( 
.A(n_1489),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1482),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1524),
.Y(n_1592)
);

INVx5_ASAP7_75t_L g1593 ( 
.A(n_1476),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1470),
.B(n_1475),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1491),
.B(n_1481),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1534),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_1507),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1533),
.B(n_1537),
.Y(n_1598)
);

AO21x1_ASAP7_75t_L g1599 ( 
.A1(n_1465),
.A2(n_1494),
.B(n_1497),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1472),
.B(n_1502),
.Y(n_1600)
);

AO21x2_ASAP7_75t_L g1601 ( 
.A1(n_1478),
.A2(n_1535),
.B(n_1501),
.Y(n_1601)
);

NOR3xp33_ASAP7_75t_L g1602 ( 
.A(n_1504),
.B(n_1503),
.C(n_1544),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_SL g1603 ( 
.A1(n_1527),
.A2(n_1528),
.B(n_1521),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1566),
.B(n_1479),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1599),
.A2(n_1583),
.B1(n_1588),
.B2(n_1602),
.Y(n_1605)
);

NOR2x1_ASAP7_75t_L g1606 ( 
.A(n_1584),
.B(n_1582),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1592),
.Y(n_1607)
);

NOR2x1p5_ASAP7_75t_L g1608 ( 
.A(n_1580),
.B(n_1556),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1566),
.B(n_1499),
.Y(n_1609)
);

INVxp67_ASAP7_75t_SL g1610 ( 
.A(n_1592),
.Y(n_1610)
);

NAND3xp33_ASAP7_75t_L g1611 ( 
.A(n_1588),
.B(n_1483),
.C(n_1495),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1564),
.B(n_1498),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1561),
.Y(n_1613)
);

INVx3_ASAP7_75t_L g1614 ( 
.A(n_1573),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1560),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1570),
.B(n_1477),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1559),
.B(n_1466),
.Y(n_1617)
);

AND2x2_ASAP7_75t_SL g1618 ( 
.A(n_1571),
.B(n_1545),
.Y(n_1618)
);

INVx3_ASAP7_75t_L g1619 ( 
.A(n_1573),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1559),
.B(n_1558),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1563),
.B(n_1555),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1592),
.Y(n_1622)
);

NAND2x1_ASAP7_75t_L g1623 ( 
.A(n_1589),
.B(n_1510),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1580),
.B(n_1549),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1564),
.B(n_1523),
.Y(n_1625)
);

AOI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1605),
.A2(n_1599),
.B1(n_1583),
.B2(n_1602),
.Y(n_1626)
);

NAND3xp33_ASAP7_75t_SL g1627 ( 
.A(n_1605),
.B(n_1599),
.C(n_1587),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_SL g1628 ( 
.A1(n_1611),
.A2(n_1601),
.B1(n_1578),
.B2(n_1587),
.Y(n_1628)
);

AOI33xp33_ASAP7_75t_L g1629 ( 
.A1(n_1604),
.A2(n_1578),
.A3(n_1577),
.B1(n_1574),
.B2(n_1569),
.B3(n_1591),
.Y(n_1629)
);

BUFx3_ASAP7_75t_L g1630 ( 
.A(n_1612),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_1612),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1611),
.A2(n_1601),
.B1(n_1578),
.B2(n_1567),
.Y(n_1632)
);

AOI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1624),
.A2(n_1601),
.B1(n_1567),
.B2(n_1594),
.Y(n_1633)
);

INVx4_ASAP7_75t_SL g1634 ( 
.A(n_1616),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1606),
.B(n_1589),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1624),
.A2(n_1601),
.B1(n_1582),
.B2(n_1571),
.Y(n_1636)
);

INVxp67_ASAP7_75t_SL g1637 ( 
.A(n_1607),
.Y(n_1637)
);

NAND4xp25_ASAP7_75t_L g1638 ( 
.A(n_1612),
.B(n_1562),
.C(n_1572),
.D(n_1595),
.Y(n_1638)
);

INVx5_ASAP7_75t_SL g1639 ( 
.A(n_1618),
.Y(n_1639)
);

NOR3xp33_ASAP7_75t_SL g1640 ( 
.A(n_1625),
.B(n_1595),
.C(n_1597),
.Y(n_1640)
);

NAND3xp33_ASAP7_75t_L g1641 ( 
.A(n_1607),
.B(n_1594),
.C(n_1572),
.Y(n_1641)
);

AOI31xp33_ASAP7_75t_L g1642 ( 
.A1(n_1610),
.A2(n_1562),
.A3(n_1596),
.B(n_1509),
.Y(n_1642)
);

OA21x2_ASAP7_75t_L g1643 ( 
.A1(n_1615),
.A2(n_1586),
.B(n_1585),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1618),
.A2(n_1601),
.B1(n_1582),
.B2(n_1571),
.Y(n_1644)
);

OAI222xp33_ASAP7_75t_L g1645 ( 
.A1(n_1604),
.A2(n_1576),
.B1(n_1589),
.B2(n_1577),
.C1(n_1581),
.C2(n_1571),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1618),
.B(n_1515),
.Y(n_1646)
);

OAI31xp33_ASAP7_75t_L g1647 ( 
.A1(n_1608),
.A2(n_1581),
.A3(n_1576),
.B(n_1600),
.Y(n_1647)
);

BUFx3_ASAP7_75t_L g1648 ( 
.A(n_1623),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1604),
.B(n_1581),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1618),
.A2(n_1582),
.B1(n_1579),
.B2(n_1577),
.Y(n_1650)
);

INVxp67_ASAP7_75t_L g1651 ( 
.A(n_1625),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1614),
.B(n_1619),
.Y(n_1652)
);

OAI211xp5_ASAP7_75t_L g1653 ( 
.A1(n_1623),
.A2(n_1603),
.B(n_1600),
.C(n_1574),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1613),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1608),
.A2(n_1584),
.B1(n_1589),
.B2(n_1593),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1616),
.A2(n_1582),
.B1(n_1579),
.B2(n_1590),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1609),
.B(n_1575),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1617),
.B(n_1598),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_1617),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_SL g1660 ( 
.A(n_1616),
.B(n_1593),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1613),
.Y(n_1661)
);

AOI31xp33_ASAP7_75t_L g1662 ( 
.A1(n_1622),
.A2(n_1596),
.A3(n_1576),
.B(n_1598),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1643),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1654),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1633),
.B(n_1621),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1654),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1634),
.B(n_1614),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1657),
.B(n_1617),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1630),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_SL g1670 ( 
.A(n_1633),
.B(n_1593),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1661),
.Y(n_1671)
);

AND2x6_ASAP7_75t_SL g1672 ( 
.A(n_1658),
.B(n_1517),
.Y(n_1672)
);

INVx4_ASAP7_75t_SL g1673 ( 
.A(n_1648),
.Y(n_1673)
);

CKINVDCx14_ASAP7_75t_R g1674 ( 
.A(n_1659),
.Y(n_1674)
);

BUFx2_ASAP7_75t_L g1675 ( 
.A(n_1634),
.Y(n_1675)
);

INVx3_ASAP7_75t_L g1676 ( 
.A(n_1643),
.Y(n_1676)
);

INVxp67_ASAP7_75t_SL g1677 ( 
.A(n_1641),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1630),
.Y(n_1678)
);

AOI21xp5_ASAP7_75t_SL g1679 ( 
.A1(n_1627),
.A2(n_1568),
.B(n_1565),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1634),
.B(n_1620),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1629),
.B(n_1621),
.Y(n_1681)
);

INVx4_ASAP7_75t_SL g1682 ( 
.A(n_1648),
.Y(n_1682)
);

BUFx3_ASAP7_75t_L g1683 ( 
.A(n_1631),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1637),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1631),
.Y(n_1685)
);

INVx4_ASAP7_75t_SL g1686 ( 
.A(n_1635),
.Y(n_1686)
);

HB1xp67_ASAP7_75t_L g1687 ( 
.A(n_1649),
.Y(n_1687)
);

INVx4_ASAP7_75t_SL g1688 ( 
.A(n_1635),
.Y(n_1688)
);

BUFx2_ASAP7_75t_L g1689 ( 
.A(n_1635),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1651),
.B(n_1621),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1638),
.B(n_1598),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1664),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1664),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1666),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1677),
.B(n_1638),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1663),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1675),
.B(n_1639),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1663),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1673),
.B(n_1660),
.Y(n_1699)
);

NOR2x1_ASAP7_75t_L g1700 ( 
.A(n_1683),
.B(n_1641),
.Y(n_1700)
);

NOR2x1_ASAP7_75t_L g1701 ( 
.A(n_1683),
.B(n_1653),
.Y(n_1701)
);

OAI222xp33_ASAP7_75t_L g1702 ( 
.A1(n_1670),
.A2(n_1626),
.B1(n_1628),
.B2(n_1632),
.C1(n_1665),
.C2(n_1681),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_SL g1703 ( 
.A(n_1691),
.B(n_1647),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1666),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1675),
.B(n_1639),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1686),
.B(n_1639),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1673),
.B(n_1652),
.Y(n_1707)
);

OAI221xp5_ASAP7_75t_L g1708 ( 
.A1(n_1679),
.A2(n_1626),
.B1(n_1636),
.B2(n_1640),
.C(n_1644),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1681),
.B(n_1620),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1686),
.B(n_1639),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1665),
.B(n_1662),
.Y(n_1711)
);

INVx1_ASAP7_75t_SL g1712 ( 
.A(n_1683),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1671),
.Y(n_1713)
);

AOI211x1_ASAP7_75t_L g1714 ( 
.A1(n_1685),
.A2(n_1662),
.B(n_1642),
.C(n_1645),
.Y(n_1714)
);

INVxp67_ASAP7_75t_L g1715 ( 
.A(n_1669),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1684),
.B(n_1642),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1676),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1688),
.B(n_1647),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1688),
.B(n_1659),
.Y(n_1719)
);

INVx2_ASAP7_75t_SL g1720 ( 
.A(n_1667),
.Y(n_1720)
);

INVx3_ASAP7_75t_L g1721 ( 
.A(n_1667),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_SL g1722 ( 
.A(n_1680),
.B(n_1646),
.Y(n_1722)
);

INVx3_ASAP7_75t_L g1723 ( 
.A(n_1699),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1717),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1692),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1717),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1706),
.B(n_1688),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1692),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1720),
.B(n_1706),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1715),
.B(n_1695),
.Y(n_1730)
);

INVxp67_ASAP7_75t_L g1731 ( 
.A(n_1701),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1715),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1712),
.B(n_1672),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1717),
.Y(n_1734)
);

AOI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1708),
.A2(n_1650),
.B1(n_1656),
.B2(n_1655),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1710),
.B(n_1688),
.Y(n_1736)
);

INVx3_ASAP7_75t_L g1737 ( 
.A(n_1699),
.Y(n_1737)
);

CKINVDCx16_ASAP7_75t_R g1738 ( 
.A(n_1701),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1693),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1693),
.Y(n_1740)
);

INVxp67_ASAP7_75t_L g1741 ( 
.A(n_1712),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1694),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1694),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1695),
.B(n_1672),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1704),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1709),
.B(n_1678),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1696),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1709),
.B(n_1668),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1710),
.B(n_1688),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1704),
.Y(n_1750)
);

AOI22xp33_ASAP7_75t_SL g1751 ( 
.A1(n_1708),
.A2(n_1674),
.B1(n_1565),
.B2(n_1689),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_SL g1752 ( 
.A(n_1700),
.B(n_1680),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1720),
.B(n_1673),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1720),
.B(n_1673),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1719),
.B(n_1673),
.Y(n_1755)
);

OAI22xp33_ASAP7_75t_L g1756 ( 
.A1(n_1711),
.A2(n_1689),
.B1(n_1690),
.B2(n_1687),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1699),
.B(n_1682),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1713),
.Y(n_1758)
);

INVxp67_ASAP7_75t_L g1759 ( 
.A(n_1732),
.Y(n_1759)
);

INVx2_ASAP7_75t_SL g1760 ( 
.A(n_1753),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1730),
.B(n_1711),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1755),
.B(n_1697),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1751),
.A2(n_1703),
.B1(n_1700),
.B2(n_1718),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1755),
.B(n_1697),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1738),
.B(n_1714),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1758),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1758),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1725),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1725),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1731),
.B(n_1714),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1723),
.Y(n_1771)
);

AND2x2_ASAP7_75t_SL g1772 ( 
.A(n_1752),
.B(n_1718),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1728),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1728),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1742),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1742),
.Y(n_1776)
);

INVx1_ASAP7_75t_SL g1777 ( 
.A(n_1727),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1727),
.B(n_1705),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1723),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1743),
.Y(n_1780)
);

CKINVDCx16_ASAP7_75t_R g1781 ( 
.A(n_1730),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1723),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1741),
.B(n_1744),
.Y(n_1783)
);

HB1xp67_ASAP7_75t_L g1784 ( 
.A(n_1737),
.Y(n_1784)
);

INVxp67_ASAP7_75t_L g1785 ( 
.A(n_1733),
.Y(n_1785)
);

OAI21xp33_ASAP7_75t_SL g1786 ( 
.A1(n_1772),
.A2(n_1749),
.B(n_1736),
.Y(n_1786)
);

INVx1_ASAP7_75t_SL g1787 ( 
.A(n_1772),
.Y(n_1787)
);

NAND2xp33_ASAP7_75t_L g1788 ( 
.A(n_1763),
.B(n_1736),
.Y(n_1788)
);

INVxp67_ASAP7_75t_SL g1789 ( 
.A(n_1784),
.Y(n_1789)
);

A2O1A1Ixp33_ASAP7_75t_L g1790 ( 
.A1(n_1765),
.A2(n_1735),
.B(n_1716),
.C(n_1757),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1766),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_L g1792 ( 
.A(n_1781),
.B(n_1702),
.Y(n_1792)
);

NAND2x1p5_ASAP7_75t_L g1793 ( 
.A(n_1772),
.B(n_1757),
.Y(n_1793)
);

AOI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1770),
.A2(n_1757),
.B1(n_1749),
.B2(n_1756),
.Y(n_1794)
);

OAI21xp33_ASAP7_75t_L g1795 ( 
.A1(n_1777),
.A2(n_1746),
.B(n_1679),
.Y(n_1795)
);

NAND2xp33_ASAP7_75t_SL g1796 ( 
.A(n_1762),
.B(n_1719),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1781),
.B(n_1729),
.Y(n_1797)
);

NAND2xp33_ASAP7_75t_L g1798 ( 
.A(n_1762),
.B(n_1705),
.Y(n_1798)
);

OAI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1785),
.A2(n_1737),
.B1(n_1722),
.B2(n_1716),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1766),
.Y(n_1800)
);

AOI21xp33_ASAP7_75t_SL g1801 ( 
.A1(n_1761),
.A2(n_1759),
.B(n_1783),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1764),
.B(n_1729),
.Y(n_1802)
);

AOI21xp5_ASAP7_75t_L g1803 ( 
.A1(n_1761),
.A2(n_1702),
.B(n_1729),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1764),
.B(n_1778),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1760),
.B(n_1737),
.Y(n_1805)
);

INVxp67_ASAP7_75t_L g1806 ( 
.A(n_1778),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1789),
.B(n_1806),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1791),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1787),
.B(n_1760),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1800),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1792),
.A2(n_1788),
.B1(n_1804),
.B2(n_1796),
.Y(n_1811)
);

BUFx6f_ASAP7_75t_L g1812 ( 
.A(n_1793),
.Y(n_1812)
);

INVxp33_ASAP7_75t_L g1813 ( 
.A(n_1793),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1805),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1797),
.B(n_1771),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1802),
.B(n_1771),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1798),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1801),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1799),
.Y(n_1819)
);

NAND3xp33_ASAP7_75t_L g1820 ( 
.A(n_1818),
.B(n_1790),
.C(n_1803),
.Y(n_1820)
);

AOI221xp5_ASAP7_75t_L g1821 ( 
.A1(n_1811),
.A2(n_1794),
.B1(n_1795),
.B2(n_1786),
.C(n_1769),
.Y(n_1821)
);

NOR2x1_ASAP7_75t_L g1822 ( 
.A(n_1807),
.B(n_1779),
.Y(n_1822)
);

AOI211xp5_ASAP7_75t_L g1823 ( 
.A1(n_1813),
.A2(n_1819),
.B(n_1817),
.C(n_1809),
.Y(n_1823)
);

OAI211xp5_ASAP7_75t_L g1824 ( 
.A1(n_1819),
.A2(n_1782),
.B(n_1779),
.C(n_1780),
.Y(n_1824)
);

AOI211xp5_ASAP7_75t_L g1825 ( 
.A1(n_1813),
.A2(n_1782),
.B(n_1754),
.C(n_1753),
.Y(n_1825)
);

NAND4xp25_ASAP7_75t_L g1826 ( 
.A(n_1815),
.B(n_1780),
.C(n_1776),
.D(n_1775),
.Y(n_1826)
);

NOR3xp33_ASAP7_75t_SL g1827 ( 
.A(n_1814),
.B(n_1768),
.C(n_1767),
.Y(n_1827)
);

AOI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1815),
.A2(n_1754),
.B1(n_1753),
.B2(n_1699),
.Y(n_1828)
);

AOI21xp5_ASAP7_75t_L g1829 ( 
.A1(n_1807),
.A2(n_1768),
.B(n_1767),
.Y(n_1829)
);

OAI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1820),
.A2(n_1816),
.B(n_1810),
.Y(n_1830)
);

OAI22xp5_ASAP7_75t_SL g1831 ( 
.A1(n_1823),
.A2(n_1812),
.B1(n_1808),
.B2(n_1754),
.Y(n_1831)
);

NAND3xp33_ASAP7_75t_L g1832 ( 
.A(n_1827),
.B(n_1812),
.C(n_1816),
.Y(n_1832)
);

INVx1_ASAP7_75t_SL g1833 ( 
.A(n_1822),
.Y(n_1833)
);

INVx1_ASAP7_75t_SL g1834 ( 
.A(n_1828),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1821),
.B(n_1812),
.Y(n_1835)
);

NOR3xp33_ASAP7_75t_L g1836 ( 
.A(n_1835),
.B(n_1824),
.C(n_1825),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1833),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1832),
.Y(n_1838)
);

AOI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1830),
.A2(n_1829),
.B(n_1812),
.Y(n_1839)
);

INVx3_ASAP7_75t_L g1840 ( 
.A(n_1834),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1831),
.B(n_1826),
.Y(n_1841)
);

OAI211xp5_ASAP7_75t_L g1842 ( 
.A1(n_1839),
.A2(n_1776),
.B(n_1775),
.C(n_1774),
.Y(n_1842)
);

XNOR2xp5_ASAP7_75t_L g1843 ( 
.A(n_1840),
.B(n_1490),
.Y(n_1843)
);

NAND4xp25_ASAP7_75t_L g1844 ( 
.A(n_1836),
.B(n_1774),
.C(n_1773),
.D(n_1769),
.Y(n_1844)
);

OAI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1838),
.A2(n_1721),
.B1(n_1773),
.B2(n_1740),
.Y(n_1845)
);

AOI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1837),
.A2(n_1739),
.B1(n_1707),
.B2(n_1750),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1843),
.Y(n_1847)
);

NOR4xp75_ASAP7_75t_L g1848 ( 
.A(n_1845),
.B(n_1841),
.C(n_1721),
.D(n_1748),
.Y(n_1848)
);

NAND4xp25_ASAP7_75t_L g1849 ( 
.A(n_1846),
.B(n_1724),
.C(n_1726),
.D(n_1734),
.Y(n_1849)
);

AND3x4_ASAP7_75t_L g1850 ( 
.A(n_1848),
.B(n_1844),
.C(n_1842),
.Y(n_1850)
);

AOI322xp5_ASAP7_75t_L g1851 ( 
.A1(n_1850),
.A2(n_1847),
.A3(n_1724),
.B1(n_1726),
.B2(n_1734),
.C1(n_1750),
.C2(n_1745),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1851),
.Y(n_1852)
);

HB1xp67_ASAP7_75t_L g1853 ( 
.A(n_1851),
.Y(n_1853)
);

AOI22xp33_ASAP7_75t_L g1854 ( 
.A1(n_1852),
.A2(n_1849),
.B1(n_1747),
.B2(n_1743),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1853),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1855),
.B(n_1721),
.Y(n_1856)
);

OAI22xp5_ASAP7_75t_SL g1857 ( 
.A1(n_1854),
.A2(n_1548),
.B1(n_1745),
.B2(n_1496),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1856),
.B(n_1721),
.Y(n_1858)
);

NAND2x1_ASAP7_75t_L g1859 ( 
.A(n_1858),
.B(n_1857),
.Y(n_1859)
);

AOI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1859),
.A2(n_1747),
.B1(n_1707),
.B2(n_1696),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1860),
.Y(n_1861)
);

AOI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1861),
.A2(n_1707),
.B1(n_1698),
.B2(n_1696),
.Y(n_1862)
);

AOI211xp5_ASAP7_75t_L g1863 ( 
.A1(n_1862),
.A2(n_1487),
.B(n_1505),
.C(n_1513),
.Y(n_1863)
);


endmodule