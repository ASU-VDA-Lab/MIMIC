module fake_ariane_1141_n_775 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_136, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_775);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_775;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_424;
wire n_584;
wire n_528;
wire n_387;
wire n_406;
wire n_139;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_138;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_140;
wire n_725;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_143;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_331;
wire n_320;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_699;
wire n_727;
wire n_590;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_141;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_616;
wire n_658;
wire n_617;
wire n_705;
wire n_630;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_769;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_147;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_47),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_3),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_123),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_137),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_55),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_8),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_126),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_18),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_121),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_87),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_30),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_27),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_83),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_21),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_106),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_84),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_59),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_116),
.Y(n_162)
);

BUFx8_ASAP7_75t_SL g163 ( 
.A(n_120),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_76),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_73),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_5),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_90),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_128),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_108),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_6),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_125),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_46),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_117),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_54),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_132),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_31),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_104),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_131),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_112),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_133),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_72),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_101),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_93),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_0),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_85),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_8),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_32),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_119),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_33),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_63),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_69),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_4),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_48),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_156),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_146),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_156),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_146),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

AND2x4_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_0),
.Y(n_203)
);

OA21x2_ASAP7_75t_L g204 ( 
.A1(n_140),
.A2(n_1),
.B(n_2),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_141),
.B(n_1),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_2),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_139),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_170),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_166),
.Y(n_211)
);

OAI22x1_ASAP7_75t_SL g212 ( 
.A1(n_194),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_143),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_171),
.Y(n_214)
);

OA21x2_ASAP7_75t_L g215 ( 
.A1(n_148),
.A2(n_6),
.B(n_7),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_170),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_163),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_149),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_145),
.B(n_7),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_178),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_170),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g223 ( 
.A(n_138),
.Y(n_223)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_145),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_157),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_158),
.B(n_9),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_159),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_170),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_160),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_164),
.B(n_9),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g232 ( 
.A(n_142),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_165),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_167),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_151),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_177),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_181),
.B(n_10),
.Y(n_237)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_144),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_223),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_223),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_234),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_234),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_232),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_232),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_234),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_218),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_238),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_234),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_238),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_225),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_206),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_238),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_209),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_234),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_211),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_201),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_201),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_213),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_213),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_196),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_207),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_214),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_214),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_196),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_198),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_207),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_199),
.B(n_184),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_198),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_R g271 ( 
.A(n_206),
.B(n_161),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_197),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_199),
.B(n_147),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_236),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_202),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_236),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_197),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_202),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_208),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_225),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_225),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_206),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_200),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_217),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_200),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_230),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_220),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_264),
.Y(n_288)
);

NOR2xp67_ASAP7_75t_SL g289 ( 
.A(n_249),
.B(n_204),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_240),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_220),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_231),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_260),
.B(n_203),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_239),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_252),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_251),
.B(n_231),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_265),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_261),
.B(n_203),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_259),
.B(n_203),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_254),
.B(n_237),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_272),
.B(n_237),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_253),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_273),
.B(n_219),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_253),
.B(n_219),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_284),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_258),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_274),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_239),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_239),
.Y(n_310)
);

NAND2x1_ASAP7_75t_L g311 ( 
.A(n_275),
.B(n_230),
.Y(n_311)
);

NOR3xp33_ASAP7_75t_L g312 ( 
.A(n_269),
.B(n_235),
.C(n_227),
.Y(n_312)
);

NOR3xp33_ASAP7_75t_L g313 ( 
.A(n_269),
.B(n_205),
.C(n_230),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_277),
.B(n_226),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_283),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_262),
.B(n_226),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_239),
.Y(n_317)
);

NAND3xp33_ASAP7_75t_L g318 ( 
.A(n_255),
.B(n_233),
.C(n_228),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_275),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_276),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_266),
.B(n_228),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_278),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_267),
.B(n_233),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_270),
.B(n_217),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_278),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_279),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_279),
.B(n_243),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_244),
.B(n_224),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_287),
.B(n_221),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_247),
.B(n_250),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_256),
.Y(n_331)
);

NAND2xp33_ASAP7_75t_L g332 ( 
.A(n_248),
.B(n_150),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_281),
.Y(n_333)
);

NAND2xp33_ASAP7_75t_L g334 ( 
.A(n_241),
.B(n_152),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_271),
.B(n_224),
.Y(n_335)
);

NOR3xp33_ASAP7_75t_L g336 ( 
.A(n_242),
.B(n_217),
.C(n_221),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_285),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_271),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_263),
.B(n_224),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_268),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_245),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_246),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_257),
.B(n_168),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_286),
.B(n_224),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_286),
.B(n_224),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_282),
.B(n_221),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_286),
.B(n_208),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_282),
.B(n_210),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_264),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_286),
.B(n_210),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_253),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_259),
.B(n_192),
.Y(n_352)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_282),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_319),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_353),
.B(n_195),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_331),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_312),
.A2(n_204),
.B1(n_215),
.B2(n_212),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_351),
.B(n_216),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_353),
.B(n_153),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_351),
.B(n_216),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_288),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_315),
.B(n_212),
.Y(n_362)
);

NOR2x2_ASAP7_75t_L g363 ( 
.A(n_340),
.B(n_11),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_329),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_298),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_349),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_307),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_315),
.B(n_154),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_319),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_348),
.B(n_313),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_306),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_331),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_348),
.B(n_222),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_307),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_308),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_320),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_319),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_296),
.B(n_155),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_326),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_300),
.B(n_204),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_329),
.B(n_204),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_352),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_L g383 ( 
.A1(n_312),
.A2(n_215),
.B1(n_229),
.B2(n_222),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_301),
.B(n_162),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_305),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_311),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_313),
.B(n_229),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_323),
.B(n_215),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_319),
.Y(n_389)
);

NOR3xp33_ASAP7_75t_SL g390 ( 
.A(n_293),
.B(n_182),
.C(n_172),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_303),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g392 ( 
.A1(n_322),
.A2(n_215),
.B1(n_193),
.B2(n_190),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_323),
.B(n_169),
.Y(n_393)
);

INVx2_ASAP7_75t_SL g394 ( 
.A(n_324),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_331),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_L g396 ( 
.A1(n_325),
.A2(n_189),
.B1(n_185),
.B2(n_183),
.Y(n_396)
);

AO22x1_ASAP7_75t_L g397 ( 
.A1(n_338),
.A2(n_180),
.B1(n_179),
.B2(n_176),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_304),
.A2(n_175),
.B1(n_174),
.B2(n_12),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_347),
.B(n_350),
.Y(n_399)
);

AND2x2_ASAP7_75t_SL g400 ( 
.A(n_337),
.B(n_13),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_330),
.Y(n_401)
);

AND2x4_ASAP7_75t_L g402 ( 
.A(n_336),
.B(n_13),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_304),
.B(n_14),
.Y(n_403)
);

CKINVDCx11_ASAP7_75t_R g404 ( 
.A(n_341),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g405 ( 
.A(n_316),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_327),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_339),
.B(n_15),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_342),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_299),
.B(n_314),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_331),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_346),
.B(n_136),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_290),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_292),
.B(n_16),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_L g414 ( 
.A1(n_336),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_414)
);

INVx5_ASAP7_75t_L g415 ( 
.A(n_294),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_321),
.B(n_302),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_R g417 ( 
.A(n_332),
.B(n_334),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_302),
.B(n_346),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_333),
.Y(n_419)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_294),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_295),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_L g422 ( 
.A1(n_318),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_L g423 ( 
.A1(n_357),
.A2(n_343),
.B1(n_291),
.B2(n_335),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_SL g424 ( 
.A1(n_400),
.A2(n_345),
.B1(n_344),
.B2(n_297),
.Y(n_424)
);

O2A1O1Ixp33_ASAP7_75t_L g425 ( 
.A1(n_364),
.A2(n_328),
.B(n_317),
.C(n_310),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_364),
.B(n_309),
.Y(n_426)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_415),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_405),
.B(n_393),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_412),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_393),
.B(n_289),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_R g431 ( 
.A(n_367),
.B(n_404),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_421),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_379),
.Y(n_433)
);

A2O1A1Ixp33_ASAP7_75t_L g434 ( 
.A1(n_370),
.A2(n_294),
.B(n_26),
.C(n_28),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_408),
.B(n_294),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_361),
.Y(n_436)
);

NAND3xp33_ASAP7_75t_L g437 ( 
.A(n_370),
.B(n_25),
.C(n_29),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_416),
.B(n_34),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_411),
.A2(n_403),
.B1(n_398),
.B2(n_388),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_L g440 ( 
.A1(n_357),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_399),
.A2(n_38),
.B(n_39),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_399),
.B(n_40),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_417),
.B(n_41),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_418),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_358),
.A2(n_45),
.B(n_49),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_403),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_374),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_382),
.B(n_135),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_385),
.B(n_53),
.Y(n_449)
);

BUFx12f_ASAP7_75t_L g450 ( 
.A(n_394),
.Y(n_450)
);

A2O1A1Ixp33_ASAP7_75t_L g451 ( 
.A1(n_409),
.A2(n_56),
.B(n_57),
.C(n_58),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_402),
.B(n_60),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_402),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_365),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_391),
.Y(n_455)
);

NAND2xp33_ASAP7_75t_L g456 ( 
.A(n_387),
.B(n_61),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_390),
.B(n_62),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_366),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_420),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_371),
.Y(n_460)
);

O2A1O1Ixp5_ASAP7_75t_L g461 ( 
.A1(n_413),
.A2(n_64),
.B(n_65),
.C(n_66),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_420),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_354),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_375),
.Y(n_464)
);

NOR3xp33_ASAP7_75t_L g465 ( 
.A(n_362),
.B(n_67),
.C(n_68),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_401),
.B(n_70),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_419),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_376),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_369),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_406),
.B(n_74),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_377),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_363),
.Y(n_472)
);

NOR3xp33_ASAP7_75t_SL g473 ( 
.A(n_368),
.B(n_77),
.C(n_78),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_358),
.A2(n_79),
.B(n_80),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_387),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_360),
.A2(n_81),
.B(n_82),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_388),
.A2(n_86),
.B1(n_88),
.B2(n_89),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_389),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_360),
.A2(n_91),
.B(n_92),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_383),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_439),
.A2(n_373),
.B(n_380),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_436),
.Y(n_482)
);

OAI21x1_ASAP7_75t_L g483 ( 
.A1(n_430),
.A2(n_373),
.B(n_356),
.Y(n_483)
);

INVx8_ASAP7_75t_L g484 ( 
.A(n_450),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_439),
.A2(n_378),
.B(n_384),
.Y(n_485)
);

AOI22x1_ASAP7_75t_L g486 ( 
.A1(n_441),
.A2(n_381),
.B1(n_386),
.B2(n_372),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_442),
.A2(n_407),
.B(n_359),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_447),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_433),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_432),
.Y(n_490)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_445),
.A2(n_395),
.B(n_356),
.Y(n_491)
);

BUFx12f_ASAP7_75t_L g492 ( 
.A(n_472),
.Y(n_492)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_431),
.Y(n_493)
);

OA21x2_ASAP7_75t_L g494 ( 
.A1(n_437),
.A2(n_392),
.B(n_414),
.Y(n_494)
);

BUFx2_ASAP7_75t_R g495 ( 
.A(n_452),
.Y(n_495)
);

INVx3_ASAP7_75t_SL g496 ( 
.A(n_435),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_429),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_454),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_427),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_467),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_427),
.Y(n_501)
);

BUFx4f_ASAP7_75t_L g502 ( 
.A(n_453),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_475),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_435),
.B(n_415),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_463),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_428),
.B(n_355),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_458),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_460),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_464),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_463),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_455),
.B(n_390),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_468),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_469),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_474),
.A2(n_372),
.B(n_410),
.Y(n_514)
);

AO21x2_ASAP7_75t_L g515 ( 
.A1(n_449),
.A2(n_354),
.B(n_410),
.Y(n_515)
);

OAI21x1_ASAP7_75t_L g516 ( 
.A1(n_476),
.A2(n_395),
.B(n_422),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_457),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_463),
.Y(n_518)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_459),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_471),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_459),
.Y(n_521)
);

OR2x6_ASAP7_75t_L g522 ( 
.A(n_448),
.B(n_354),
.Y(n_522)
);

CKINVDCx6p67_ASAP7_75t_R g523 ( 
.A(n_443),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_478),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_473),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_426),
.Y(n_526)
);

INVx6_ASAP7_75t_L g527 ( 
.A(n_462),
.Y(n_527)
);

AO21x2_ASAP7_75t_L g528 ( 
.A1(n_438),
.A2(n_397),
.B(n_415),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_506),
.A2(n_423),
.B1(n_440),
.B2(n_424),
.Y(n_529)
);

OAI22x1_ASAP7_75t_L g530 ( 
.A1(n_506),
.A2(n_526),
.B1(n_503),
.B2(n_511),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_503),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_482),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_483),
.A2(n_479),
.B(n_425),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_497),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_497),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_496),
.Y(n_536)
);

OAI21x1_ASAP7_75t_L g537 ( 
.A1(n_483),
.A2(n_461),
.B(n_477),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_498),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_502),
.B(n_465),
.Y(n_539)
);

INVx1_ASAP7_75t_SL g540 ( 
.A(n_488),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_493),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_507),
.Y(n_542)
);

CKINVDCx11_ASAP7_75t_R g543 ( 
.A(n_484),
.Y(n_543)
);

OAI22xp33_ASAP7_75t_L g544 ( 
.A1(n_525),
.A2(n_480),
.B1(n_444),
.B2(n_437),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_508),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_504),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_502),
.B(n_396),
.Y(n_547)
);

INVx8_ASAP7_75t_L g548 ( 
.A(n_484),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_494),
.A2(n_480),
.B1(n_446),
.B2(n_466),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_484),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_492),
.Y(n_551)
);

CKINVDCx11_ASAP7_75t_R g552 ( 
.A(n_492),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_490),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_490),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_509),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_489),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_L g557 ( 
.A1(n_481),
.A2(n_470),
.B(n_434),
.Y(n_557)
);

OAI21x1_ASAP7_75t_SL g558 ( 
.A1(n_485),
.A2(n_446),
.B(n_456),
.Y(n_558)
);

INVx1_ASAP7_75t_SL g559 ( 
.A(n_496),
.Y(n_559)
);

BUFx2_ASAP7_75t_R g560 ( 
.A(n_505),
.Y(n_560)
);

INVx6_ASAP7_75t_L g561 ( 
.A(n_504),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_504),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_512),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_489),
.B(n_500),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_500),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_524),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_513),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_524),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_518),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_SL g570 ( 
.A1(n_525),
.A2(n_462),
.B1(n_451),
.B2(n_415),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_515),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_571),
.Y(n_572)
);

OR2x6_ASAP7_75t_L g573 ( 
.A(n_548),
.B(n_522),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_531),
.B(n_505),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_531),
.B(n_510),
.Y(n_575)
);

AND2x4_ASAP7_75t_SL g576 ( 
.A(n_541),
.B(n_518),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_571),
.Y(n_577)
);

OR2x2_ASAP7_75t_L g578 ( 
.A(n_566),
.B(n_568),
.Y(n_578)
);

NAND3xp33_ASAP7_75t_SL g579 ( 
.A(n_529),
.B(n_517),
.C(n_487),
.Y(n_579)
);

AO31x2_ASAP7_75t_L g580 ( 
.A1(n_530),
.A2(n_513),
.A3(n_520),
.B(n_515),
.Y(n_580)
);

OR2x6_ASAP7_75t_L g581 ( 
.A(n_548),
.B(n_522),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_553),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_546),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_547),
.B(n_536),
.Y(n_584)
);

CKINVDCx16_ASAP7_75t_R g585 ( 
.A(n_550),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_553),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_536),
.B(n_510),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_540),
.B(n_495),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_L g589 ( 
.A1(n_557),
.A2(n_494),
.B(n_516),
.Y(n_589)
);

OR2x6_ASAP7_75t_L g590 ( 
.A(n_548),
.B(n_522),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_559),
.B(n_518),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_564),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_532),
.B(n_518),
.Y(n_593)
);

CKINVDCx16_ASAP7_75t_R g594 ( 
.A(n_539),
.Y(n_594)
);

CKINVDCx14_ASAP7_75t_R g595 ( 
.A(n_543),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_543),
.Y(n_596)
);

AND2x6_ASAP7_75t_L g597 ( 
.A(n_546),
.B(n_501),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g598 ( 
.A(n_569),
.Y(n_598)
);

NAND2xp33_ASAP7_75t_R g599 ( 
.A(n_551),
.B(n_494),
.Y(n_599)
);

NOR3xp33_ASAP7_75t_SL g600 ( 
.A(n_544),
.B(n_517),
.C(n_523),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_552),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_538),
.B(n_521),
.Y(n_602)
);

NOR2x1p5_ASAP7_75t_L g603 ( 
.A(n_569),
.B(n_523),
.Y(n_603)
);

BUFx8_ASAP7_75t_L g604 ( 
.A(n_542),
.Y(n_604)
);

INVx4_ASAP7_75t_L g605 ( 
.A(n_546),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_545),
.B(n_520),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_555),
.B(n_521),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_563),
.B(n_527),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_546),
.B(n_527),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_562),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_562),
.B(n_560),
.Y(n_611)
);

A2O1A1Ixp33_ASAP7_75t_L g612 ( 
.A1(n_529),
.A2(n_516),
.B(n_491),
.C(n_514),
.Y(n_612)
);

NAND2xp33_ASAP7_75t_R g613 ( 
.A(n_565),
.B(n_499),
.Y(n_613)
);

NAND3xp33_ASAP7_75t_SL g614 ( 
.A(n_549),
.B(n_519),
.C(n_527),
.Y(n_614)
);

INVxp67_ASAP7_75t_L g615 ( 
.A(n_562),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_554),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_552),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_544),
.A2(n_519),
.B1(n_486),
.B2(n_501),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_562),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_578),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_584),
.B(n_549),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_582),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_582),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_586),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_574),
.Y(n_625)
);

OR2x2_ASAP7_75t_L g626 ( 
.A(n_594),
.B(n_554),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_586),
.Y(n_627)
);

AOI221xp5_ASAP7_75t_L g628 ( 
.A1(n_579),
.A2(n_558),
.B1(n_570),
.B2(n_556),
.C(n_534),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_606),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_600),
.A2(n_519),
.B1(n_561),
.B2(n_501),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_593),
.B(n_556),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_616),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_572),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g634 ( 
.A(n_608),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_575),
.B(n_567),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_594),
.A2(n_561),
.B1(n_528),
.B2(n_499),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_602),
.B(n_567),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_572),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_577),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_589),
.B(n_577),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_592),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_591),
.B(n_535),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_607),
.B(n_535),
.Y(n_643)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_585),
.B(n_534),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_583),
.B(n_528),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_618),
.A2(n_561),
.B1(n_514),
.B2(n_491),
.Y(n_646)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_587),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_580),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_580),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_583),
.B(n_533),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_610),
.B(n_537),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_619),
.B(n_97),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_604),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_580),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_598),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_619),
.B(n_98),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_638),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_638),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_633),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_633),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_639),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_640),
.B(n_612),
.Y(n_662)
);

AND2x4_ASAP7_75t_SL g663 ( 
.A(n_642),
.B(n_573),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_640),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_625),
.B(n_611),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_647),
.B(n_576),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_621),
.B(n_588),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_621),
.B(n_596),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_639),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_620),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_624),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_635),
.B(n_614),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_632),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_634),
.B(n_644),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_627),
.B(n_604),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_655),
.B(n_595),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_622),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_629),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_622),
.Y(n_679)
);

OR2x6_ASAP7_75t_L g680 ( 
.A(n_626),
.B(n_573),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_650),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_677),
.Y(n_682)
);

NAND2x1p5_ASAP7_75t_L g683 ( 
.A(n_665),
.B(n_636),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_664),
.B(n_650),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_664),
.B(n_643),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_681),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_668),
.B(n_653),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_681),
.B(n_645),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_657),
.B(n_643),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_677),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_658),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_659),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_662),
.B(n_645),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_665),
.B(n_642),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_660),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_662),
.B(n_651),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_671),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_673),
.Y(n_698)
);

NAND4xp75_ASAP7_75t_L g699 ( 
.A(n_696),
.B(n_675),
.C(n_667),
.D(n_672),
.Y(n_699)
);

AOI32xp33_ASAP7_75t_L g700 ( 
.A1(n_696),
.A2(n_674),
.A3(n_675),
.B1(n_617),
.B2(n_670),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_693),
.B(n_672),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_697),
.Y(n_702)
);

NAND2x1p5_ASAP7_75t_L g703 ( 
.A(n_697),
.B(n_666),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_697),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_693),
.B(n_691),
.Y(n_705)
);

HB1xp67_ASAP7_75t_L g706 ( 
.A(n_684),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_692),
.Y(n_707)
);

AOI21xp33_ASAP7_75t_L g708 ( 
.A1(n_707),
.A2(n_599),
.B(n_683),
.Y(n_708)
);

OAI221xp5_ASAP7_75t_L g709 ( 
.A1(n_700),
.A2(n_683),
.B1(n_678),
.B2(n_695),
.C(n_689),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_699),
.A2(n_613),
.B1(n_694),
.B2(n_680),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_705),
.Y(n_711)
);

OAI21xp5_ASAP7_75t_SL g712 ( 
.A1(n_703),
.A2(n_687),
.B(n_686),
.Y(n_712)
);

INVx1_ASAP7_75t_SL g713 ( 
.A(n_711),
.Y(n_713)
);

OAI21xp5_ASAP7_75t_L g714 ( 
.A1(n_709),
.A2(n_701),
.B(n_704),
.Y(n_714)
);

NAND3x2_ASAP7_75t_L g715 ( 
.A(n_712),
.B(n_676),
.C(n_684),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_710),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_708),
.A2(n_694),
.B1(n_680),
.B2(n_661),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_711),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_718),
.Y(n_719)
);

NOR3x1_ASAP7_75t_L g720 ( 
.A(n_716),
.B(n_702),
.C(n_601),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_717),
.A2(n_694),
.B1(n_669),
.B2(n_631),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_713),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_722),
.Y(n_723)
);

OA22x2_ASAP7_75t_L g724 ( 
.A1(n_721),
.A2(n_714),
.B1(n_715),
.B2(n_706),
.Y(n_724)
);

OAI221xp5_ASAP7_75t_L g725 ( 
.A1(n_724),
.A2(n_719),
.B1(n_720),
.B2(n_703),
.C(n_685),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_723),
.Y(n_726)
);

AOI222xp33_ASAP7_75t_L g727 ( 
.A1(n_723),
.A2(n_628),
.B1(n_641),
.B2(n_637),
.C1(n_648),
.C2(n_654),
.Y(n_727)
);

NOR2x1_ASAP7_75t_L g728 ( 
.A(n_726),
.B(n_725),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_727),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_726),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_726),
.Y(n_731)
);

OR2x2_ASAP7_75t_L g732 ( 
.A(n_726),
.B(n_686),
.Y(n_732)
);

HB1xp67_ASAP7_75t_L g733 ( 
.A(n_726),
.Y(n_733)
);

NOR3xp33_ASAP7_75t_SL g734 ( 
.A(n_730),
.B(n_630),
.C(n_646),
.Y(n_734)
);

AOI21xp33_ASAP7_75t_SL g735 ( 
.A1(n_733),
.A2(n_590),
.B(n_581),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_731),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_732),
.Y(n_737)
);

AOI221xp5_ASAP7_75t_L g738 ( 
.A1(n_729),
.A2(n_649),
.B1(n_698),
.B2(n_688),
.C(n_682),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_728),
.Y(n_739)
);

AND2x4_ASAP7_75t_L g740 ( 
.A(n_730),
.B(n_686),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_739),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_736),
.B(n_688),
.Y(n_742)
);

NAND2xp33_ASAP7_75t_R g743 ( 
.A(n_734),
.B(n_590),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_737),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_740),
.Y(n_745)
);

BUFx2_ASAP7_75t_L g746 ( 
.A(n_738),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_735),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_744),
.B(n_741),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_SL g749 ( 
.A1(n_746),
.A2(n_581),
.B1(n_609),
.B2(n_652),
.Y(n_749)
);

HB1xp67_ASAP7_75t_L g750 ( 
.A(n_745),
.Y(n_750)
);

XNOR2x1_ASAP7_75t_L g751 ( 
.A(n_747),
.B(n_603),
.Y(n_751)
);

NOR2xp67_ASAP7_75t_L g752 ( 
.A(n_742),
.B(n_99),
.Y(n_752)
);

OAI22x1_ASAP7_75t_L g753 ( 
.A1(n_743),
.A2(n_603),
.B1(n_652),
.B2(n_656),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_744),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_744),
.B(n_656),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_741),
.A2(n_680),
.B1(n_690),
.B2(n_682),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_750),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_752),
.A2(n_649),
.B1(n_631),
.B2(n_698),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_754),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_748),
.A2(n_597),
.B1(n_690),
.B2(n_615),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_755),
.A2(n_605),
.B1(n_663),
.B2(n_679),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_751),
.B(n_605),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_SL g763 ( 
.A1(n_753),
.A2(n_597),
.B1(n_649),
.B2(n_663),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_749),
.A2(n_597),
.B1(n_632),
.B2(n_623),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_759),
.Y(n_765)
);

OA22x2_ASAP7_75t_L g766 ( 
.A1(n_757),
.A2(n_756),
.B1(n_623),
.B2(n_597),
.Y(n_766)
);

XOR2xp5_ASAP7_75t_L g767 ( 
.A(n_760),
.B(n_134),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_762),
.Y(n_768)
);

BUFx2_ASAP7_75t_L g769 ( 
.A(n_761),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_765),
.Y(n_770)
);

OAI22xp33_ASAP7_75t_L g771 ( 
.A1(n_768),
.A2(n_764),
.B1(n_763),
.B2(n_758),
.Y(n_771)
);

OAI22xp33_ASAP7_75t_L g772 ( 
.A1(n_770),
.A2(n_769),
.B1(n_766),
.B2(n_767),
.Y(n_772)
);

AOI222xp33_ASAP7_75t_L g773 ( 
.A1(n_772),
.A2(n_771),
.B1(n_102),
.B2(n_103),
.C1(n_105),
.C2(n_107),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_SL g774 ( 
.A1(n_773),
.A2(n_100),
.B1(n_109),
.B2(n_110),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_774),
.A2(n_111),
.B1(n_114),
.B2(n_115),
.Y(n_775)
);


endmodule