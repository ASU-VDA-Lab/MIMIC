module fake_jpeg_20115_n_132 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_132);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_23),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_13),
.B(n_29),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

INVx11_ASAP7_75t_SL g55 ( 
.A(n_36),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_30),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_18),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_20),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_28),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_71),
.Y(n_76)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_2),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_74),
.Y(n_83)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_62),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_71),
.A2(n_50),
.B1(n_63),
.B2(n_64),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_78),
.B1(n_84),
.B2(n_73),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_78)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_61),
.B1(n_59),
.B2(n_57),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_56),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_45),
.Y(n_91)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_89),
.Y(n_101)
);

OAI32xp33_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_48),
.A3(n_51),
.B1(n_47),
.B2(n_46),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_91),
.B(n_94),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_49),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_19),
.B(n_22),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_48),
.B1(n_49),
.B2(n_4),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_93),
.A2(n_95),
.B1(n_3),
.B2(n_4),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_52),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_21),
.B1(n_39),
.B2(n_35),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_96),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_2),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_97),
.B(n_16),
.Y(n_109)
);

BUFx2_ASAP7_75t_SL g98 ( 
.A(n_80),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_103),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_92),
.A2(n_3),
.B(n_5),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_102),
.A2(n_105),
.B(n_111),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_6),
.B(n_9),
.C(n_11),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_93),
.A2(n_6),
.B1(n_12),
.B2(n_14),
.Y(n_104)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_88),
.B(n_15),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_109),
.B(n_31),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_108),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_118),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_116),
.B(n_106),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_107),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_119),
.B(n_117),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_103),
.B(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_113),
.Y(n_123)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_122),
.A2(n_123),
.B(n_113),
.C(n_102),
.D(n_120),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_104),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_125),
.A2(n_112),
.B(n_33),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_32),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_127),
.B(n_34),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_43),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_100),
.C(n_90),
.Y(n_130)
);

BUFx24_ASAP7_75t_SL g131 ( 
.A(n_130),
.Y(n_131)
);

BUFx24_ASAP7_75t_SL g132 ( 
.A(n_131),
.Y(n_132)
);


endmodule