module fake_jpeg_13884_n_139 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_139);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_4),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_40),
.B(n_10),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_18),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_22),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_11),
.B(n_15),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_0),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_61),
.Y(n_72)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_2),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_3),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_65),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g63 ( 
.A(n_45),
.B(n_3),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_55),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_43),
.A2(n_23),
.B1(n_38),
.B2(n_37),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_44),
.B1(n_42),
.B2(n_53),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_4),
.Y(n_65)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_76),
.Y(n_94)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

NOR2x1_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_57),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_77),
.Y(n_83)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_75),
.Y(n_96)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_46),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_80),
.B(n_81),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_51),
.Y(n_81)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

OAI32xp33_ASAP7_75t_L g84 ( 
.A1(n_79),
.A2(n_63),
.A3(n_64),
.B1(n_61),
.B2(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_98),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_68),
.A2(n_74),
.B(n_71),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_90),
.B(n_12),
.C(n_14),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_88),
.B(n_91),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_55),
.B1(n_46),
.B2(n_57),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_95),
.B1(n_9),
.B2(n_10),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_70),
.A2(n_58),
.B1(n_54),
.B2(n_50),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_49),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_73),
.A2(n_54),
.B(n_47),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_7),
.C(n_8),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_5),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_97),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_21),
.B1(n_36),
.B2(n_34),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_76),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_86),
.B(n_6),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_99),
.B(n_105),
.Y(n_117)
);

AO22x1_ASAP7_75t_SL g102 ( 
.A1(n_94),
.A2(n_20),
.B1(n_33),
.B2(n_31),
.Y(n_102)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_6),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_107),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_9),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_111),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_25),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_16),
.Y(n_118)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_12),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_17),
.B1(n_24),
.B2(n_26),
.Y(n_120)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_98),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_87),
.B(n_82),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_114),
.A2(n_109),
.B(n_101),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_104),
.A2(n_85),
.B1(n_98),
.B2(n_19),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_116),
.A2(n_112),
.B1(n_100),
.B2(n_106),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_121),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_102),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_128),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_125),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_126),
.B(n_119),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_114),
.A2(n_108),
.B1(n_102),
.B2(n_30),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_130),
.A2(n_123),
.B1(n_131),
.B2(n_129),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_132),
.A2(n_133),
.B1(n_125),
.B2(n_115),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_117),
.Y(n_133)
);

OAI31xp33_ASAP7_75t_SL g135 ( 
.A1(n_134),
.A2(n_128),
.A3(n_127),
.B(n_118),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_122),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_136),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_27),
.C(n_29),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_41),
.Y(n_139)
);


endmodule