module fake_jpeg_5352_n_61 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_61);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_61;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_56;
wire n_25;
wire n_37;
wire n_43;
wire n_50;
wire n_29;
wire n_32;

INVx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx4f_ASAP7_75t_SL g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_5),
.B(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_30),
.A2(n_0),
.B1(n_35),
.B2(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_40),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_34),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_42),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_18),
.B1(n_26),
.B2(n_24),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_32),
.B(n_37),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_18),
.A2(n_24),
.B1(n_26),
.B2(n_23),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_45),
.B1(n_39),
.B2(n_43),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_49),
.A2(n_46),
.B1(n_31),
.B2(n_43),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_47),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g51 ( 
.A(n_50),
.B(n_36),
.Y(n_51)
);

XOR2x1_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_28),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_47),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_56),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_25),
.Y(n_56)
);

NOR2x1_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_29),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_44),
.C(n_27),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_58),
.Y(n_61)
);


endmodule