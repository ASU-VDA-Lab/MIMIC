module fake_jpeg_952_n_713 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_713);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_713;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_704;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_710;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_709;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_708;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_703;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_702;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_707;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_705;
wire n_665;
wire n_706;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_712;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_711;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVxp33_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_7),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_61),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_62),
.Y(n_142)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_63),
.Y(n_164)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_64),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_65),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_66),
.Y(n_169)
);

NAND2x1_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_10),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_67),
.B(n_51),
.C(n_41),
.Y(n_191)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_68),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_69),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_70),
.B(n_89),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_71),
.Y(n_220)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_72),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_73),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_74),
.Y(n_144)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_75),
.Y(n_165)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_57),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_76),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_78),
.Y(n_140)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_80),
.Y(n_225)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_81),
.Y(n_170)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_82),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_43),
.Y(n_83)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_83),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_84),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_29),
.B(n_19),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_85),
.B(n_108),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_86),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_88),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_46),
.B(n_10),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_91),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_94),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_95),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_96),
.Y(n_201)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_97),
.Y(n_183)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_98),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_99),
.Y(n_179)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_100),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_20),
.B(n_10),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_101),
.B(n_109),
.Y(n_163)
);

BUFx8_ASAP7_75t_L g102 ( 
.A(n_22),
.Y(n_102)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_102),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_103),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_50),
.Y(n_104)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_104),
.Y(n_204)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_105),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_106),
.Y(n_205)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_107),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_21),
.B(n_10),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_20),
.B(n_9),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_22),
.Y(n_110)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_110),
.Y(n_211)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_25),
.Y(n_111)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_25),
.B(n_9),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_112),
.B(n_117),
.Y(n_197)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_22),
.Y(n_113)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_45),
.Y(n_114)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_114),
.Y(n_229)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_24),
.Y(n_115)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_40),
.Y(n_116)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_116),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_28),
.B(n_12),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_31),
.Y(n_118)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_27),
.A2(n_12),
.B1(n_17),
.B2(n_16),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_119),
.A2(n_21),
.B1(n_48),
.B2(n_49),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_31),
.Y(n_121)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_28),
.Y(n_122)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_24),
.Y(n_123)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_123),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_124),
.Y(n_188)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_27),
.Y(n_125)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_125),
.Y(n_210)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_24),
.Y(n_126)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_126),
.Y(n_187)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_22),
.Y(n_127)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_127),
.Y(n_223)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_40),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_24),
.Y(n_129)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_129),
.Y(n_192)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_40),
.Y(n_130)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_130),
.Y(n_182)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_50),
.Y(n_131)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_131),
.Y(n_196)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_50),
.Y(n_132)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_132),
.Y(n_200)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_40),
.Y(n_133)
);

BUFx4f_ASAP7_75t_L g180 ( 
.A(n_133),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_67),
.B(n_47),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_149),
.B(n_203),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_76),
.B(n_33),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_151),
.B(n_162),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_65),
.A2(n_47),
.B1(n_33),
.B2(n_38),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_153),
.A2(n_186),
.B1(n_213),
.B2(n_218),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_80),
.A2(n_30),
.B1(n_58),
.B2(n_32),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_161),
.B(n_189),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_104),
.B(n_38),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_168),
.A2(n_171),
.B1(n_178),
.B2(n_181),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_103),
.A2(n_48),
.B1(n_58),
.B2(n_49),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_L g178 ( 
.A1(n_64),
.A2(n_97),
.B1(n_100),
.B2(n_72),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_66),
.A2(n_59),
.B1(n_40),
.B2(n_52),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_69),
.A2(n_53),
.B1(n_41),
.B2(n_51),
.Y(n_186)
);

OA22x2_ASAP7_75t_L g189 ( 
.A1(n_83),
.A2(n_56),
.B1(n_53),
.B2(n_52),
.Y(n_189)
);

NAND3xp33_ASAP7_75t_L g261 ( 
.A(n_191),
.B(n_8),
.C(n_1),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_120),
.B(n_34),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_193),
.B(n_199),
.Y(n_256)
);

OA22x2_ASAP7_75t_L g194 ( 
.A1(n_68),
.A2(n_56),
.B1(n_52),
.B2(n_34),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_194),
.A2(n_88),
.B1(n_121),
.B2(n_118),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_124),
.B(n_32),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_63),
.Y(n_202)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_106),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_102),
.A2(n_52),
.B1(n_30),
.B2(n_13),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_206),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_114),
.B(n_52),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_207),
.B(n_208),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_62),
.B(n_102),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_71),
.A2(n_93),
.B1(n_92),
.B2(n_74),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_61),
.B(n_12),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_214),
.B(n_179),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_62),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_215),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_84),
.A2(n_12),
.B1(n_17),
.B2(n_16),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_73),
.Y(n_219)
);

BUFx4f_ASAP7_75t_L g263 ( 
.A(n_219),
.Y(n_263)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_75),
.Y(n_221)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_81),
.Y(n_222)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_86),
.A2(n_6),
.B1(n_15),
.B2(n_14),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_227),
.A2(n_228),
.B1(n_3),
.B2(n_4),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_95),
.A2(n_18),
.B1(n_14),
.B2(n_13),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_133),
.Y(n_230)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_230),
.Y(n_258)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_159),
.Y(n_233)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_233),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_234),
.B(n_279),
.Y(n_337)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_155),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_235),
.Y(n_315)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_175),
.Y(n_237)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_237),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_145),
.B(n_113),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_238),
.B(n_240),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_L g239 ( 
.A1(n_206),
.A2(n_96),
.B1(n_130),
.B2(n_116),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_239),
.A2(n_265),
.B1(n_282),
.B2(n_176),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_145),
.B(n_8),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_204),
.Y(n_241)
);

INVx4_ASAP7_75t_SL g318 ( 
.A(n_241),
.Y(n_318)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_242),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_215),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_243),
.B(n_273),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_155),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_244),
.Y(n_347)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_187),
.Y(n_245)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_245),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_148),
.Y(n_246)
);

BUFx4f_ASAP7_75t_L g329 ( 
.A(n_246),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_247),
.A2(n_259),
.B1(n_308),
.B2(n_309),
.Y(n_340)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_192),
.Y(n_249)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_249),
.Y(n_371)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_169),
.Y(n_250)
);

INVx8_ASAP7_75t_L g359 ( 
.A(n_250),
.Y(n_359)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g366 ( 
.A(n_251),
.Y(n_366)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_169),
.Y(n_252)
);

INVx5_ASAP7_75t_L g363 ( 
.A(n_252),
.Y(n_363)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_253),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_217),
.Y(n_254)
);

INVx6_ASAP7_75t_L g338 ( 
.A(n_254),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_208),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g374 ( 
.A(n_255),
.Y(n_374)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_217),
.Y(n_257)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_257),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_157),
.A2(n_8),
.B1(n_18),
.B2(n_2),
.Y(n_259)
);

OAI21xp33_ASAP7_75t_L g328 ( 
.A1(n_261),
.A2(n_268),
.B(n_271),
.Y(n_328)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_138),
.Y(n_262)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_262),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_180),
.Y(n_264)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_264),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_171),
.A2(n_178),
.B1(n_213),
.B2(n_194),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_147),
.B(n_4),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_142),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g326 ( 
.A(n_269),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_219),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_270),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_163),
.B(n_0),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_167),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_272),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_136),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_183),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_274),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_163),
.B(n_1),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_276),
.B(n_307),
.Y(n_341)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_164),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_277),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_139),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_278),
.B(n_286),
.Y(n_322)
);

NAND2xp33_ASAP7_75t_SL g279 ( 
.A(n_210),
.B(n_1),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_195),
.Y(n_280)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_280),
.Y(n_333)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_196),
.Y(n_281)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_281),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_194),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_220),
.Y(n_283)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_283),
.Y(n_370)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_165),
.Y(n_284)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_284),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_220),
.Y(n_285)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_285),
.Y(n_376)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_170),
.Y(n_286)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_158),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_287),
.Y(n_372)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_200),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_288),
.B(n_289),
.Y(n_325)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_223),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_141),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_290),
.B(n_292),
.Y(n_336)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_143),
.Y(n_291)
);

INVx13_ASAP7_75t_L g358 ( 
.A(n_291),
.Y(n_358)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_152),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_172),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_293),
.B(n_294),
.Y(n_342)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_174),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_295),
.B(n_296),
.Y(n_348)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_184),
.Y(n_296)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_182),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_298),
.B(n_299),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_197),
.B(n_3),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_198),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_300),
.B(n_301),
.Y(n_354)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_182),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_139),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_302),
.B(n_304),
.Y(n_355)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_135),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_216),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_305),
.B(n_306),
.Y(n_356)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_137),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_197),
.B(n_140),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_211),
.A2(n_3),
.B1(n_4),
.B2(n_156),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_173),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_310),
.B(n_313),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_144),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_311),
.A2(n_312),
.B1(n_314),
.B2(n_209),
.Y(n_346)
);

INVx8_ASAP7_75t_L g312 ( 
.A(n_144),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_150),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_176),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_267),
.A2(n_189),
.B(n_177),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_321),
.A2(n_246),
.B(n_259),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_303),
.A2(n_189),
.B1(n_209),
.B2(n_188),
.Y(n_323)
);

OAI22xp33_ASAP7_75t_SL g418 ( 
.A1(n_323),
.A2(n_327),
.B1(n_241),
.B2(n_298),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_260),
.B(n_146),
.C(n_212),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_324),
.B(n_304),
.C(n_242),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_256),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_232),
.B(n_229),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_330),
.B(n_349),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_282),
.A2(n_185),
.B(n_205),
.Y(n_332)
);

NOR3xp33_ASAP7_75t_L g424 ( 
.A(n_332),
.B(n_353),
.C(n_317),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_339),
.A2(n_352),
.B1(n_368),
.B2(n_239),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_346),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_268),
.B(n_224),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_299),
.B(n_224),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_351),
.B(n_364),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_247),
.A2(n_154),
.B1(n_190),
.B2(n_201),
.Y(n_352)
);

NAND2xp33_ASAP7_75t_SL g353 ( 
.A(n_270),
.B(n_173),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_353),
.B(n_297),
.Y(n_388)
);

O2A1O1Ixp33_ASAP7_75t_L g364 ( 
.A1(n_275),
.A2(n_185),
.B(n_212),
.C(n_158),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_263),
.A2(n_180),
.B1(n_264),
.B2(n_291),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g426 ( 
.A1(n_365),
.A2(n_318),
.B1(n_366),
.B2(n_317),
.Y(n_426)
);

OAI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_309),
.A2(n_154),
.B1(n_134),
.B2(n_160),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_231),
.B(n_134),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_369),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_261),
.B(n_190),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_377),
.B(n_287),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_378),
.A2(n_390),
.B1(n_406),
.B2(n_407),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_342),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_379),
.B(n_380),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_356),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_336),
.Y(n_381)
);

CKINVDCx14_ASAP7_75t_R g469 ( 
.A(n_381),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_331),
.Y(n_382)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_382),
.Y(n_430)
);

NAND3xp33_ASAP7_75t_L g383 ( 
.A(n_357),
.B(n_341),
.C(n_348),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_383),
.B(n_408),
.Y(n_429)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_331),
.Y(n_384)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_384),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_357),
.B(n_319),
.Y(n_385)
);

CKINVDCx14_ASAP7_75t_R g444 ( 
.A(n_385),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_339),
.A2(n_321),
.B1(n_337),
.B2(n_330),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_386),
.A2(n_393),
.B1(n_398),
.B2(n_318),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_324),
.B(n_258),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_387),
.B(n_403),
.C(n_420),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_388),
.B(n_424),
.Y(n_462)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_320),
.Y(n_389)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_389),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_337),
.A2(n_160),
.B1(n_166),
.B2(n_201),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_341),
.B(n_349),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_391),
.B(n_395),
.Y(n_443)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_329),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_392),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_337),
.A2(n_312),
.B1(n_311),
.B2(n_314),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_394),
.A2(n_372),
.B(n_375),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_351),
.B(n_248),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_374),
.B(n_236),
.Y(n_396)
);

CKINVDCx14_ASAP7_75t_R g454 ( 
.A(n_396),
.Y(n_454)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_329),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_397),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_352),
.A2(n_166),
.B1(n_285),
.B2(n_283),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_329),
.Y(n_399)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_399),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_320),
.B(n_297),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_401),
.B(n_416),
.Y(n_445)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_355),
.Y(n_402)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_402),
.Y(n_451)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_344),
.Y(n_404)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_404),
.Y(n_456)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_344),
.Y(n_405)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_405),
.Y(n_458)
);

OAI22x1_ASAP7_75t_SL g406 ( 
.A1(n_340),
.A2(n_364),
.B1(n_377),
.B2(n_332),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_350),
.A2(n_250),
.B1(n_235),
.B2(n_257),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_345),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_345),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_409),
.B(n_411),
.Y(n_450)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_366),
.Y(n_410)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_410),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_322),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_318),
.Y(n_414)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_414),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_361),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_328),
.A2(n_252),
.B1(n_244),
.B2(n_254),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_417),
.A2(n_418),
.B1(n_422),
.B2(n_376),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_419),
.B(n_421),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_325),
.B(n_263),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_354),
.B(n_301),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_373),
.A2(n_4),
.B1(n_362),
.B2(n_376),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_329),
.Y(n_423)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_423),
.Y(n_464)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_366),
.Y(n_425)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_425),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_SL g441 ( 
.A1(n_426),
.A2(n_372),
.B1(n_326),
.B2(n_316),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_358),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_427),
.Y(n_440)
);

AND2x2_ASAP7_75t_SL g431 ( 
.A(n_386),
.B(n_373),
.Y(n_431)
);

CKINVDCx14_ASAP7_75t_R g502 ( 
.A(n_431),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_387),
.B(n_333),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_433),
.B(n_434),
.C(n_453),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_403),
.B(n_333),
.C(n_375),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_436),
.A2(n_410),
.B(n_423),
.Y(n_492)
);

OAI21xp33_ASAP7_75t_SL g505 ( 
.A1(n_439),
.A2(n_441),
.B(n_460),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_394),
.A2(n_316),
.B(n_358),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_446),
.A2(n_452),
.B(n_421),
.Y(n_481)
);

NAND2x1_ASAP7_75t_L g447 ( 
.A(n_394),
.B(n_388),
.Y(n_447)
);

OAI21xp33_ASAP7_75t_L g494 ( 
.A1(n_447),
.A2(n_422),
.B(n_399),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_413),
.A2(n_358),
.B(n_334),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_391),
.B(n_360),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_412),
.B(n_371),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_457),
.B(n_463),
.C(n_465),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_SL g461 ( 
.A1(n_400),
.A2(n_390),
.B1(n_388),
.B2(n_417),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_461),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_412),
.B(n_371),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_402),
.B(n_360),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_401),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_466),
.B(n_381),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_380),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_470),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_428),
.B(n_420),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_471),
.B(n_434),
.C(n_465),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_437),
.A2(n_378),
.B1(n_419),
.B2(n_413),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_472),
.A2(n_474),
.B1(n_477),
.B2(n_493),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_468),
.B(n_385),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_473),
.B(n_486),
.Y(n_523)
);

OAI22x1_ASAP7_75t_SL g474 ( 
.A1(n_437),
.A2(n_406),
.B1(n_393),
.B2(n_398),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_431),
.A2(n_379),
.B1(n_411),
.B2(n_395),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_432),
.Y(n_478)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_478),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_445),
.B(n_416),
.Y(n_479)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_479),
.Y(n_515)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_432),
.Y(n_480)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_480),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_481),
.A2(n_483),
.B(n_492),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_466),
.B(n_415),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_482),
.B(n_491),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_447),
.A2(n_396),
.B(n_408),
.Y(n_483)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_484),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_428),
.B(n_389),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_485),
.B(n_488),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_451),
.B(n_409),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_469),
.B(n_334),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_487),
.B(n_496),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_433),
.B(n_404),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_446),
.A2(n_407),
.B1(n_405),
.B2(n_384),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_489),
.A2(n_495),
.B1(n_440),
.B2(n_467),
.Y(n_513)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_435),
.Y(n_490)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_490),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_445),
.B(n_425),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_431),
.A2(n_370),
.B1(n_362),
.B2(n_315),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_494),
.A2(n_442),
.B(n_448),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_439),
.A2(n_370),
.B1(n_338),
.B2(n_414),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_435),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_456),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_497),
.B(n_498),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_454),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_447),
.A2(n_427),
.B(n_414),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_499),
.A2(n_462),
.B(n_455),
.Y(n_518)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_456),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_500),
.B(n_501),
.Y(n_522)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_458),
.Y(n_501)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_458),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_503),
.B(n_504),
.Y(n_529)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_459),
.Y(n_504)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_459),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_506),
.B(n_508),
.Y(n_530)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_430),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_491),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_509),
.B(n_533),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_502),
.A2(n_436),
.B1(n_460),
.B2(n_452),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_510),
.A2(n_517),
.B1(n_527),
.B2(n_535),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_512),
.B(n_526),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_513),
.B(n_531),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_481),
.A2(n_455),
.B1(n_444),
.B2(n_443),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_SL g552 ( 
.A1(n_518),
.A2(n_519),
.B(n_520),
.Y(n_552)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_492),
.A2(n_462),
.B(n_450),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_483),
.A2(n_462),
.B(n_443),
.Y(n_520)
);

AOI21xp33_ASAP7_75t_L g524 ( 
.A1(n_507),
.A2(n_429),
.B(n_453),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_524),
.A2(n_532),
.B(n_495),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_SL g525 ( 
.A(n_471),
.B(n_463),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_SL g554 ( 
.A(n_525),
.B(n_543),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_485),
.B(n_457),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_479),
.A2(n_430),
.B1(n_467),
.B2(n_442),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_507),
.A2(n_448),
.B(n_438),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_484),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_474),
.A2(n_440),
.B1(n_464),
.B2(n_449),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_475),
.B(n_367),
.C(n_335),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_537),
.B(n_476),
.C(n_475),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_489),
.A2(n_438),
.B1(n_449),
.B2(n_464),
.Y(n_540)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_540),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_482),
.B(n_397),
.Y(n_541)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_541),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_SL g543 ( 
.A(n_476),
.B(n_367),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_472),
.A2(n_392),
.B1(n_363),
.B2(n_315),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_544),
.B(n_493),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_498),
.B(n_363),
.Y(n_545)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_545),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_508),
.B(n_315),
.Y(n_546)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_546),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_522),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_548),
.B(n_549),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_522),
.Y(n_549)
);

CKINVDCx16_ASAP7_75t_R g550 ( 
.A(n_542),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_550),
.B(n_569),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_551),
.B(n_562),
.C(n_574),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_536),
.B(n_473),
.Y(n_556)
);

INVxp33_ASAP7_75t_SL g607 ( 
.A(n_556),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_529),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g587 ( 
.A1(n_558),
.A2(n_582),
.B1(n_515),
.B2(n_534),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_533),
.B(n_477),
.Y(n_560)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_560),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_512),
.B(n_488),
.C(n_499),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_SL g563 ( 
.A(n_525),
.B(n_505),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_563),
.B(n_566),
.Y(n_595)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_565),
.Y(n_591)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_538),
.B(n_504),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_538),
.B(n_506),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_567),
.B(n_516),
.Y(n_593)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_542),
.Y(n_568)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_568),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_SL g569 ( 
.A(n_523),
.B(n_480),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_534),
.B(n_343),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_570),
.B(n_577),
.Y(n_598)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_543),
.B(n_490),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_571),
.B(n_524),
.Y(n_605)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_545),
.Y(n_572)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_572),
.Y(n_608)
);

OAI21xp5_ASAP7_75t_L g601 ( 
.A1(n_573),
.A2(n_531),
.B(n_532),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_537),
.B(n_478),
.C(n_501),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_543),
.B(n_503),
.C(n_500),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_575),
.B(n_581),
.C(n_520),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_SL g577 ( 
.A(n_523),
.B(n_497),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_509),
.B(n_496),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_579),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_516),
.B(n_338),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_580),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_526),
.B(n_335),
.C(n_343),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_529),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g584 ( 
.A1(n_552),
.A2(n_514),
.B(n_576),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_SL g630 ( 
.A1(n_584),
.A2(n_596),
.B(n_601),
.Y(n_630)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_587),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_553),
.A2(n_539),
.B1(n_535),
.B2(n_517),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_588),
.A2(n_600),
.B1(n_602),
.B2(n_611),
.Y(n_633)
);

XNOR2xp5_ASAP7_75t_L g617 ( 
.A(n_589),
.B(n_593),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_551),
.B(n_519),
.C(n_518),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_590),
.B(n_597),
.C(n_606),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_552),
.A2(n_514),
.B(n_510),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_564),
.B(n_540),
.C(n_527),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_559),
.A2(n_539),
.B1(n_515),
.B2(n_568),
.Y(n_599)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_599),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_SL g600 ( 
.A1(n_559),
.A2(n_553),
.B1(n_573),
.B2(n_582),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_548),
.A2(n_513),
.B1(n_541),
.B2(n_528),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g604 ( 
.A(n_564),
.B(n_566),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_604),
.B(n_567),
.Y(n_622)
);

XNOR2xp5_ASAP7_75t_SL g613 ( 
.A(n_605),
.B(n_563),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_562),
.B(n_530),
.C(n_544),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_574),
.B(n_530),
.C(n_528),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_610),
.B(n_571),
.C(n_581),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_549),
.A2(n_511),
.B1(n_521),
.B2(n_547),
.Y(n_611)
);

XOR2xp5_ASAP7_75t_L g649 ( 
.A(n_613),
.B(n_605),
.Y(n_649)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_592),
.Y(n_614)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_614),
.Y(n_650)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_592),
.Y(n_615)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_615),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_600),
.B(n_576),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_616),
.B(n_625),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_607),
.B(n_578),
.Y(n_618)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_618),
.Y(n_657)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_585),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_619),
.B(n_624),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_SL g620 ( 
.A1(n_594),
.A2(n_576),
.B1(n_558),
.B2(n_578),
.Y(n_620)
);

XNOR2xp5_ASAP7_75t_L g641 ( 
.A(n_620),
.B(n_622),
.Y(n_641)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_609),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_621),
.B(n_623),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_597),
.B(n_575),
.Y(n_623)
);

CKINVDCx16_ASAP7_75t_R g624 ( 
.A(n_598),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_611),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_609),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_626),
.B(n_631),
.Y(n_647)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_602),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_628),
.B(n_591),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g651 ( 
.A(n_629),
.Y(n_651)
);

INVxp67_ASAP7_75t_L g631 ( 
.A(n_610),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_586),
.B(n_579),
.Y(n_632)
);

XNOR2xp5_ASAP7_75t_L g642 ( 
.A(n_632),
.B(n_635),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_591),
.A2(n_572),
.B1(n_557),
.B2(n_555),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_SL g637 ( 
.A1(n_634),
.A2(n_608),
.B1(n_603),
.B2(n_561),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_SL g635 ( 
.A1(n_584),
.A2(n_557),
.B(n_555),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_637),
.A2(n_654),
.B1(n_511),
.B2(n_547),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_639),
.Y(n_670)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_617),
.B(n_583),
.C(n_631),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_640),
.B(n_644),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_617),
.B(n_583),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_636),
.A2(n_608),
.B1(n_601),
.B2(n_588),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g665 ( 
.A1(n_645),
.A2(n_655),
.B1(n_647),
.B2(n_657),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_612),
.B(n_606),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_646),
.B(n_648),
.Y(n_674)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_627),
.B(n_604),
.C(n_589),
.Y(n_648)
);

XOR2xp5_ASAP7_75t_L g671 ( 
.A(n_649),
.B(n_554),
.Y(n_671)
);

OAI22xp5_ASAP7_75t_SL g654 ( 
.A1(n_633),
.A2(n_596),
.B1(n_561),
.B2(n_580),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_626),
.A2(n_590),
.B1(n_593),
.B2(n_595),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_627),
.B(n_521),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_SL g660 ( 
.A1(n_656),
.A2(n_618),
.B(n_632),
.Y(n_660)
);

XNOR2xp5_ASAP7_75t_L g658 ( 
.A(n_648),
.B(n_620),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_658),
.B(n_659),
.Y(n_680)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_640),
.B(n_629),
.C(n_633),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_660),
.B(n_661),
.Y(n_684)
);

MAJIxp5_ASAP7_75t_L g661 ( 
.A(n_651),
.B(n_625),
.C(n_622),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_SL g662 ( 
.A1(n_653),
.A2(n_630),
.B(n_635),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_662),
.A2(n_664),
.B(n_666),
.Y(n_681)
);

MAJIxp5_ASAP7_75t_L g663 ( 
.A(n_655),
.B(n_616),
.C(n_630),
.Y(n_663)
);

MAJIxp5_ASAP7_75t_L g677 ( 
.A(n_663),
.B(n_673),
.C(n_641),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_L g664 ( 
.A1(n_647),
.A2(n_616),
.B(n_634),
.Y(n_664)
);

XNOR2xp5_ASAP7_75t_L g676 ( 
.A(n_665),
.B(n_667),
.Y(n_676)
);

OAI21xp5_ASAP7_75t_SL g666 ( 
.A1(n_638),
.A2(n_613),
.B(n_546),
.Y(n_666)
);

XOR2xp5_ASAP7_75t_SL g667 ( 
.A(n_649),
.B(n_595),
.Y(n_667)
);

XNOR2xp5_ASAP7_75t_L g683 ( 
.A(n_669),
.B(n_642),
.Y(n_683)
);

XOR2xp5_ASAP7_75t_L g682 ( 
.A(n_671),
.B(n_642),
.Y(n_682)
);

AOI211xp5_ASAP7_75t_L g672 ( 
.A1(n_637),
.A2(n_554),
.B(n_347),
.C(n_326),
.Y(n_672)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_672),
.A2(n_650),
.B(n_652),
.Y(n_686)
);

MAJIxp5_ASAP7_75t_L g673 ( 
.A(n_641),
.B(n_347),
.C(n_359),
.Y(n_673)
);

INVx6_ASAP7_75t_L g675 ( 
.A(n_674),
.Y(n_675)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_675),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_677),
.B(n_679),
.Y(n_693)
);

MAJIxp5_ASAP7_75t_L g678 ( 
.A(n_659),
.B(n_643),
.C(n_654),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_678),
.B(n_683),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_SL g679 ( 
.A(n_668),
.B(n_670),
.Y(n_679)
);

XNOR2xp5_ASAP7_75t_L g689 ( 
.A(n_682),
.B(n_664),
.Y(n_689)
);

OAI21xp5_ASAP7_75t_L g685 ( 
.A1(n_658),
.A2(n_645),
.B(n_643),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_685),
.B(n_686),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g687 ( 
.A1(n_663),
.A2(n_338),
.B(n_359),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_687),
.B(n_673),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_SL g688 ( 
.A(n_684),
.B(n_661),
.Y(n_688)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_688),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_689),
.B(n_694),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_675),
.B(n_669),
.Y(n_691)
);

NOR3xp33_ASAP7_75t_L g699 ( 
.A(n_691),
.B(n_695),
.C(n_681),
.Y(n_699)
);

XNOR2xp5_ASAP7_75t_L g694 ( 
.A(n_682),
.B(n_667),
.Y(n_694)
);

NOR2x1_ASAP7_75t_L g695 ( 
.A(n_683),
.B(n_672),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_SL g700 ( 
.A(n_697),
.B(n_680),
.Y(n_700)
);

AO21x1_ASAP7_75t_L g705 ( 
.A1(n_699),
.A2(n_700),
.B(n_702),
.Y(n_705)
);

OAI21xp5_ASAP7_75t_L g701 ( 
.A1(n_692),
.A2(n_676),
.B(n_678),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_SL g706 ( 
.A1(n_701),
.A2(n_695),
.B(n_691),
.Y(n_706)
);

BUFx24_ASAP7_75t_SL g702 ( 
.A(n_696),
.Y(n_702)
);

MAJIxp5_ASAP7_75t_L g704 ( 
.A(n_703),
.B(n_693),
.C(n_690),
.Y(n_704)
);

INVxp67_ASAP7_75t_L g708 ( 
.A(n_704),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_SL g707 ( 
.A1(n_706),
.A2(n_698),
.B(n_705),
.Y(n_707)
);

INVxp67_ASAP7_75t_L g709 ( 
.A(n_707),
.Y(n_709)
);

AOI221xp5_ASAP7_75t_L g710 ( 
.A1(n_709),
.A2(n_708),
.B1(n_677),
.B2(n_676),
.C(n_671),
.Y(n_710)
);

OAI21xp5_ASAP7_75t_SL g711 ( 
.A1(n_710),
.A2(n_347),
.B(n_359),
.Y(n_711)
);

MAJIxp5_ASAP7_75t_L g712 ( 
.A(n_711),
.B(n_326),
.C(n_696),
.Y(n_712)
);

INVxp67_ASAP7_75t_L g713 ( 
.A(n_712),
.Y(n_713)
);


endmodule