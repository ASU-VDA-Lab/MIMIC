module fake_jpeg_13712_n_246 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_246);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_246;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_43),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_24),
.B(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_59),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_19),
.B(n_0),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_17),
.B(n_0),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_65),
.Y(n_96)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_24),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_33),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_67),
.B(n_69),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_33),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_21),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_71),
.B(n_86),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_43),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_75),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_44),
.B(n_37),
.Y(n_75)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_37),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_79),
.B(n_99),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_22),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_41),
.A2(n_39),
.B1(n_18),
.B2(n_36),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_88),
.A2(n_90),
.B1(n_94),
.B2(n_102),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_42),
.A2(n_18),
.B1(n_36),
.B2(n_26),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_46),
.A2(n_50),
.B1(n_51),
.B2(n_48),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_29),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_56),
.A2(n_38),
.B1(n_35),
.B2(n_20),
.Y(n_102)
);

AO22x1_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_98),
.B1(n_88),
.B2(n_43),
.Y(n_103)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_106),
.Y(n_160)
);

INVx3_ASAP7_75t_SL g109 ( 
.A(n_80),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_112),
.Y(n_154)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_99),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_124),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_55),
.Y(n_112)
);

INVx4_ASAP7_75t_SL g113 ( 
.A(n_92),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_113),
.B(n_114),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_26),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_34),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_115),
.B(n_133),
.Y(n_162)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_22),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_117),
.B(n_122),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_73),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_119),
.A2(n_101),
.B1(n_95),
.B2(n_85),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_93),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_120),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_20),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_71),
.B(n_15),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_123),
.B(n_127),
.Y(n_147)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_0),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_130),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_70),
.B(n_15),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_97),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_101),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_66),
.B(n_13),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_129),
.B(n_132),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_84),
.B(n_1),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_131),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

NOR2x1_ASAP7_75t_L g133 ( 
.A(n_68),
.B(n_74),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_133),
.B(n_103),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_81),
.B(n_10),
.Y(n_134)
);

NAND3xp33_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_2),
.C(n_5),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_74),
.C(n_9),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_162),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_138),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_143),
.B(n_161),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_125),
.A2(n_95),
.B1(n_85),
.B2(n_84),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_145),
.A2(n_146),
.B1(n_151),
.B2(n_152),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_76),
.B1(n_5),
.B2(n_6),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_121),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_149),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_76),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_157),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_103),
.A2(n_7),
.B1(n_8),
.B2(n_130),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_108),
.A2(n_7),
.B1(n_8),
.B2(n_112),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_114),
.B(n_107),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_115),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_104),
.B(n_106),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_160),
.Y(n_164)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_160),
.Y(n_166)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_166),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_168),
.B(n_179),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_153),
.A2(n_136),
.B(n_149),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_169),
.A2(n_182),
.B(n_120),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_115),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_183),
.Y(n_187)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_148),
.B(n_142),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_174),
.B(n_175),
.Y(n_198)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_135),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_177),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_140),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_108),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_178),
.B(n_180),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_159),
.B(n_113),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_128),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_136),
.A2(n_153),
.B(n_154),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_156),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_110),
.Y(n_193)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_120),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_182),
.A2(n_169),
.B(n_185),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_188),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_174),
.A2(n_151),
.B1(n_145),
.B2(n_154),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_189),
.A2(n_192),
.B1(n_179),
.B2(n_173),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_163),
.A2(n_158),
.B(n_162),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_191),
.B(n_202),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_158),
.B1(n_137),
.B2(n_109),
.Y(n_192)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_193),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_158),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_195),
.B(n_203),
.Y(n_216)
);

OAI32xp33_ASAP7_75t_L g215 ( 
.A1(n_200),
.A2(n_164),
.A3(n_166),
.B1(n_167),
.B2(n_173),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_177),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_163),
.A2(n_113),
.B(n_124),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_170),
.B(n_155),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_181),
.C(n_172),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_209),
.C(n_210),
.Y(n_220)
);

NOR3xp33_ASAP7_75t_SL g207 ( 
.A(n_199),
.B(n_168),
.C(n_165),
.Y(n_207)
);

AOI322xp5_ASAP7_75t_L g222 ( 
.A1(n_207),
.A2(n_197),
.A3(n_186),
.B1(n_198),
.B2(n_199),
.C1(n_196),
.C2(n_203),
.Y(n_222)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_208),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_181),
.C(n_175),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_183),
.C(n_184),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_190),
.Y(n_211)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_211),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_212),
.A2(n_200),
.B(n_187),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_214),
.A2(n_215),
.B1(n_201),
.B2(n_213),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_210),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_219),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_204),
.Y(n_219)
);

AOI31xp67_ASAP7_75t_L g230 ( 
.A1(n_222),
.A2(n_207),
.A3(n_197),
.B(n_216),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_225),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_224),
.A2(n_225),
.B(n_213),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_202),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_209),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_228),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_227),
.B(n_229),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_206),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_214),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_232),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_231),
.A2(n_223),
.B1(n_224),
.B2(n_189),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_234),
.A2(n_194),
.B(n_171),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_228),
.A2(n_221),
.B1(n_217),
.B2(n_194),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_236),
.B(n_221),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_238),
.A2(n_240),
.B(n_237),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_217),
.Y(n_239)
);

AOI21x1_ASAP7_75t_L g243 ( 
.A1(n_239),
.A2(n_241),
.B(n_105),
.Y(n_243)
);

AOI31xp67_ASAP7_75t_SL g241 ( 
.A1(n_234),
.A2(n_226),
.A3(n_155),
.B(n_116),
.Y(n_241)
);

NOR3xp33_ASAP7_75t_SL g244 ( 
.A(n_242),
.B(n_243),
.C(n_119),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_244),
.A2(n_109),
.B1(n_105),
.B2(n_233),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_245),
.B(n_233),
.Y(n_246)
);


endmodule