module fake_jpeg_23586_n_231 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_231);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_56;
wire n_131;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_41),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_31),
.B(n_1),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_33),
.A2(n_25),
.B1(n_31),
.B2(n_28),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_28),
.B1(n_21),
.B2(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_44),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_31),
.B1(n_25),
.B2(n_30),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_47),
.A2(n_48),
.B1(n_19),
.B2(n_22),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_25),
.B1(n_30),
.B2(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_35),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_16),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_24),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_39),
.Y(n_83)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_58),
.B(n_59),
.Y(n_112)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_62),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_61),
.A2(n_71),
.B1(n_78),
.B2(n_81),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_49),
.B(n_26),
.Y(n_62)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_64),
.B(n_65),
.Y(n_113)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_68),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_46),
.Y(n_68)
);

O2A1O1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_48),
.A2(n_40),
.B(n_33),
.C(n_29),
.Y(n_69)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_73),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_45),
.A2(n_33),
.B1(n_38),
.B2(n_37),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_16),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_72),
.B(n_75),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_50),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_77),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_18),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g77 ( 
.A(n_52),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_29),
.B1(n_24),
.B2(n_26),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_56),
.B(n_18),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_83),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_91),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_56),
.A2(n_37),
.B1(n_40),
.B2(n_23),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_85),
.B1(n_90),
.B2(n_36),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_53),
.A2(n_23),
.B1(n_22),
.B2(n_19),
.Y(n_85)
);

FAx1_ASAP7_75t_SL g98 ( 
.A(n_87),
.B(n_36),
.CI(n_54),
.CON(n_98),
.SN(n_98)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_44),
.A2(n_19),
.B1(n_2),
.B2(n_3),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_17),
.B(n_4),
.Y(n_108)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_23),
.Y(n_91)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_94),
.B(n_103),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_96),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_102),
.B1(n_108),
.B2(n_90),
.Y(n_124)
);

FAx1_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_39),
.CI(n_36),
.CON(n_101),
.SN(n_101)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_101),
.B(n_89),
.Y(n_137)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_10),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_64),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_110),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_69),
.A2(n_88),
.B(n_81),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_3),
.B(n_5),
.Y(n_138)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_118),
.B(n_119),
.Y(n_151)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_125),
.Y(n_143)
);

AO21x1_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_115),
.B(n_101),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_122),
.A2(n_136),
.B(n_138),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_137),
.B1(n_94),
.B2(n_114),
.Y(n_153)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_39),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_134),
.Y(n_156)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_85),
.B1(n_86),
.B2(n_84),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_114),
.B1(n_100),
.B2(n_86),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_111),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_133),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_117),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_39),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_93),
.C(n_117),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_93),
.C(n_92),
.Y(n_145)
);

OAI21x1_ASAP7_75t_SL g136 ( 
.A1(n_108),
.A2(n_68),
.B(n_4),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_92),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_139),
.A2(n_94),
.B1(n_103),
.B2(n_110),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_141),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_142),
.B(n_144),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_146),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_101),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_122),
.A2(n_97),
.B1(n_98),
.B2(n_104),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_147),
.A2(n_154),
.B1(n_158),
.B2(n_161),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_98),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_159),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

INVxp67_ASAP7_75t_SL g175 ( 
.A(n_152),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_153),
.Y(n_168)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_100),
.B1(n_116),
.B2(n_82),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_125),
.A2(n_116),
.B(n_8),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_118),
.A2(n_107),
.B1(n_8),
.B2(n_6),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_160),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_121),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_143),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_165),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_152),
.A2(n_140),
.B1(n_119),
.B2(n_129),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_166),
.A2(n_154),
.B(n_139),
.Y(n_193)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_177),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_157),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_170),
.Y(n_184)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_162),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_172),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_159),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_174),
.B(n_148),
.Y(n_183)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_150),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_182),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_146),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_183),
.A2(n_191),
.B1(n_193),
.B2(n_166),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_156),
.C(n_145),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_190),
.C(n_193),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_156),
.C(n_147),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_176),
.A2(n_161),
.B1(n_140),
.B2(n_148),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_164),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_204),
.C(n_190),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_196),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_197),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_188),
.A2(n_176),
.B1(n_168),
.B2(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_198),
.Y(n_209)
);

MAJx2_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_174),
.C(n_121),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_202),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_191),
.A2(n_169),
.B1(n_177),
.B2(n_178),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_201),
.A2(n_187),
.B1(n_173),
.B2(n_181),
.Y(n_210)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_186),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_170),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_164),
.C(n_167),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_195),
.C(n_200),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_204),
.B(n_184),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_208),
.B(n_194),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_198),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_199),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_216),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_210),
.B(n_165),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_214),
.B(n_211),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_217),
.Y(n_220)
);

OAI221xp5_ASAP7_75t_L g218 ( 
.A1(n_212),
.A2(n_172),
.B1(n_128),
.B2(n_120),
.C(n_195),
.Y(n_218)
);

NOR2xp67_ASAP7_75t_SL g222 ( 
.A(n_218),
.B(n_207),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_219),
.B(n_222),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_205),
.C(n_206),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_223),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_180),
.Y(n_224)
);

NOR2x1_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_209),
.Y(n_226)
);

AOI322xp5_ASAP7_75t_L g228 ( 
.A1(n_226),
.A2(n_225),
.A3(n_126),
.B1(n_123),
.B2(n_131),
.C1(n_13),
.C2(n_11),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_227),
.C(n_123),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_229),
.A2(n_13),
.B(n_14),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_6),
.Y(n_231)
);


endmodule