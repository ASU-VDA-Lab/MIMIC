module fake_jpeg_2948_n_42 (n_3, n_2, n_1, n_0, n_4, n_5, n_42);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_42;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx3_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

BUFx2_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx8_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_4),
.B(n_2),
.Y(n_9)
);

BUFx2_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_2),
.B(n_3),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_4),
.B(n_3),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_14),
.A2(n_18),
.B1(n_9),
.B2(n_7),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_0),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_19),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_12),
.B(n_4),
.C(n_5),
.Y(n_16)
);

NOR2x1_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_19),
.Y(n_20)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g18 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_9),
.A2(n_0),
.B1(n_5),
.B2(n_12),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_15),
.C(n_16),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_25),
.Y(n_29)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_20),
.B(n_16),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_26),
.A2(n_22),
.B(n_23),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_28),
.C(n_21),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_21),
.B(n_18),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_31),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_23),
.C(n_24),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_33),
.B(n_17),
.Y(n_35)
);

A2O1A1O1Ixp25_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_24),
.B(n_14),
.C(n_13),
.D(n_17),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_7),
.B(n_10),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_7),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_38),
.B(n_34),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_36),
.C(n_7),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_10),
.C(n_6),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_8),
.C(n_23),
.Y(n_42)
);


endmodule