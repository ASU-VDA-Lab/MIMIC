module real_jpeg_818_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_228;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_1),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_2),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_2),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_2),
.A2(n_53),
.B1(n_68),
.B2(n_69),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_2),
.A2(n_33),
.B1(n_36),
.B2(n_53),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_53),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_5),
.A2(n_68),
.B1(n_69),
.B2(n_72),
.Y(n_67)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_5),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_72),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_5),
.A2(n_33),
.B1(n_36),
.B2(n_72),
.Y(n_272)
);

BUFx16f_ASAP7_75t_L g90 ( 
.A(n_6),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_8),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_32)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_8),
.B(n_33),
.C(n_48),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_8),
.A2(n_35),
.B1(n_51),
.B2(n_54),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_8),
.B(n_46),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_8),
.A2(n_35),
.B1(n_68),
.B2(n_69),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_8),
.B(n_26),
.C(n_28),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_8),
.B(n_69),
.C(n_89),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_8),
.B(n_24),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_8),
.B(n_66),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_8),
.B(n_140),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_10),
.A2(n_33),
.B1(n_36),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_10),
.A2(n_41),
.B1(n_51),
.B2(n_54),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_41),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_10),
.A2(n_41),
.B1(n_68),
.B2(n_69),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_254),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_231),
.B(n_252),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_208),
.B(n_228),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_125),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_109),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_18),
.B(n_109),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_76),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_19),
.B(n_77),
.C(n_101),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_60),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_44),
.B2(n_59),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_21),
.B(n_59),
.C(n_60),
.Y(n_211)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_37),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_32),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_24),
.B(n_40),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_24),
.A2(n_32),
.B(n_158),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_24),
.A2(n_97),
.B(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_25),
.B(n_98),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_31),
.Y(n_25)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_26),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_26),
.A2(n_31),
.B1(n_33),
.B2(n_36),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_27),
.A2(n_28),
.B1(n_88),
.B2(n_89),
.Y(n_93)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_28),
.B(n_167),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_32),
.B(n_158),
.Y(n_157)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_36),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_33),
.B(n_135),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_38),
.B(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_42),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_42),
.B(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_42),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_55),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_50),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_58),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_46),
.B(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_46),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_48),
.B1(n_51),
.B2(n_54),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_50),
.B(n_56),
.Y(n_218)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_63),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_55),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_58),
.Y(n_55)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_64),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_67),
.B(n_73),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_65),
.B(n_74),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_65),
.A2(n_75),
.B(n_124),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_65),
.B(n_175),
.Y(n_189)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_66),
.B(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_67),
.A2(n_75),
.B(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_68),
.A2(n_69),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_69),
.B(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_73),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_73),
.B(n_171),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_75),
.B(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_75),
.B(n_175),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_101),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_84),
.C(n_96),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

INVxp33_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_80),
.B(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_82),
.A2(n_83),
.B(n_267),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_83),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_84),
.A2(n_85),
.B1(n_96),
.B2(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI21x1_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_91),
.B(n_94),
.Y(n_85)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_86),
.A2(n_155),
.B(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_87),
.B(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_91),
.A2(n_107),
.B(n_225),
.Y(n_249)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_95),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_92),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_92),
.B(n_108),
.Y(n_155)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_95),
.B(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_100),
.B(n_157),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_102),
.B(n_105),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_104),
.B(n_174),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_106),
.B(n_154),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_107),
.B(n_141),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.C(n_116),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_110),
.A2(n_111),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_116),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_119),
.C(n_120),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_118),
.B(n_246),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_119),
.A2(n_120),
.B1(n_121),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_123),
.B(n_189),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_124),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_146),
.B(n_207),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_143),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_127),
.B(n_143),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_132),
.C(n_137),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_128),
.A2(n_129),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_132),
.A2(n_137),
.B1(n_138),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_133),
.A2(n_134),
.B1(n_136),
.B2(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_136),
.A2(n_160),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_136),
.B(n_249),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_136),
.A2(n_160),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_139),
.B(n_155),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_140),
.B(n_142),
.Y(n_154)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

AOI21x1_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_161),
.B(n_206),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_152),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_148),
.B(n_152),
.Y(n_206)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_149),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.C(n_159),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_153),
.B(n_156),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

INVxp33_ASAP7_75t_L g246 ( 
.A(n_157),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_159),
.B(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_201),
.B(n_205),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_183),
.B(n_200),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_169),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_169),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_165),
.A2(n_166),
.B1(n_168),
.B2(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_176),
.B1(n_177),
.B2(n_182),
.Y(n_169)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_170),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_178),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_179),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_180),
.C(n_182),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_190),
.B(n_199),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_187),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_187),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_195),
.B(n_198),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_196),
.B(n_197),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_203),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_229),
.B(n_230),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_227),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_227),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_211),
.B(n_213),
.C(n_223),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_222),
.B2(n_223),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_219),
.C(n_220),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_216)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_217),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_219),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_226),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_251),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_251),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_236),
.C(n_248),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_247),
.B2(n_248),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_240),
.C(n_245),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_244),
.B2(n_245),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_249),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_274),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_258),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_268),
.B2(n_269),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_271),
.B(n_273),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_270),
.B(n_271),
.Y(n_273)
);


endmodule