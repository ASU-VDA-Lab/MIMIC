module fake_jpeg_6146_n_40 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_40);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_40;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

AND2x2_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_7),
.Y(n_20)
);

OAI21xp33_ASAP7_75t_SL g21 ( 
.A1(n_3),
.A2(n_8),
.B(n_6),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_11),
.C(n_19),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_20),
.A2(n_9),
.B1(n_1),
.B2(n_2),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_29),
.C(n_30),
.Y(n_34)
);

AO21x2_ASAP7_75t_L g29 ( 
.A1(n_22),
.A2(n_21),
.B(n_23),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_0),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_32),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_24),
.B(n_5),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_36),
.B(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_34),
.Y(n_39)
);

AOI221xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_35),
.B1(n_17),
.B2(n_15),
.C(n_27),
.Y(n_40)
);


endmodule