module real_jpeg_24218_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_4),
.A2(n_40),
.B1(n_79),
.B2(n_144),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_4),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_4),
.A2(n_52),
.B1(n_55),
.B2(n_144),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_144),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_4),
.A2(n_25),
.B1(n_28),
.B2(n_144),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_5),
.A2(n_52),
.B1(n_55),
.B2(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_5),
.A2(n_63),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_63),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_5),
.A2(n_25),
.B1(n_28),
.B2(n_63),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_6),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_6),
.B(n_51),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_6),
.B(n_32),
.C(n_67),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_6),
.A2(n_52),
.B1(n_55),
.B2(n_186),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_6),
.B(n_70),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_186),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_6),
.B(n_25),
.C(n_27),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_6),
.A2(n_102),
.B(n_276),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_7),
.A2(n_40),
.B1(n_57),
.B2(n_59),
.Y(n_56)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_7),
.A2(n_52),
.B1(n_55),
.B2(n_59),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_59),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_7),
.A2(n_25),
.B1(n_28),
.B2(n_59),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_9),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_38)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_9),
.A2(n_43),
.B1(n_52),
.B2(n_55),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_43),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_9),
.A2(n_25),
.B1(n_28),
.B2(n_43),
.Y(n_226)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_11),
.A2(n_41),
.B1(n_42),
.B2(n_160),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_11),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_11),
.A2(n_52),
.B1(n_55),
.B2(n_160),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_160),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_11),
.A2(n_25),
.B1(n_28),
.B2(n_160),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_13),
.A2(n_36),
.B1(n_52),
.B2(n_55),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_13),
.A2(n_25),
.B1(n_28),
.B2(n_36),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_14),
.A2(n_47),
.B1(n_80),
.B2(n_115),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_14),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_14),
.A2(n_52),
.B1(n_55),
.B2(n_115),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_115),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_14),
.A2(n_25),
.B1(n_28),
.B2(n_115),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_15),
.A2(n_52),
.B1(n_55),
.B2(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_73),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_15),
.A2(n_25),
.B1(n_28),
.B2(n_73),
.Y(n_131)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_16),
.Y(n_103)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_16),
.Y(n_104)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_16),
.Y(n_134)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_16),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_118),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_116),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_87),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_20),
.B(n_87),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_74),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_37),
.C(n_60),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_22),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_81)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_22),
.A2(n_60),
.B1(n_85),
.B2(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_29),
.B(n_34),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_23),
.A2(n_29),
.B1(n_99),
.B2(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_23),
.A2(n_29),
.B1(n_109),
.B2(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_23),
.A2(n_29),
.B1(n_248),
.B2(n_250),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_23),
.B(n_214),
.Y(n_264)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_24),
.A2(n_35),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_24),
.A2(n_97),
.B1(n_138),
.B2(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_24),
.A2(n_172),
.B(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_24),
.A2(n_213),
.B(n_249),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_24),
.B(n_186),
.Y(n_296)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_24)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_25),
.B(n_103),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_28),
.B(n_301),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_29),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_29),
.B(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_31),
.A2(n_32),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_32),
.B(n_284),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_37),
.A2(n_75),
.B1(n_76),
.B2(n_86),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_37),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_37),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_44),
.B1(n_50),
.B2(n_56),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_38),
.A2(n_50),
.B(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_42),
.B(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_44),
.A2(n_50),
.B1(n_56),
.B2(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_44),
.A2(n_142),
.B(n_145),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_45),
.B(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_45),
.A2(n_51),
.B1(n_143),
.B2(n_159),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_45),
.A2(n_146),
.B(n_216),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_50),
.Y(n_45)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_48),
.A2(n_49),
.B1(n_52),
.B2(n_55),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_48),
.A2(n_52),
.B(n_185),
.C(n_187),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_SL g187 ( 
.A(n_49),
.B(n_55),
.C(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_50),
.B(n_114),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_50),
.A2(n_112),
.B(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_55),
.B1(n_67),
.B2(n_68),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_52),
.B(n_241),
.Y(n_240)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_57),
.Y(n_188)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_60),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_64),
.B1(n_70),
.B2(n_71),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_62),
.A2(n_65),
.B1(n_66),
.B2(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_64),
.B(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_64),
.A2(n_70),
.B1(n_180),
.B2(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_65),
.A2(n_66),
.B1(n_72),
.B2(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_65),
.A2(n_66),
.B1(n_95),
.B2(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_65),
.A2(n_179),
.B(n_181),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_L g252 ( 
.A1(n_65),
.A2(n_181),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_66),
.A2(n_140),
.B(n_163),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_66),
.A2(n_163),
.B(n_222),
.Y(n_221)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_70),
.B(n_164),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_81),
.Y(n_76)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_92),
.C(n_100),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_88),
.A2(n_92),
.B1(n_93),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_93),
.A2(n_94),
.B(n_96),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_97),
.A2(n_263),
.B(n_264),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_97),
.A2(n_264),
.B(n_282),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_100),
.B(n_148),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_106),
.B(n_110),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_110),
.B1(n_111),
.B2(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_101),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_101),
.A2(n_107),
.B1(n_108),
.B2(n_123),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_104),
.B(n_105),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_102),
.A2(n_105),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_102),
.A2(n_131),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_102),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_102),
.A2(n_192),
.B1(n_194),
.B2(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_102),
.B(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_102),
.A2(n_275),
.B(n_276),
.Y(n_274)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_103),
.Y(n_290)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_104),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_150),
.B(n_334),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_147),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_120),
.B(n_147),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.C(n_126),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_121),
.A2(n_124),
.B1(n_125),
.B2(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_121),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_126),
.A2(n_127),
.B1(n_329),
.B2(n_331),
.Y(n_328)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_139),
.C(n_141),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_128),
.A2(n_129),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_135),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_130),
.A2(n_135),
.B1(n_136),
.B2(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_130),
.Y(n_174)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_SL g244 ( 
.A(n_134),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_139),
.B(n_141),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_327),
.B(n_333),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_202),
.B(n_326),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_195),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_153),
.B(n_195),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_173),
.C(n_175),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_154),
.A2(n_155),
.B1(n_173),
.B2(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_165),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_161),
.B2(n_162),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_161),
.C(n_165),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_159),
.Y(n_177)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_171),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_166),
.B(n_171),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_168),
.A2(n_190),
.B1(n_191),
.B2(n_193),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_169),
.B(n_186),
.Y(n_301)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_173),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_175),
.B(n_323),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.C(n_182),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_176),
.B(n_178),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_182),
.B(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_189),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_183),
.A2(n_184),
.B1(n_189),
.B2(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g216 ( 
.A1(n_185),
.A2(n_186),
.B(n_188),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_190),
.A2(n_288),
.B1(n_290),
.B2(n_291),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_194),
.A2(n_289),
.B(n_298),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_201),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_197),
.B(n_198),
.C(n_201),
.Y(n_332)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

O2A1O1Ixp33_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_233),
.B(n_320),
.C(n_325),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_227),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_227),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_217),
.C(n_220),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_205),
.A2(n_206),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_215),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_211),
.B2(n_212),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_211),
.C(n_215),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_210),
.Y(n_222)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_217),
.A2(n_218),
.B1(n_220),
.B2(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_220),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.C(n_225),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_221),
.B(n_257),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_226),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_228),
.B(n_231),
.C(n_232),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_313),
.B(n_319),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_265),
.B(n_312),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_254),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_238),
.B(n_254),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_247),
.C(n_251),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_239),
.B(n_308),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_242),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B(n_245),
.Y(n_242)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_245),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_246),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_247),
.A2(n_251),
.B1(n_252),
.B2(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_247),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_250),
.Y(n_263)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_259),
.B2(n_260),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_255),
.B(n_261),
.C(n_262),
.Y(n_318)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_306),
.B(n_311),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_285),
.B(n_305),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_279),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_268),
.B(n_279),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_274),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_270),
.B(n_273),
.C(n_274),
.Y(n_310)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_275),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_283),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_280),
.A2(n_281),
.B1(n_283),
.B2(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_283),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_294),
.B(n_304),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_292),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_292),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_299),
.B(n_303),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_297),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_302),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_310),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_310),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_318),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_318),
.Y(n_319)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_322),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_332),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_332),
.Y(n_333)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_329),
.Y(n_331)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);


endmodule