module real_jpeg_14414_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_1),
.A2(n_33),
.B1(n_70),
.B2(n_72),
.Y(n_94)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g92 ( 
.A(n_3),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_4),
.A2(n_37),
.B(n_38),
.C(n_44),
.Y(n_36)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_4),
.A2(n_40),
.B1(n_44),
.B2(n_45),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_4),
.B(n_108),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_4),
.A2(n_40),
.B1(n_70),
.B2(n_72),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_4),
.A2(n_82),
.B1(n_86),
.B2(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_4),
.B(n_75),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_5),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_5),
.A2(n_41),
.B1(n_42),
.B2(n_57),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_5),
.A2(n_57),
.B1(n_70),
.B2(n_72),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_57),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_10),
.A2(n_41),
.B1(n_42),
.B2(n_60),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_10),
.A2(n_60),
.B1(n_70),
.B2(n_72),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_60),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_12),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_12),
.A2(n_70),
.B1(n_72),
.B2(n_88),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_13),
.A2(n_41),
.B1(n_42),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_13),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_13),
.A2(n_70),
.B1(n_72),
.B2(n_77),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_77),
.Y(n_137)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_15),
.A2(n_41),
.B1(n_42),
.B2(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_15),
.A2(n_64),
.B1(n_70),
.B2(n_72),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_64),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_126),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_124),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_109),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_20),
.B(n_109),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_79),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_48),
.B1(n_49),
.B2(n_78),
.Y(n_21)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_23),
.A2(n_24),
.B1(n_36),
.B2(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_24)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_25),
.B(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_25),
.A2(n_85),
.B(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_25),
.A2(n_30),
.B1(n_165),
.B2(n_167),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_26),
.A2(n_27),
.B1(n_91),
.B2(n_93),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_26),
.B(n_40),
.C(n_91),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_26),
.B(n_172),
.Y(n_171)
);

CKINVDCx6p67_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_30),
.B(n_137),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_32),
.A2(n_86),
.B(n_116),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_34),
.Y(n_83)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_36),
.Y(n_113)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B(n_41),
.Y(n_38)
);

HAxp5_ASAP7_75t_SL g134 ( 
.A(n_40),
.B(n_42),
.CON(n_134),
.SN(n_134)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_40),
.B(n_86),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_40),
.B(n_90),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_41),
.A2(n_42),
.B1(n_68),
.B2(n_69),
.Y(n_73)
);

NOR3xp33_ASAP7_75t_L g135 ( 
.A(n_41),
.B(n_69),
.C(n_70),
.Y(n_135)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_61),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_54),
.B1(n_55),
.B2(n_58),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_52),
.A2(n_56),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_65),
.B(n_74),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_63),
.A2(n_66),
.B1(n_75),
.B2(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_65),
.A2(n_67),
.B1(n_121),
.B2(n_123),
.Y(n_120)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_66),
.A2(n_75),
.B1(n_122),
.B2(n_134),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_73),
.Y(n_66)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

OA22x2_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_67)
);

O2A1O1Ixp33_ASAP7_75t_SL g132 ( 
.A1(n_68),
.A2(n_72),
.B(n_133),
.C(n_135),
.Y(n_132)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_70),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_70),
.A2(n_72),
.B1(n_91),
.B2(n_93),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_72),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_100),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_89),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B(n_84),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_82),
.A2(n_86),
.B1(n_166),
.B2(n_174),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_82),
.A2(n_168),
.B(n_184),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_94),
.B(n_95),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_97),
.Y(n_103)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_90),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_SL g93 ( 
.A(n_91),
.Y(n_93)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_98),
.A2(n_102),
.B(n_103),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_98),
.A2(n_141),
.B1(n_143),
.B2(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_98),
.A2(n_143),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_98),
.A2(n_143),
.B1(n_151),
.B2(n_161),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_104),
.C(n_106),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_104),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_143),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_105),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.C(n_114),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_110),
.B(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_112),
.B(n_114),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.C(n_120),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_118),
.B1(n_119),
.B2(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_120),
.B(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_197),
.B(n_201),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_152),
.B(n_196),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_147),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_129),
.B(n_147),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_144),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_138),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_131),
.B(n_138),
.C(n_144),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_136),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_132),
.B(n_136),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_140),
.B(n_142),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.C(n_150),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_150),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_191),
.B(n_195),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_180),
.B(n_190),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_169),
.B(n_179),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_164),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_164),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_159),
.B1(n_162),
.B2(n_163),
.Y(n_156)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_157),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_159),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_162),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_175),
.B(n_178),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_177),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_182),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_186),
.C(n_189),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_188),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_194),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_200),
.Y(n_201)
);


endmodule