module fake_jpeg_15083_n_317 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx8_ASAP7_75t_SL g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_34),
.Y(n_40)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_30),
.A2(n_27),
.B1(n_23),
.B2(n_25),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_41),
.A2(n_44),
.B1(n_16),
.B2(n_28),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_52),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_27),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_18),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_30),
.A2(n_23),
.B1(n_15),
.B2(n_25),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_49),
.B(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_19),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_19),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_51),
.B(n_35),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_34),
.B(n_28),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_33),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_20),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_33),
.A2(n_23),
.B1(n_18),
.B2(n_21),
.Y(n_57)
);

OAI32xp33_ASAP7_75t_L g77 ( 
.A1(n_57),
.A2(n_29),
.A3(n_33),
.B1(n_28),
.B2(n_16),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_56),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_59),
.Y(n_83)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_23),
.B1(n_32),
.B2(n_36),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_61),
.A2(n_65),
.B1(n_68),
.B2(n_79),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_64),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_67),
.Y(n_81)
);

OR2x2_ASAP7_75t_SL g64 ( 
.A(n_40),
.B(n_23),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_32),
.B1(n_23),
.B2(n_36),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_38),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_32),
.B1(n_38),
.B2(n_36),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_73),
.B1(n_16),
.B2(n_67),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_38),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_74),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_47),
.A2(n_16),
.B1(n_28),
.B2(n_14),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_37),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_37),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_76),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_37),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_48),
.B1(n_53),
.B2(n_57),
.Y(n_91)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_41),
.A2(n_45),
.B1(n_48),
.B2(n_53),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_84),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_62),
.A2(n_79),
.B1(n_77),
.B2(n_59),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_91),
.B1(n_98),
.B2(n_100),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_95),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_54),
.C(n_33),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_101),
.C(n_29),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_102),
.B1(n_57),
.B2(n_29),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_50),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_75),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_70),
.A2(n_48),
.B1(n_53),
.B2(n_46),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_74),
.A2(n_46),
.B1(n_39),
.B2(n_57),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_55),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_63),
.A2(n_46),
.B1(n_39),
.B2(n_57),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_77),
.A2(n_60),
.B1(n_66),
.B2(n_65),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_104),
.A2(n_76),
.B1(n_64),
.B2(n_68),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_88),
.A2(n_60),
.B1(n_80),
.B2(n_58),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_124),
.B1(n_88),
.B2(n_85),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_110),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_96),
.B(n_75),
.Y(n_110)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_80),
.B(n_73),
.C(n_39),
.Y(n_113)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_72),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_116),
.Y(n_149)
);

OA21x2_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_76),
.B(n_66),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_118),
.B1(n_94),
.B2(n_90),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_72),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_103),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_97),
.A2(n_64),
.B(n_65),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_126),
.B(n_127),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_91),
.A2(n_80),
.B1(n_57),
.B2(n_58),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_120),
.A2(n_100),
.B1(n_85),
.B2(n_93),
.Y(n_145)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_56),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_0),
.Y(n_126)
);

AND2x2_ASAP7_75t_SL g127 ( 
.A(n_99),
.B(n_58),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_56),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_129),
.B(n_86),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_131),
.A2(n_145),
.B1(n_151),
.B2(n_141),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_141),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_81),
.C(n_108),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_153),
.C(n_127),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_138),
.A2(n_110),
.B1(n_113),
.B2(n_107),
.Y(n_161)
);

NOR3xp33_ASAP7_75t_SL g141 ( 
.A(n_115),
.B(n_104),
.C(n_89),
.Y(n_141)
);

OAI32xp33_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_81),
.A3(n_118),
.B1(n_116),
.B2(n_114),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_154),
.Y(n_162)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_148),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_124),
.A2(n_93),
.B1(n_90),
.B2(n_92),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_107),
.B1(n_120),
.B2(n_115),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_121),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_122),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_152),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_101),
.B1(n_20),
.B2(n_14),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

OAI32xp33_ASAP7_75t_L g154 ( 
.A1(n_109),
.A2(n_113),
.A3(n_115),
.B1(n_111),
.B2(n_126),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_152),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_161),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_119),
.B(n_105),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_160),
.A2(n_165),
.B(n_136),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_143),
.A2(n_126),
.B(n_105),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_132),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_166),
.B(n_170),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_167),
.A2(n_180),
.B1(n_139),
.B2(n_26),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_175),
.C(n_178),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_132),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_149),
.B(n_127),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_171),
.B(n_174),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_172),
.A2(n_26),
.B1(n_21),
.B2(n_17),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_112),
.Y(n_173)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_117),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_137),
.B(n_127),
.C(n_126),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_130),
.A2(n_117),
.B1(n_56),
.B2(n_20),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_176),
.A2(n_177),
.B1(n_133),
.B2(n_146),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_136),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_140),
.C(n_138),
.Y(n_178)
);

AOI322xp5_ASAP7_75t_L g179 ( 
.A1(n_142),
.A2(n_24),
.A3(n_26),
.B1(n_21),
.B2(n_17),
.C1(n_18),
.C2(n_13),
.Y(n_179)
);

NAND3xp33_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_18),
.C(n_13),
.Y(n_191)
);

AOI22x1_ASAP7_75t_L g180 ( 
.A1(n_154),
.A2(n_26),
.B1(n_24),
.B2(n_21),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_26),
.Y(n_181)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_181),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_145),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_167),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_133),
.Y(n_183)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_185),
.B(n_158),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_206),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_168),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_187),
.B(n_196),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_192),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_163),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_155),
.Y(n_195)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_195),
.Y(n_211)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_156),
.Y(n_198)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_198),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_178),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_201),
.C(n_171),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_139),
.Y(n_201)
);

NAND2x1_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_159),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_202),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_203),
.A2(n_207),
.B1(n_180),
.B2(n_177),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_162),
.A2(n_0),
.B(n_1),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_204),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_164),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_205),
.B(n_170),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_24),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_165),
.A2(n_0),
.B(n_1),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_162),
.B(n_161),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_160),
.Y(n_217)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_209),
.Y(n_214)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_210),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_198),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_213),
.Y(n_251)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_219),
.Y(n_232)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_218),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_206),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_197),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_220),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_157),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_223),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_157),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_224),
.A2(n_176),
.B1(n_203),
.B2(n_207),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_164),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_226),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_229),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_184),
.B(n_158),
.C(n_166),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_231),
.B(n_184),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_226),
.A2(n_200),
.B1(n_202),
.B2(n_186),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_234),
.A2(n_250),
.B1(n_188),
.B2(n_216),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_202),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_237),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_244),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_201),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_248),
.C(n_249),
.Y(n_258)
);

BUFx24_ASAP7_75t_SL g244 ( 
.A(n_228),
.Y(n_244)
);

HAxp5_ASAP7_75t_SL g245 ( 
.A(n_225),
.B(n_185),
.CON(n_245),
.SN(n_245)
);

XNOR2x1_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_227),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_246),
.A2(n_214),
.B1(n_230),
.B2(n_222),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_217),
.A2(n_208),
.B(n_197),
.Y(n_247)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_247),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_209),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_227),
.A2(n_188),
.B1(n_183),
.B2(n_190),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_252),
.A2(n_4),
.B(n_5),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_253),
.A2(n_236),
.B1(n_239),
.B2(n_250),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_243),
.B(n_210),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_260),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_224),
.Y(n_256)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_256),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_257),
.A2(n_261),
.B1(n_237),
.B2(n_235),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_233),
.C(n_249),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_265),
.C(n_266),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_219),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_242),
.A2(n_216),
.B1(n_4),
.B2(n_5),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_234),
.B(n_3),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_237),
.Y(n_273)
);

BUFx4f_ASAP7_75t_SL g263 ( 
.A(n_245),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_268),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_21),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_18),
.C(n_17),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_21),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_269),
.A2(n_282),
.B1(n_262),
.B2(n_263),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_273),
.B(n_274),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_232),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_275),
.C(n_279),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_252),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_279),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_254),
.B(n_18),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_281),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_3),
.Y(n_279)
);

A2O1A1Ixp33_ASAP7_75t_L g280 ( 
.A1(n_267),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_280),
.A2(n_8),
.B(n_9),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_264),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_258),
.Y(n_284)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_284),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_266),
.Y(n_286)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_286),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_272),
.B(n_263),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_288),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_283),
.C(n_290),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_273),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_294),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_18),
.C(n_21),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_292),
.B(n_293),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_270),
.B(n_17),
.C(n_21),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_277),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_303),
.C(n_17),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_283),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_301),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_280),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_296),
.A2(n_8),
.B(n_10),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_305),
.A2(n_306),
.B(n_307),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_17),
.C(n_11),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_298),
.C(n_295),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_308),
.A2(n_10),
.B(n_11),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_17),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_309),
.A2(n_302),
.B(n_11),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_311),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_312),
.A2(n_10),
.B1(n_12),
.B2(n_304),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_310),
.C(n_17),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_313),
.C(n_12),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_12),
.Y(n_317)
);


endmodule