module fake_aes_7558_n_22 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_22);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_22;
wire n_20;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
wire n_7;
INVx1_ASAP7_75t_L g7 ( .A(n_6), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_4), .Y(n_8) );
AND2x4_ASAP7_75t_L g9 ( .A(n_3), .B(n_0), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_0), .Y(n_10) );
AND2x2_ASAP7_75t_SL g11 ( .A(n_4), .B(n_1), .Y(n_11) );
BUFx6f_ASAP7_75t_L g12 ( .A(n_7), .Y(n_12) );
INVx3_ASAP7_75t_L g13 ( .A(n_9), .Y(n_13) );
AOI22xp33_ASAP7_75t_L g14 ( .A1(n_9), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_14) );
BUFx2_ASAP7_75t_L g15 ( .A(n_13), .Y(n_15) );
AOI211xp5_ASAP7_75t_L g16 ( .A1(n_13), .A2(n_8), .B(n_10), .C(n_9), .Y(n_16) );
INVxp67_ASAP7_75t_L g17 ( .A(n_15), .Y(n_17) );
NOR3xp33_ASAP7_75t_SL g18 ( .A(n_16), .B(n_7), .C(n_11), .Y(n_18) );
AOI211xp5_ASAP7_75t_L g19 ( .A1(n_17), .A2(n_12), .B(n_11), .C(n_14), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
OAI21xp5_ASAP7_75t_L g21 ( .A1(n_19), .A2(n_18), .B(n_14), .Y(n_21) );
AOI222xp33_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_2), .B1(n_5), .B2(n_12), .C1(n_20), .C2(n_11), .Y(n_22) );
endmodule