module fake_ibex_1269_n_184 (n_7, n_20, n_40, n_17, n_25, n_36, n_18, n_3, n_22, n_28, n_32, n_39, n_4, n_33, n_5, n_11, n_30, n_6, n_29, n_13, n_2, n_8, n_26, n_35, n_14, n_0, n_9, n_34, n_12, n_38, n_15, n_37, n_24, n_31, n_10, n_23, n_21, n_27, n_19, n_16, n_1, n_184);

input n_7;
input n_20;
input n_40;
input n_17;
input n_25;
input n_36;
input n_18;
input n_3;
input n_22;
input n_28;
input n_32;
input n_39;
input n_4;
input n_33;
input n_5;
input n_11;
input n_30;
input n_6;
input n_29;
input n_13;
input n_2;
input n_8;
input n_26;
input n_35;
input n_14;
input n_0;
input n_9;
input n_34;
input n_12;
input n_38;
input n_15;
input n_37;
input n_24;
input n_31;
input n_10;
input n_23;
input n_21;
input n_27;
input n_19;
input n_16;
input n_1;

output n_184;

wire n_151;
wire n_147;
wire n_85;
wire n_167;
wire n_128;
wire n_84;
wire n_64;
wire n_73;
wire n_152;
wire n_171;
wire n_145;
wire n_65;
wire n_103;
wire n_95;
wire n_139;
wire n_55;
wire n_130;
wire n_63;
wire n_98;
wire n_129;
wire n_161;
wire n_143;
wire n_106;
wire n_177;
wire n_148;
wire n_76;
wire n_118;
wire n_183;
wire n_67;
wire n_164;
wire n_124;
wire n_110;
wire n_47;
wire n_169;
wire n_108;
wire n_82;
wire n_165;
wire n_78;
wire n_60;
wire n_86;
wire n_70;
wire n_87;
wire n_69;
wire n_75;
wire n_109;
wire n_127;
wire n_121;
wire n_175;
wire n_137;
wire n_48;
wire n_57;
wire n_59;
wire n_125;
wire n_178;
wire n_62;
wire n_71;
wire n_153;
wire n_173;
wire n_120;
wire n_93;
wire n_168;
wire n_155;
wire n_162;
wire n_180;
wire n_122;
wire n_116;
wire n_61;
wire n_94;
wire n_134;
wire n_42;
wire n_77;
wire n_112;
wire n_150;
wire n_88;
wire n_133;
wire n_44;
wire n_142;
wire n_51;
wire n_46;
wire n_80;
wire n_172;
wire n_49;
wire n_66;
wire n_74;
wire n_90;
wire n_176;
wire n_58;
wire n_43;
wire n_140;
wire n_136;
wire n_119;
wire n_100;
wire n_179;
wire n_72;
wire n_166;
wire n_163;
wire n_114;
wire n_97;
wire n_102;
wire n_181;
wire n_131;
wire n_123;
wire n_52;
wire n_99;
wire n_135;
wire n_105;
wire n_156;
wire n_126;
wire n_154;
wire n_182;
wire n_111;
wire n_104;
wire n_41;
wire n_141;
wire n_89;
wire n_83;
wire n_53;
wire n_107;
wire n_115;
wire n_149;
wire n_54;
wire n_50;
wire n_92;
wire n_144;
wire n_170;
wire n_101;
wire n_113;
wire n_138;
wire n_96;
wire n_68;
wire n_117;
wire n_79;
wire n_81;
wire n_159;
wire n_158;
wire n_132;
wire n_174;
wire n_157;
wire n_160;
wire n_56;
wire n_146;
wire n_91;
wire n_45;

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

INVxp33_ASAP7_75t_SL g44 ( 
.A(n_4),
.Y(n_44)
);

INVxp33_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_27),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_20),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

NOR2xp67_ASAP7_75t_L g50 ( 
.A(n_6),
.B(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVxp67_ASAP7_75t_SL g52 ( 
.A(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_30),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_0),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_8),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_2),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_5),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_35),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_37),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_19),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_3),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_34),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_R g70 ( 
.A(n_7),
.B(n_38),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_6),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_24),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_23),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_13),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_10),
.Y(n_76)
);

INVxp67_ASAP7_75t_SL g77 ( 
.A(n_9),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_11),
.Y(n_79)
);

AND2x4_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_1),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_57),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_42),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_41),
.B(n_1),
.Y(n_83)
);

CKINVDCx8_ASAP7_75t_R g84 ( 
.A(n_58),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_69),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_44),
.A2(n_4),
.B1(n_9),
.B2(n_12),
.Y(n_88)
);

AND2x6_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_16),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_17),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_25),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_79),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_78),
.Y(n_93)
);

NAND3xp33_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_39),
.C(n_71),
.Y(n_94)
);

NOR3xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_61),
.C(n_50),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_47),
.B(n_73),
.Y(n_97)
);

OR2x6_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_67),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_43),
.B(n_66),
.Y(n_99)
);

NAND2xp33_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_72),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_70),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_43),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_67),
.B(n_49),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

OR2x6_ASAP7_75t_L g108 ( 
.A(n_54),
.B(n_76),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_54),
.B(n_66),
.Y(n_109)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_64),
.B(n_41),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_85),
.B(n_87),
.C(n_83),
.Y(n_115)
);

NAND3xp33_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_105),
.C(n_81),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_113),
.A2(n_90),
.B(n_93),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_113),
.A2(n_90),
.B(n_93),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_97),
.B(n_100),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_92),
.A2(n_97),
.B(n_86),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_82),
.B1(n_98),
.B2(n_80),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_96),
.A2(n_91),
.B(n_101),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_84),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_89),
.A2(n_94),
.B(n_80),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_89),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_98),
.A2(n_99),
.B1(n_88),
.B2(n_110),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_98),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_112),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_99),
.A2(n_110),
.B1(n_108),
.B2(n_111),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_111),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_111),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_89),
.A2(n_109),
.B(n_106),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_109),
.A2(n_87),
.B(n_92),
.C(n_93),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_108),
.A2(n_113),
.B(n_90),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_104),
.A2(n_113),
.B(n_90),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_90),
.B(n_93),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_82),
.Y(n_140)
);

NAND2xp33_ASAP7_75t_L g141 ( 
.A(n_89),
.B(n_91),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_113),
.A2(n_90),
.B(n_93),
.Y(n_143)
);

OR2x6_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_128),
.Y(n_144)
);

INVx3_ASAP7_75t_SL g145 ( 
.A(n_134),
.Y(n_145)
);

AND2x4_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_140),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

AND2x4_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_137),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_121),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_141),
.A2(n_143),
.B(n_139),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_129),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_117),
.A2(n_118),
.B(n_120),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_119),
.B(n_135),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_115),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_126),
.A2(n_136),
.B(n_133),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_136),
.Y(n_157)
);

OR2x6_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_124),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_148),
.Y(n_162)
);

AND2x4_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_158),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_158),
.Y(n_164)
);

AO21x2_ASAP7_75t_L g165 ( 
.A1(n_154),
.A2(n_151),
.B(n_156),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_146),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_146),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_150),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_163),
.A2(n_144),
.B1(n_145),
.B2(n_158),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_147),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_144),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_144),
.Y(n_172)
);

NAND3xp33_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_153),
.C(n_155),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_153),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_163),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_175),
.Y(n_176)
);

NAND3xp33_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_173),
.C(n_169),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_177),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_178),
.Y(n_179)
);

XNOR2x1_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_172),
.Y(n_180)
);

AND4x1_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_170),
.C(n_171),
.D(n_167),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_164),
.B1(n_165),
.B2(n_163),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_174),
.B(n_167),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_183),
.A2(n_164),
.B1(n_163),
.B2(n_165),
.Y(n_184)
);


endmodule