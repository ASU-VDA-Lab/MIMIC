module fake_jpeg_1779_n_298 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_1),
.B(n_5),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_40),
.B(n_30),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_15),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_28),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_60),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_32),
.B1(n_16),
.B2(n_18),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_57),
.A2(n_78),
.B1(n_90),
.B2(n_100),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_35),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_58),
.B(n_84),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_29),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_25),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_25),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_61),
.B(n_65),
.Y(n_107)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_62),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_45),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_69),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_24),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_43),
.A2(n_16),
.B1(n_19),
.B2(n_36),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_70),
.A2(n_96),
.B1(n_92),
.B2(n_55),
.Y(n_113)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_73),
.Y(n_132)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_42),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_75),
.Y(n_103)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_42),
.A2(n_32),
.B1(n_18),
.B2(n_22),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_38),
.B(n_34),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_79),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_46),
.B(n_34),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_80),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_44),
.B(n_33),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_83),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_33),
.Y(n_84)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_46),
.B(n_22),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_88),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_24),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_43),
.B(n_24),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_21),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_36),
.C(n_23),
.Y(n_112)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

BUFx12_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

AO22x1_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_96),
.B1(n_98),
.B2(n_101),
.Y(n_108)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_47),
.A2(n_20),
.B1(n_19),
.B2(n_23),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_27),
.B1(n_1),
.B2(n_2),
.Y(n_116)
);

INVxp67_ASAP7_75t_SL g100 ( 
.A(n_50),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_SL g105 ( 
.A1(n_75),
.A2(n_27),
.B(n_20),
.C(n_2),
.Y(n_105)
);

OA21x2_ASAP7_75t_L g166 ( 
.A1(n_105),
.A2(n_121),
.B(n_126),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_36),
.B1(n_23),
.B2(n_27),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_106),
.A2(n_116),
.B1(n_123),
.B2(n_124),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_62),
.C(n_72),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_128),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_58),
.A2(n_27),
.B1(n_1),
.B2(n_2),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_69),
.A2(n_0),
.B(n_3),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_122),
.A2(n_62),
.B(n_72),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_89),
.A2(n_14),
.B1(n_9),
.B2(n_6),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_89),
.A2(n_10),
.B1(n_13),
.B2(n_7),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_82),
.A2(n_55),
.B1(n_69),
.B2(n_77),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_82),
.A2(n_11),
.B1(n_13),
.B2(n_7),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_67),
.A2(n_0),
.B1(n_3),
.B2(n_7),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_0),
.Y(n_154)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_74),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_136),
.Y(n_170)
);

AO21x1_ASAP7_75t_L g179 ( 
.A1(n_135),
.A2(n_141),
.B(n_165),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_74),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_129),
.B(n_81),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_137),
.B(n_138),
.Y(n_167)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_110),
.A2(n_81),
.B(n_67),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_142),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_98),
.C(n_64),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_149),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_145),
.Y(n_195)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_146),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_147),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_112),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_152),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_102),
.B(n_64),
.C(n_71),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_107),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_153),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_86),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_156),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_102),
.B(n_71),
.C(n_94),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_158),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_125),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_111),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_157),
.A2(n_162),
.B1(n_125),
.B2(n_103),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_95),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_130),
.B(n_63),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_159),
.B(n_103),
.Y(n_175)
);

MAJx2_ASAP7_75t_L g160 ( 
.A(n_102),
.B(n_130),
.C(n_120),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_164),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_161),
.Y(n_168)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_163),
.Y(n_177)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_108),
.Y(n_164)
);

AND2x4_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_95),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_166),
.A2(n_144),
.B1(n_148),
.B2(n_165),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_172),
.A2(n_180),
.B1(n_189),
.B2(n_196),
.Y(n_204)
);

OAI22x1_ASAP7_75t_L g173 ( 
.A1(n_165),
.A2(n_105),
.B1(n_120),
.B2(n_104),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_173),
.A2(n_188),
.B1(n_192),
.B2(n_186),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_175),
.B(n_181),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_166),
.A2(n_113),
.B1(n_121),
.B2(n_116),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_143),
.B(n_104),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_122),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_190),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_144),
.A2(n_150),
.B1(n_166),
.B2(n_135),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_188),
.A2(n_63),
.B1(n_101),
.B2(n_73),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_144),
.A2(n_105),
.B1(n_128),
.B2(n_124),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_138),
.B(n_126),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_165),
.A2(n_132),
.B1(n_93),
.B2(n_97),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_149),
.A2(n_108),
.B1(n_123),
.B2(n_132),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_118),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_197),
.B(n_118),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_145),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_147),
.Y(n_215)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_199),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_195),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_208),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_193),
.B(n_155),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_207),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_179),
.A2(n_141),
.B(n_156),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_206),
.A2(n_209),
.B(n_210),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_193),
.B(n_133),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_162),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_180),
.A2(n_157),
.B1(n_161),
.B2(n_163),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_212),
.A2(n_198),
.B1(n_177),
.B2(n_168),
.Y(n_228)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_215),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_175),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_214),
.Y(n_238)
);

NOR2xp67_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_185),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_219),
.A2(n_221),
.B1(n_206),
.B2(n_196),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_184),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_220),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_189),
.A2(n_77),
.B1(n_68),
.B2(n_85),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_181),
.B(n_94),
.C(n_54),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_190),
.C(n_183),
.Y(n_232)
);

INVxp33_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_228),
.A2(n_236),
.B1(n_221),
.B2(n_209),
.Y(n_244)
);

A2O1A1O1Ixp25_ASAP7_75t_L g229 ( 
.A1(n_217),
.A2(n_176),
.B(n_178),
.C(n_172),
.D(n_167),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_232),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_217),
.B(n_176),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_235),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_167),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_240),
.C(n_241),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_211),
.B(n_178),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_204),
.A2(n_173),
.B1(n_185),
.B2(n_177),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_208),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_174),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_174),
.Y(n_241)
);

INVxp33_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_223),
.A2(n_214),
.B(n_240),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_245),
.A2(n_255),
.B(n_223),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_242),
.B(n_222),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_250),
.Y(n_265)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_247),
.Y(n_257)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_226),
.Y(n_248)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_236),
.A2(n_218),
.B1(n_219),
.B2(n_202),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_233),
.C(n_241),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_253),
.C(n_254),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_214),
.C(n_209),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_200),
.C(n_213),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_226),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_225),
.C(n_224),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_253),
.C(n_252),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_260),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_229),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_252),
.B(n_238),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_267),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_225),
.C(n_227),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_254),
.C(n_245),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_234),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_270),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_265),
.A2(n_257),
.B(n_266),
.Y(n_271)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_271),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_264),
.A2(n_249),
.B1(n_218),
.B2(n_234),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_272),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_249),
.C(n_239),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_274),
.C(n_275),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_231),
.C(n_202),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_231),
.C(n_203),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_263),
.C(n_267),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_281),
.C(n_194),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_269),
.A2(n_264),
.B(n_262),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_169),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_228),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_283),
.A2(n_199),
.B1(n_168),
.B2(n_194),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_287),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_286),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_280),
.A2(n_195),
.B1(n_169),
.B2(n_97),
.Y(n_286)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_281),
.Y(n_288)
);

OAI221xp5_ASAP7_75t_L g291 ( 
.A1(n_288),
.A2(n_279),
.B1(n_282),
.B2(n_277),
.C(n_278),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_291),
.B(n_277),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_292),
.A2(n_293),
.B(n_289),
.Y(n_294)
);

AO21x1_ASAP7_75t_L g293 ( 
.A1(n_290),
.A2(n_287),
.B(n_288),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_54),
.Y(n_295)
);

AOI321xp33_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_93),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C(n_8),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_12),
.C(n_68),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_12),
.Y(n_298)
);


endmodule