module real_aes_7710_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_725;
wire n_504;
wire n_119;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g474 ( .A1(n_0), .A2(n_164), .B(n_475), .C(n_478), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_1), .B(n_469), .Y(n_479) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_2), .B(n_109), .C(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g124 ( .A(n_2), .Y(n_124) );
INVx1_ASAP7_75t_L g162 ( .A(n_3), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_4), .B(n_165), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_5), .A2(n_464), .B(n_537), .Y(n_536) );
AO21x2_ASAP7_75t_L g544 ( .A1(n_6), .A2(n_187), .B(n_545), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_7), .A2(n_40), .B1(n_152), .B2(n_210), .Y(n_250) );
AOI222xp33_ASAP7_75t_L g439 ( .A1(n_8), .A2(n_20), .B1(n_440), .B2(n_725), .C1(n_726), .C2(n_729), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_8), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_9), .B(n_187), .Y(n_195) );
AND2x6_ASAP7_75t_L g167 ( .A(n_10), .B(n_168), .Y(n_167) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_11), .A2(n_167), .B(n_455), .C(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g106 ( .A(n_12), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_12), .B(n_41), .Y(n_125) );
INVx1_ASAP7_75t_L g146 ( .A(n_13), .Y(n_146) );
INVx1_ASAP7_75t_L g143 ( .A(n_14), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_15), .B(n_148), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_16), .B(n_165), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_17), .B(n_139), .Y(n_197) );
AO32x2_ASAP7_75t_L g248 ( .A1(n_18), .A2(n_138), .A3(n_181), .B1(n_187), .B2(n_249), .Y(n_248) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_19), .A2(n_30), .B1(n_128), .B2(n_129), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_19), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_21), .B(n_152), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_22), .B(n_139), .Y(n_169) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_23), .A2(n_55), .B1(n_152), .B2(n_210), .Y(n_251) );
AOI22xp33_ASAP7_75t_SL g212 ( .A1(n_24), .A2(n_80), .B1(n_148), .B2(n_152), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_25), .B(n_152), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_L g485 ( .A1(n_26), .A2(n_181), .B(n_455), .C(n_486), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g547 ( .A1(n_27), .A2(n_181), .B(n_455), .C(n_548), .Y(n_547) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_28), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_29), .B(n_183), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_30), .Y(n_129) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_30), .A2(n_129), .B1(n_130), .B2(n_131), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_31), .A2(n_464), .B(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_32), .B(n_183), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_33), .B(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g150 ( .A(n_34), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_35), .A2(n_461), .B(n_504), .C(n_505), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_36), .B(n_152), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_37), .B(n_183), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g100 ( .A1(n_38), .A2(n_101), .B1(n_113), .B2(n_733), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_39), .B(n_232), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_41), .B(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_42), .B(n_484), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_43), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_44), .B(n_165), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_45), .B(n_464), .Y(n_546) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_46), .A2(n_461), .B(n_504), .C(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_47), .B(n_152), .Y(n_190) );
INVx1_ASAP7_75t_L g476 ( .A(n_48), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_49), .A2(n_89), .B1(n_210), .B2(n_211), .Y(n_209) );
INVx1_ASAP7_75t_L g529 ( .A(n_50), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_51), .B(n_152), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_52), .B(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_53), .B(n_464), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_54), .B(n_160), .Y(n_194) );
AOI22xp33_ASAP7_75t_SL g201 ( .A1(n_56), .A2(n_60), .B1(n_148), .B2(n_152), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_57), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_58), .B(n_152), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_59), .B(n_152), .Y(n_229) );
INVx1_ASAP7_75t_L g168 ( .A(n_61), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_62), .B(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_63), .B(n_469), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g539 ( .A1(n_64), .A2(n_154), .B(n_160), .C(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_65), .B(n_152), .Y(n_163) );
INVx1_ASAP7_75t_L g142 ( .A(n_66), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_67), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_68), .B(n_165), .Y(n_507) );
AO32x2_ASAP7_75t_L g207 ( .A1(n_69), .A2(n_181), .A3(n_187), .B1(n_208), .B2(n_213), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_70), .B(n_166), .Y(n_520) );
INVx1_ASAP7_75t_L g177 ( .A(n_71), .Y(n_177) );
INVx1_ASAP7_75t_L g220 ( .A(n_72), .Y(n_220) );
CKINVDCx16_ASAP7_75t_R g472 ( .A(n_73), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_74), .B(n_488), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_L g454 ( .A1(n_75), .A2(n_455), .B(n_457), .C(n_461), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_76), .B(n_148), .Y(n_221) );
CKINVDCx16_ASAP7_75t_R g538 ( .A(n_77), .Y(n_538) );
INVx1_ASAP7_75t_L g112 ( .A(n_78), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_79), .B(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_81), .B(n_210), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_82), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_83), .B(n_148), .Y(n_224) );
INVx2_ASAP7_75t_L g140 ( .A(n_84), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_85), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_86), .B(n_180), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_87), .B(n_148), .Y(n_191) );
INVx2_ASAP7_75t_L g109 ( .A(n_88), .Y(n_109) );
OR2x2_ASAP7_75t_L g121 ( .A(n_88), .B(n_122), .Y(n_121) );
OR2x2_ASAP7_75t_L g443 ( .A(n_88), .B(n_123), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_90), .A2(n_99), .B1(n_148), .B2(n_149), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_91), .B(n_464), .Y(n_502) );
INVx1_ASAP7_75t_L g506 ( .A(n_92), .Y(n_506) );
INVxp67_ASAP7_75t_L g541 ( .A(n_93), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_94), .B(n_148), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_95), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g458 ( .A(n_96), .Y(n_458) );
INVx1_ASAP7_75t_L g516 ( .A(n_97), .Y(n_516) );
AND2x2_ASAP7_75t_L g531 ( .A(n_98), .B(n_183), .Y(n_531) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_SL g733 ( .A(n_103), .Y(n_733) );
AND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_107), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OR2x2_ASAP7_75t_L g446 ( .A(n_109), .B(n_123), .Y(n_446) );
NOR2x2_ASAP7_75t_L g728 ( .A(n_109), .B(n_122), .Y(n_728) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OA21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_119), .B(n_438), .Y(n_113) );
BUFx2_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g732 ( .A(n_118), .Y(n_732) );
OAI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_126), .B(n_435), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g437 ( .A(n_121), .Y(n_437) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
AOI22xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_130), .B1(n_131), .B2(n_434), .Y(n_126) );
INVx1_ASAP7_75t_L g434 ( .A(n_127), .Y(n_434) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OR5x1_ASAP7_75t_L g131 ( .A(n_132), .B(n_325), .C(n_383), .D(n_419), .E(n_426), .Y(n_131) );
NAND3xp33_ASAP7_75t_SL g132 ( .A(n_133), .B(n_271), .C(n_295), .Y(n_132) );
AOI221xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_203), .B1(n_237), .B2(n_242), .C(n_252), .Y(n_133) );
OAI21xp5_ASAP7_75t_SL g405 ( .A1(n_134), .A2(n_406), .B(n_408), .Y(n_405) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_184), .Y(n_134) );
NAND2x1p5_ASAP7_75t_L g395 ( .A(n_135), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_170), .Y(n_135) );
INVx2_ASAP7_75t_L g241 ( .A(n_136), .Y(n_241) );
AND2x2_ASAP7_75t_L g254 ( .A(n_136), .B(n_186), .Y(n_254) );
AND2x2_ASAP7_75t_L g308 ( .A(n_136), .B(n_185), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_136), .B(n_171), .Y(n_323) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_144), .B(n_169), .Y(n_136) );
OA21x2_ASAP7_75t_L g171 ( .A1(n_137), .A2(n_172), .B(n_182), .Y(n_171) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_138), .B(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_139), .Y(n_187) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x2_ASAP7_75t_SL g183 ( .A(n_140), .B(n_141), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
OAI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_158), .B(n_167), .Y(n_144) );
O2A1O1Ixp33_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_151), .C(n_154), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_147), .A2(n_520), .B(n_521), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_147), .A2(n_549), .B(n_550), .Y(n_548) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g153 ( .A(n_150), .Y(n_153) );
INVx1_ASAP7_75t_L g161 ( .A(n_150), .Y(n_161) );
INVx3_ASAP7_75t_L g219 ( .A(n_152), .Y(n_219) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_152), .Y(n_460) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g210 ( .A(n_153), .Y(n_210) );
BUFx3_ASAP7_75t_L g211 ( .A(n_153), .Y(n_211) );
AND2x6_ASAP7_75t_L g455 ( .A(n_153), .B(n_456), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_L g457 ( .A1(n_154), .A2(n_458), .B(n_459), .C(n_460), .Y(n_457) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_155), .A2(n_223), .B(n_224), .Y(n_222) );
INVx4_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g488 ( .A(n_156), .Y(n_488) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx3_ASAP7_75t_L g166 ( .A(n_157), .Y(n_166) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_157), .Y(n_180) );
INVx1_ASAP7_75t_L g232 ( .A(n_157), .Y(n_232) );
INVx1_ASAP7_75t_L g456 ( .A(n_157), .Y(n_456) );
AND2x2_ASAP7_75t_L g465 ( .A(n_157), .B(n_161), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_162), .B(n_163), .C(n_164), .Y(n_158) );
O2A1O1Ixp5_ASAP7_75t_L g176 ( .A1(n_159), .A2(n_177), .B(n_178), .C(n_179), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_159), .A2(n_487), .B(n_489), .Y(n_486) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_164), .A2(n_193), .B(n_194), .Y(n_192) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_164), .A2(n_180), .B1(n_200), .B2(n_201), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_164), .A2(n_180), .B1(n_250), .B2(n_251), .Y(n_249) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_165), .A2(n_174), .B(n_175), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_165), .A2(n_190), .B(n_191), .Y(n_189) );
O2A1O1Ixp5_ASAP7_75t_SL g218 ( .A1(n_165), .A2(n_219), .B(n_220), .C(n_221), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_165), .B(n_541), .Y(n_540) );
INVx5_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
OAI22xp5_ASAP7_75t_SL g208 ( .A1(n_166), .A2(n_180), .B1(n_209), .B2(n_212), .Y(n_208) );
BUFx3_ASAP7_75t_L g181 ( .A(n_167), .Y(n_181) );
OAI21xp5_ASAP7_75t_L g188 ( .A1(n_167), .A2(n_189), .B(n_192), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g217 ( .A1(n_167), .A2(n_218), .B(n_222), .Y(n_217) );
OAI21xp5_ASAP7_75t_L g227 ( .A1(n_167), .A2(n_228), .B(n_233), .Y(n_227) );
INVx4_ASAP7_75t_SL g462 ( .A(n_167), .Y(n_462) );
AND2x4_ASAP7_75t_L g464 ( .A(n_167), .B(n_465), .Y(n_464) );
NAND2x1p5_ASAP7_75t_L g517 ( .A(n_167), .B(n_465), .Y(n_517) );
AND2x2_ASAP7_75t_L g341 ( .A(n_170), .B(n_282), .Y(n_341) );
AND2x2_ASAP7_75t_L g374 ( .A(n_170), .B(n_186), .Y(n_374) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
OR2x2_ASAP7_75t_L g281 ( .A(n_171), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g294 ( .A(n_171), .B(n_186), .Y(n_294) );
AND2x2_ASAP7_75t_L g301 ( .A(n_171), .B(n_282), .Y(n_301) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_171), .Y(n_310) );
AND2x2_ASAP7_75t_L g317 ( .A(n_171), .B(n_185), .Y(n_317) );
INVx1_ASAP7_75t_L g348 ( .A(n_171), .Y(n_348) );
OAI21xp5_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_176), .B(n_181), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_179), .A2(n_234), .B(n_235), .Y(n_233) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx4_ASAP7_75t_L g477 ( .A(n_180), .Y(n_477) );
NAND3xp33_ASAP7_75t_L g198 ( .A(n_181), .B(n_199), .C(n_202), .Y(n_198) );
INVx2_ASAP7_75t_L g213 ( .A(n_183), .Y(n_213) );
OA21x2_ASAP7_75t_L g216 ( .A1(n_183), .A2(n_217), .B(n_225), .Y(n_216) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_183), .A2(n_227), .B(n_236), .Y(n_226) );
INVx1_ASAP7_75t_L g494 ( .A(n_183), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_183), .A2(n_502), .B(n_503), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_183), .A2(n_526), .B(n_527), .Y(n_525) );
INVx1_ASAP7_75t_L g324 ( .A(n_184), .Y(n_324) );
AND2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_196), .Y(n_184) );
INVx2_ASAP7_75t_L g280 ( .A(n_185), .Y(n_280) );
AND2x2_ASAP7_75t_L g302 ( .A(n_185), .B(n_241), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_185), .B(n_348), .Y(n_353) );
INVx3_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_186), .B(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g425 ( .A(n_186), .B(n_389), .Y(n_425) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_195), .Y(n_186) );
INVx4_ASAP7_75t_L g202 ( .A(n_187), .Y(n_202) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_187), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_187), .A2(n_546), .B(n_547), .Y(n_545) );
INVx2_ASAP7_75t_L g239 ( .A(n_196), .Y(n_239) );
INVx3_ASAP7_75t_L g340 ( .A(n_196), .Y(n_340) );
OR2x2_ASAP7_75t_L g370 ( .A(n_196), .B(n_371), .Y(n_370) );
NOR2x1_ASAP7_75t_L g396 ( .A(n_196), .B(n_280), .Y(n_396) );
AND2x4_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
INVx1_ASAP7_75t_L g283 ( .A(n_197), .Y(n_283) );
AO21x1_ASAP7_75t_L g282 ( .A1(n_199), .A2(n_202), .B(n_283), .Y(n_282) );
AO21x2_ASAP7_75t_L g452 ( .A1(n_202), .A2(n_453), .B(n_466), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_202), .B(n_467), .Y(n_466) );
INVx3_ASAP7_75t_L g469 ( .A(n_202), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_202), .B(n_510), .Y(n_509) );
AO21x2_ASAP7_75t_L g514 ( .A1(n_202), .A2(n_515), .B(n_522), .Y(n_514) );
AOI33xp33_ASAP7_75t_L g416 ( .A1(n_203), .A2(n_254), .A3(n_268), .B1(n_340), .B2(n_417), .B3(n_418), .Y(n_416) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
OR2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_214), .Y(n_204) );
OR2x2_ASAP7_75t_L g269 ( .A(n_205), .B(n_270), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_205), .B(n_266), .Y(n_328) );
OR2x2_ASAP7_75t_L g381 ( .A(n_205), .B(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g307 ( .A(n_206), .B(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g332 ( .A(n_206), .B(n_214), .Y(n_332) );
AND2x2_ASAP7_75t_L g399 ( .A(n_206), .B(n_244), .Y(n_399) );
AOI21xp5_ASAP7_75t_L g424 ( .A1(n_206), .A2(n_299), .B(n_425), .Y(n_424) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g246 ( .A(n_207), .Y(n_246) );
INVx1_ASAP7_75t_L g259 ( .A(n_207), .Y(n_259) );
AND2x2_ASAP7_75t_L g278 ( .A(n_207), .B(n_248), .Y(n_278) );
AND2x2_ASAP7_75t_L g327 ( .A(n_207), .B(n_247), .Y(n_327) );
INVx2_ASAP7_75t_L g478 ( .A(n_211), .Y(n_478) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_211), .Y(n_508) );
INVx1_ASAP7_75t_L g491 ( .A(n_213), .Y(n_491) );
INVx2_ASAP7_75t_SL g369 ( .A(n_214), .Y(n_369) );
OR2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_226), .Y(n_214) );
INVx2_ASAP7_75t_L g289 ( .A(n_215), .Y(n_289) );
INVx1_ASAP7_75t_L g420 ( .A(n_215), .Y(n_420) );
AND2x2_ASAP7_75t_L g433 ( .A(n_215), .B(n_314), .Y(n_433) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g260 ( .A(n_216), .Y(n_260) );
OR2x2_ASAP7_75t_L g266 ( .A(n_216), .B(n_267), .Y(n_266) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_216), .Y(n_277) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_226), .Y(n_244) );
AND2x2_ASAP7_75t_L g261 ( .A(n_226), .B(n_247), .Y(n_261) );
INVx1_ASAP7_75t_L g267 ( .A(n_226), .Y(n_267) );
INVx1_ASAP7_75t_L g274 ( .A(n_226), .Y(n_274) );
AND2x2_ASAP7_75t_L g299 ( .A(n_226), .B(n_248), .Y(n_299) );
INVx2_ASAP7_75t_L g315 ( .A(n_226), .Y(n_315) );
AND2x2_ASAP7_75t_L g408 ( .A(n_226), .B(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_226), .B(n_289), .Y(n_429) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_231), .Y(n_228) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_SL g237 ( .A(n_238), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
INVx2_ASAP7_75t_L g263 ( .A(n_239), .Y(n_263) );
INVx1_ASAP7_75t_L g292 ( .A(n_239), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_239), .B(n_323), .Y(n_389) );
INVx1_ASAP7_75t_SL g349 ( .A(n_240), .Y(n_349) );
INVx2_ASAP7_75t_L g270 ( .A(n_241), .Y(n_270) );
AND2x2_ASAP7_75t_L g339 ( .A(n_241), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g355 ( .A(n_241), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_245), .Y(n_242) );
INVx1_ASAP7_75t_L g417 ( .A(n_243), .Y(n_417) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g272 ( .A(n_245), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g375 ( .A(n_245), .B(n_365), .Y(n_375) );
AOI21xp5_ASAP7_75t_L g427 ( .A1(n_245), .A2(n_386), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
AND2x2_ASAP7_75t_L g288 ( .A(n_246), .B(n_289), .Y(n_288) );
BUFx2_ASAP7_75t_L g313 ( .A(n_246), .Y(n_313) );
INVx1_ASAP7_75t_L g337 ( .A(n_246), .Y(n_337) );
OR2x2_ASAP7_75t_L g401 ( .A(n_247), .B(n_260), .Y(n_401) );
NOR2xp67_ASAP7_75t_L g409 ( .A(n_247), .B(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g314 ( .A(n_248), .B(n_315), .Y(n_314) );
BUFx2_ASAP7_75t_L g321 ( .A(n_248), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_255), .B1(n_262), .B2(n_264), .Y(n_252) );
OR2x2_ASAP7_75t_L g331 ( .A(n_253), .B(n_281), .Y(n_331) );
INVx1_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
AOI222xp33_ASAP7_75t_L g372 ( .A1(n_254), .A2(n_373), .B1(n_375), .B2(n_376), .C1(n_377), .C2(n_380), .Y(n_372) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_261), .Y(n_256) );
INVx1_ASAP7_75t_SL g257 ( .A(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g319 ( .A(n_258), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
AND2x2_ASAP7_75t_SL g273 ( .A(n_260), .B(n_274), .Y(n_273) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_260), .Y(n_344) );
AND2x2_ASAP7_75t_L g392 ( .A(n_260), .B(n_261), .Y(n_392) );
INVx1_ASAP7_75t_L g410 ( .A(n_260), .Y(n_410) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g376 ( .A(n_263), .B(n_302), .Y(n_376) );
AND2x2_ASAP7_75t_L g418 ( .A(n_263), .B(n_294), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_268), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_265), .B(n_313), .Y(n_400) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_266), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g293 ( .A(n_270), .B(n_294), .Y(n_293) );
INVx3_ASAP7_75t_L g361 ( .A(n_270), .Y(n_361) );
O2A1O1Ixp33_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_275), .B(n_279), .C(n_284), .Y(n_271) );
INVxp67_ASAP7_75t_L g285 ( .A(n_272), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_273), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_273), .B(n_320), .Y(n_415) );
BUFx3_ASAP7_75t_L g379 ( .A(n_274), .Y(n_379) );
INVx1_ASAP7_75t_L g286 ( .A(n_275), .Y(n_286) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g305 ( .A(n_277), .B(n_299), .Y(n_305) );
INVx1_ASAP7_75t_SL g345 ( .A(n_278), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g335 ( .A(n_280), .Y(n_335) );
AND2x2_ASAP7_75t_L g358 ( .A(n_280), .B(n_341), .Y(n_358) );
INVx1_ASAP7_75t_SL g329 ( .A(n_281), .Y(n_329) );
INVx1_ASAP7_75t_L g356 ( .A(n_282), .Y(n_356) );
AOI31xp33_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_286), .A3(n_287), .B(n_290), .Y(n_284) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g377 ( .A(n_288), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g351 ( .A(n_289), .Y(n_351) );
BUFx2_ASAP7_75t_L g365 ( .A(n_289), .Y(n_365) );
AND2x2_ASAP7_75t_L g393 ( .A(n_289), .B(n_314), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_SL g366 ( .A(n_293), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_294), .B(n_361), .Y(n_407) );
AND2x2_ASAP7_75t_L g414 ( .A(n_294), .B(n_340), .Y(n_414) );
AOI211xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_300), .B(n_303), .C(n_318), .Y(n_295) );
INVxp67_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AOI221xp5_ASAP7_75t_L g326 ( .A1(n_300), .A2(n_327), .B1(n_328), .B2(n_329), .C(n_330), .Y(n_326) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
AND2x2_ASAP7_75t_L g334 ( .A(n_301), .B(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g371 ( .A(n_302), .Y(n_371) );
OAI32xp33_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_306), .A3(n_309), .B1(n_311), .B2(n_316), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
O2A1O1Ixp33_ASAP7_75t_L g357 ( .A1(n_305), .A2(n_358), .B(n_359), .C(n_362), .Y(n_357) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
OAI21xp5_ASAP7_75t_SL g421 ( .A1(n_313), .A2(n_422), .B(n_423), .Y(n_421) );
INVx1_ASAP7_75t_L g382 ( .A(n_314), .Y(n_382) );
INVxp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_319), .B(n_322), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_320), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g368 ( .A(n_320), .B(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g385 ( .A(n_322), .Y(n_385) );
OR2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
NAND4xp25_ASAP7_75t_SL g325 ( .A(n_326), .B(n_338), .C(n_357), .D(n_372), .Y(n_325) );
AND2x2_ASAP7_75t_L g364 ( .A(n_327), .B(n_365), .Y(n_364) );
AND2x4_ASAP7_75t_L g386 ( .A(n_327), .B(n_379), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_329), .B(n_361), .Y(n_360) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_332), .B1(n_333), .B2(n_336), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_331), .A2(n_382), .B1(n_413), .B2(n_415), .Y(n_412) );
O2A1O1Ixp33_ASAP7_75t_L g419 ( .A1(n_331), .A2(n_420), .B(n_421), .C(n_424), .Y(n_419) );
INVx2_ASAP7_75t_L g390 ( .A(n_332), .Y(n_390) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AOI222xp33_ASAP7_75t_L g384 ( .A1(n_334), .A2(n_368), .B1(n_385), .B2(n_386), .C1(n_387), .C2(n_390), .Y(n_384) );
O2A1O1Ixp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_341), .B(n_342), .C(n_346), .Y(n_338) );
INVx1_ASAP7_75t_L g404 ( .A(n_339), .Y(n_404) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OAI22xp33_ASAP7_75t_L g346 ( .A1(n_343), .A2(n_347), .B1(n_350), .B2(n_352), .Y(n_346) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
OR2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g373 ( .A(n_355), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g431 ( .A(n_358), .Y(n_431) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OAI22xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_366), .B1(n_367), .B2(n_370), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_365), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g422 ( .A(n_370), .Y(n_422) );
INVx1_ASAP7_75t_L g403 ( .A(n_374), .Y(n_403) );
CKINVDCx16_ASAP7_75t_R g430 ( .A(n_376), .Y(n_430) );
INVxp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND5xp2_ASAP7_75t_L g383 ( .A(n_384), .B(n_391), .C(n_405), .D(n_411), .E(n_416), .Y(n_383) );
INVx1_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
O2A1O1Ixp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B(n_394), .C(n_397), .Y(n_391) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AOI31xp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_400), .A3(n_401), .B(n_402), .Y(n_397) );
INVx1_ASAP7_75t_L g423 ( .A(n_399), .Y(n_423) );
OR2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OAI222xp33_ASAP7_75t_L g426 ( .A1(n_413), .A2(n_415), .B1(n_427), .B2(n_430), .C1(n_431), .C2(n_432), .Y(n_426) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
NAND3xp33_ASAP7_75t_L g438 ( .A(n_435), .B(n_439), .C(n_732), .Y(n_438) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_444), .B1(n_445), .B2(n_447), .Y(n_441) );
INVx2_ASAP7_75t_L g730 ( .A(n_442), .Y(n_730) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OAI22xp5_ASAP7_75t_SL g729 ( .A1(n_444), .A2(n_447), .B1(n_730), .B2(n_731), .Y(n_729) );
INVx2_ASAP7_75t_L g731 ( .A(n_445), .Y(n_731) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OR3x1_ASAP7_75t_L g447 ( .A(n_448), .B(n_633), .C(n_682), .Y(n_447) );
NAND5xp2_ASAP7_75t_L g448 ( .A(n_449), .B(n_567), .C(n_596), .D(n_604), .E(n_619), .Y(n_448) );
O2A1O1Ixp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_495), .B(n_511), .C(n_551), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_451), .B(n_480), .Y(n_450) );
AND2x2_ASAP7_75t_L g562 ( .A(n_451), .B(n_559), .Y(n_562) );
AND2x2_ASAP7_75t_L g595 ( .A(n_451), .B(n_481), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_451), .B(n_499), .Y(n_688) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_468), .Y(n_451) );
INVx2_ASAP7_75t_L g498 ( .A(n_452), .Y(n_498) );
BUFx2_ASAP7_75t_L g662 ( .A(n_452), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_463), .Y(n_453) );
INVx5_ASAP7_75t_L g473 ( .A(n_455), .Y(n_473) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_SL g471 ( .A1(n_462), .A2(n_472), .B(n_473), .C(n_474), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g537 ( .A1(n_462), .A2(n_473), .B(n_538), .C(n_539), .Y(n_537) );
BUFx2_ASAP7_75t_L g484 ( .A(n_464), .Y(n_484) );
AND2x2_ASAP7_75t_L g480 ( .A(n_468), .B(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g560 ( .A(n_468), .Y(n_560) );
AND2x2_ASAP7_75t_L g646 ( .A(n_468), .B(n_559), .Y(n_646) );
AND2x2_ASAP7_75t_L g701 ( .A(n_468), .B(n_498), .Y(n_701) );
OA21x2_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_470), .B(n_479), .Y(n_468) );
INVx2_ASAP7_75t_L g504 ( .A(n_473), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
INVx1_ASAP7_75t_L g618 ( .A(n_480), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_480), .B(n_499), .Y(n_665) );
INVx5_ASAP7_75t_L g559 ( .A(n_481), .Y(n_559) );
AND2x4_ASAP7_75t_L g580 ( .A(n_481), .B(n_560), .Y(n_580) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_481), .Y(n_602) );
AND2x2_ASAP7_75t_L g677 ( .A(n_481), .B(n_662), .Y(n_677) );
AND2x2_ASAP7_75t_L g680 ( .A(n_481), .B(n_500), .Y(n_680) );
OR2x6_ASAP7_75t_L g481 ( .A(n_482), .B(n_492), .Y(n_481) );
AOI21xp5_ASAP7_75t_SL g482 ( .A1(n_483), .A2(n_485), .B(n_491), .Y(n_482) );
INVx2_ASAP7_75t_L g490 ( .A(n_488), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_L g505 ( .A1(n_490), .A2(n_506), .B(n_507), .C(n_508), .Y(n_505) );
O2A1O1Ixp33_ASAP7_75t_L g528 ( .A1(n_490), .A2(n_508), .B(n_529), .C(n_530), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_495), .B(n_560), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_495), .B(n_691), .Y(n_690) );
INVx2_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_499), .Y(n_496) );
AND2x2_ASAP7_75t_L g585 ( .A(n_497), .B(n_560), .Y(n_585) );
AND2x2_ASAP7_75t_L g603 ( .A(n_497), .B(n_500), .Y(n_603) );
INVx1_ASAP7_75t_L g623 ( .A(n_497), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_497), .B(n_559), .Y(n_668) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_497), .Y(n_710) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_498), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_499), .B(n_558), .Y(n_557) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_499), .Y(n_612) );
O2A1O1Ixp33_ASAP7_75t_L g615 ( .A1(n_499), .A2(n_555), .B(n_616), .C(n_618), .Y(n_615) );
AND2x2_ASAP7_75t_L g622 ( .A(n_499), .B(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g631 ( .A(n_499), .B(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g635 ( .A(n_499), .B(n_559), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_499), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g650 ( .A(n_499), .B(n_560), .Y(n_650) );
AND2x2_ASAP7_75t_L g700 ( .A(n_499), .B(n_701), .Y(n_700) );
INVx5_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx2_ASAP7_75t_L g564 ( .A(n_500), .Y(n_564) );
AND2x2_ASAP7_75t_L g605 ( .A(n_500), .B(n_558), .Y(n_605) );
AND2x2_ASAP7_75t_L g617 ( .A(n_500), .B(n_592), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_500), .B(n_646), .Y(n_664) );
OR2x6_ASAP7_75t_L g500 ( .A(n_501), .B(n_509), .Y(n_500) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_532), .Y(n_511) );
INVx1_ASAP7_75t_L g553 ( .A(n_512), .Y(n_553) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_524), .Y(n_512) );
OR2x2_ASAP7_75t_L g555 ( .A(n_513), .B(n_524), .Y(n_555) );
NAND3xp33_ASAP7_75t_L g561 ( .A(n_513), .B(n_562), .C(n_563), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_513), .B(n_534), .Y(n_572) );
OR2x2_ASAP7_75t_L g587 ( .A(n_513), .B(n_575), .Y(n_587) );
AND2x2_ASAP7_75t_L g593 ( .A(n_513), .B(n_543), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_513), .B(n_724), .Y(n_723) );
INVx5_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_514), .B(n_534), .Y(n_590) );
AND2x2_ASAP7_75t_L g629 ( .A(n_514), .B(n_544), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g657 ( .A(n_514), .B(n_543), .Y(n_657) );
OR2x2_ASAP7_75t_L g660 ( .A(n_514), .B(n_543), .Y(n_660) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_517), .B(n_518), .Y(n_515) );
INVx5_ASAP7_75t_SL g575 ( .A(n_524), .Y(n_575) );
OR2x2_ASAP7_75t_L g581 ( .A(n_524), .B(n_533), .Y(n_581) );
AND2x2_ASAP7_75t_L g597 ( .A(n_524), .B(n_598), .Y(n_597) );
AOI321xp33_ASAP7_75t_L g604 ( .A1(n_524), .A2(n_605), .A3(n_606), .B1(n_607), .B2(n_613), .C(n_615), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_524), .B(n_532), .Y(n_614) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_524), .Y(n_627) );
OR2x2_ASAP7_75t_L g674 ( .A(n_524), .B(n_572), .Y(n_674) );
AND2x2_ASAP7_75t_L g696 ( .A(n_524), .B(n_593), .Y(n_696) );
AND2x2_ASAP7_75t_L g715 ( .A(n_524), .B(n_534), .Y(n_715) );
OR2x6_ASAP7_75t_L g524 ( .A(n_525), .B(n_531), .Y(n_524) );
INVx1_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_543), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_534), .B(n_543), .Y(n_556) );
AND2x2_ASAP7_75t_L g565 ( .A(n_534), .B(n_566), .Y(n_565) );
INVx3_ASAP7_75t_L g592 ( .A(n_534), .Y(n_592) );
AND2x2_ASAP7_75t_L g598 ( .A(n_534), .B(n_593), .Y(n_598) );
INVxp67_ASAP7_75t_L g628 ( .A(n_534), .Y(n_628) );
OR2x2_ASAP7_75t_L g670 ( .A(n_534), .B(n_575), .Y(n_670) );
OA21x2_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_536), .B(n_542), .Y(n_534) );
OR2x2_ASAP7_75t_L g552 ( .A(n_543), .B(n_553), .Y(n_552) );
INVx1_ASAP7_75t_SL g566 ( .A(n_543), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_543), .B(n_555), .Y(n_599) );
AND2x2_ASAP7_75t_L g648 ( .A(n_543), .B(n_592), .Y(n_648) );
AND2x2_ASAP7_75t_L g686 ( .A(n_543), .B(n_575), .Y(n_686) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_544), .B(n_575), .Y(n_574) );
A2O1A1Ixp33_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_554), .B(n_557), .C(n_561), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_552), .A2(n_554), .B1(n_679), .B2(n_681), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_554), .A2(n_577), .B1(n_632), .B2(n_718), .Y(n_717) );
OR2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
INVx1_ASAP7_75t_SL g706 ( .A(n_555), .Y(n_706) );
INVx1_ASAP7_75t_SL g606 ( .A(n_556), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_558), .B(n_578), .Y(n_608) );
AOI222xp33_ASAP7_75t_L g619 ( .A1(n_558), .A2(n_599), .B1(n_606), .B2(n_620), .C1(n_624), .C2(n_630), .Y(n_619) );
AND2x2_ASAP7_75t_L g709 ( .A(n_558), .B(n_710), .Y(n_709) );
AND2x4_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
INVx2_ASAP7_75t_L g584 ( .A(n_559), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_559), .B(n_579), .Y(n_654) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_559), .Y(n_691) );
AND2x2_ASAP7_75t_L g694 ( .A(n_559), .B(n_603), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_559), .B(n_710), .Y(n_720) );
INVx1_ASAP7_75t_L g611 ( .A(n_560), .Y(n_611) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_560), .Y(n_639) );
O2A1O1Ixp33_ASAP7_75t_L g702 ( .A1(n_562), .A2(n_703), .B(n_704), .C(n_707), .Y(n_702) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
NAND3xp33_ASAP7_75t_L g625 ( .A(n_564), .B(n_626), .C(n_629), .Y(n_625) );
OR2x2_ASAP7_75t_L g653 ( .A(n_564), .B(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_564), .B(n_580), .Y(n_681) );
OR2x2_ASAP7_75t_L g586 ( .A(n_566), .B(n_587), .Y(n_586) );
AOI211xp5_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_570), .B(n_576), .C(n_588), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_569), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g675 ( .A(n_570), .B(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_571), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g589 ( .A(n_574), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_575), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g643 ( .A(n_575), .B(n_593), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_575), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_575), .B(n_592), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_581), .B1(n_582), .B2(n_586), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_578), .B(n_650), .Y(n_649) );
BUFx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_580), .B(n_622), .Y(n_621) );
OAI221xp5_ASAP7_75t_SL g644 ( .A1(n_581), .A2(n_645), .B1(n_647), .B2(n_649), .C(n_651), .Y(n_644) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
AND2x2_ASAP7_75t_L g699 ( .A(n_584), .B(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g712 ( .A(n_584), .B(n_701), .Y(n_712) );
INVx1_ASAP7_75t_L g632 ( .A(n_585), .Y(n_632) );
INVx1_ASAP7_75t_L g703 ( .A(n_586), .Y(n_703) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_587), .A2(n_670), .B(n_693), .Y(n_692) );
AOI21xp33_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_591), .B(n_594), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OAI21xp5_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_599), .B(n_600), .Y(n_596) );
INVx1_ASAP7_75t_L g636 ( .A(n_597), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_598), .A2(n_684), .B1(n_687), .B2(n_689), .C(n_692), .Y(n_683) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_606), .A2(n_696), .B1(n_697), .B2(n_699), .Y(n_695) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_608), .B(n_609), .Y(n_607) );
INVx1_ASAP7_75t_L g672 ( .A(n_608), .Y(n_672) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NOR2xp67_ASAP7_75t_SL g610 ( .A(n_611), .B(n_612), .Y(n_610) );
AND2x2_ASAP7_75t_L g676 ( .A(n_612), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g641 ( .A(n_617), .Y(n_641) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_622), .B(n_646), .Y(n_698) );
INVxp67_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_628), .B(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g714 ( .A(n_629), .B(n_715), .Y(n_714) );
AND2x4_ASAP7_75t_L g721 ( .A(n_629), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OAI211xp5_ASAP7_75t_SL g633 ( .A1(n_634), .A2(n_636), .B(n_637), .C(n_671), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AOI211xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_640), .B(n_644), .C(n_663), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_SL g724 ( .A(n_648), .Y(n_724) );
AND2x2_ASAP7_75t_L g661 ( .A(n_650), .B(n_662), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_655), .B1(n_659), .B2(n_661), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OR2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
OR2x2_ASAP7_75t_L g669 ( .A(n_657), .B(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g722 ( .A(n_658), .Y(n_722) );
INVxp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AOI31xp33_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .A3(n_666), .B(n_669), .Y(n_663) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AOI211xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .B(n_675), .C(n_678), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
CKINVDCx16_ASAP7_75t_R g679 ( .A(n_680), .Y(n_679) );
NAND5xp2_ASAP7_75t_L g682 ( .A(n_683), .B(n_695), .C(n_702), .D(n_716), .E(n_719), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_694), .A2(n_720), .B1(n_721), .B2(n_723), .Y(n_719) );
INVx1_ASAP7_75t_SL g718 ( .A(n_696), .Y(n_718) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AOI21xp33_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_711), .B(n_713), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVxp67_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
endmodule