module fake_jpeg_2195_n_288 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_288);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_118;
wire n_128;
wire n_82;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_15),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_45),
.B(n_53),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_46),
.B(n_33),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx2_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_61),
.Y(n_92)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_18),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_18),
.B(n_15),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_13),
.Y(n_90)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_22),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

NAND3xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_33),
.C(n_31),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_70),
.B(n_77),
.Y(n_119)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_73),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_52),
.B(n_37),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_83),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_91),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_37),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_59),
.B(n_20),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_97),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_34),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_105),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_46),
.B(n_20),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_26),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_100),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_47),
.A2(n_23),
.B1(n_30),
.B2(n_28),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g136 ( 
.A1(n_99),
.A2(n_22),
.B1(n_29),
.B2(n_57),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_34),
.Y(n_100)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

CKINVDCx12_ASAP7_75t_R g104 ( 
.A(n_51),
.Y(n_104)
);

BUFx4f_ASAP7_75t_SL g141 ( 
.A(n_104),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_31),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_69),
.A2(n_30),
.B1(n_21),
.B2(n_26),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_106),
.A2(n_69),
.B1(n_58),
.B2(n_65),
.Y(n_120)
);

INVx6_ASAP7_75t_SL g107 ( 
.A(n_51),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_107),
.Y(n_112)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_92),
.A2(n_44),
.B1(n_48),
.B2(n_61),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_111),
.A2(n_117),
.B1(n_131),
.B2(n_133),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_50),
.B(n_64),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_113),
.A2(n_135),
.B(n_144),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_70),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_114),
.B(n_140),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_99),
.A2(n_49),
.B1(n_68),
.B2(n_43),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_120),
.A2(n_125),
.B1(n_127),
.B2(n_128),
.Y(n_171)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_76),
.A2(n_60),
.B1(n_66),
.B2(n_41),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_126),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_28),
.B1(n_41),
.B2(n_21),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_87),
.A2(n_41),
.B1(n_19),
.B2(n_27),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_129),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_87),
.A2(n_19),
.B1(n_27),
.B2(n_36),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_72),
.A2(n_78),
.B1(n_108),
.B2(n_103),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_132),
.A2(n_144),
.B1(n_81),
.B2(n_24),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_72),
.A2(n_27),
.B1(n_36),
.B2(n_24),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_88),
.B(n_27),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_102),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_79),
.B(n_50),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_135),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_139),
.Y(n_151)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_71),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_109),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_142),
.B(n_143),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_109),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_78),
.A2(n_24),
.B1(n_22),
.B2(n_29),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_86),
.B(n_0),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_0),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_114),
.A2(n_102),
.B(n_79),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_154),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_85),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_156),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_95),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_113),
.A2(n_85),
.B(n_101),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_164),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_88),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_157),
.B(n_165),
.Y(n_194)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_158),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_108),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_160),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_112),
.A2(n_84),
.B(n_73),
.Y(n_160)
);

BUFx24_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

INVx13_ASAP7_75t_L g200 ( 
.A(n_162),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_84),
.C(n_103),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_121),
.B(n_80),
.C(n_110),
.Y(n_165)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

O2A1O1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_112),
.A2(n_24),
.B(n_81),
.C(n_80),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_172),
.Y(n_190)
);

AO21x2_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_117),
.B(n_120),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_141),
.Y(n_170)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_130),
.B(n_1),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_141),
.Y(n_176)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_176),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_191),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_153),
.A2(n_131),
.B1(n_128),
.B2(n_134),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_174),
.A2(n_143),
.B1(n_136),
.B2(n_129),
.Y(n_179)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_151),
.A2(n_136),
.B1(n_133),
.B2(n_135),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_189),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_149),
.A2(n_136),
.B1(n_124),
.B2(n_118),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_171),
.A2(n_115),
.B1(n_139),
.B2(n_140),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_193),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_151),
.A2(n_115),
.B1(n_122),
.B2(n_138),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_151),
.A2(n_137),
.B1(n_24),
.B2(n_5),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_195),
.Y(n_204)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_163),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_197),
.B(n_199),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_12),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_172),
.Y(n_210)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_167),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_207),
.Y(n_229)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

OAI32xp33_ASAP7_75t_L g207 ( 
.A1(n_180),
.A2(n_159),
.A3(n_150),
.B1(n_165),
.B2(n_164),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_SL g208 ( 
.A1(n_185),
.A2(n_190),
.B(n_182),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_208),
.A2(n_219),
.B(n_222),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_217),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_154),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_213),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_161),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_175),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_200),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_220),
.Y(n_234)
);

AOI21x1_ASAP7_75t_L g219 ( 
.A1(n_186),
.A2(n_147),
.B(n_155),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_146),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_179),
.A2(n_152),
.B1(n_169),
.B2(n_168),
.Y(n_221)
);

AO21x1_ASAP7_75t_L g232 ( 
.A1(n_221),
.A2(n_185),
.B(n_186),
.Y(n_232)
);

A2O1A1O1Ixp25_ASAP7_75t_L g222 ( 
.A1(n_183),
.A2(n_160),
.B(n_162),
.C(n_146),
.D(n_166),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_158),
.Y(n_223)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_223),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_196),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_224),
.Y(n_226)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

AOI21x1_ASAP7_75t_L g250 ( 
.A1(n_232),
.A2(n_233),
.B(n_204),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_219),
.A2(n_183),
.B(n_193),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_217),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_235),
.B(n_228),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_212),
.A2(n_191),
.B(n_190),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_236),
.A2(n_241),
.B(n_209),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_189),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_204),
.C(n_221),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_216),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_216),
.Y(n_246)
);

AOI322xp5_ASAP7_75t_L g239 ( 
.A1(n_209),
.A2(n_177),
.A3(n_203),
.B1(n_195),
.B2(n_192),
.C1(n_200),
.C2(n_201),
.Y(n_239)
);

AOI322xp5_ASAP7_75t_L g253 ( 
.A1(n_239),
.A2(n_214),
.A3(n_224),
.B1(n_177),
.B2(n_162),
.C1(n_201),
.C2(n_196),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_222),
.A2(n_203),
.B(n_162),
.Y(n_241)
);

NAND3xp33_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_251),
.C(n_231),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_234),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_243),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_244),
.A2(n_247),
.B1(n_252),
.B2(n_253),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_250),
.Y(n_256)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_227),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_223),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_249),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_226),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_229),
.A2(n_177),
.B1(n_214),
.B2(n_210),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_237),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_257),
.B(n_258),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_225),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_233),
.C(n_230),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_260),
.B(n_262),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_261),
.A2(n_225),
.B1(n_242),
.B2(n_240),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_230),
.C(n_238),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_245),
.C(n_252),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_241),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_264),
.B(n_267),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_259),
.A2(n_250),
.B1(n_244),
.B2(n_251),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_266),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_227),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_268),
.B(n_269),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_240),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_236),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_1),
.Y(n_277)
);

AOI322xp5_ASAP7_75t_L g273 ( 
.A1(n_265),
.A2(n_232),
.A3(n_254),
.B1(n_257),
.B2(n_260),
.C1(n_256),
.C2(n_177),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_273),
.A2(n_274),
.B1(n_266),
.B2(n_7),
.Y(n_280)
);

AOI322xp5_ASAP7_75t_L g274 ( 
.A1(n_270),
.A2(n_254),
.A3(n_148),
.B1(n_5),
.B2(n_7),
.C1(n_8),
.C2(n_1),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_277),
.B(n_4),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_268),
.Y(n_278)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_278),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_279),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_281),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_276),
.A2(n_4),
.B(n_8),
.Y(n_281)
);

O2A1O1Ixp33_ASAP7_75t_L g285 ( 
.A1(n_282),
.A2(n_275),
.B(n_8),
.C(n_9),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_286),
.Y(n_287)
);

AOI322xp5_ASAP7_75t_L g286 ( 
.A1(n_284),
.A2(n_4),
.A3(n_10),
.B1(n_11),
.B2(n_275),
.C1(n_282),
.C2(n_276),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_283),
.Y(n_288)
);


endmodule