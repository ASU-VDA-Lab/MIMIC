module real_aes_7033_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_551;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_725;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_0), .B(n_88), .C(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g127 ( .A(n_0), .Y(n_127) );
A2O1A1Ixp33_ASAP7_75t_L g466 ( .A1(n_1), .A2(n_155), .B(n_167), .C(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g274 ( .A(n_2), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_3), .A2(n_182), .B(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_4), .B(n_178), .Y(n_511) );
AOI21xp33_ASAP7_75t_L g181 ( .A1(n_5), .A2(n_182), .B(n_183), .Y(n_181) );
AND2x6_ASAP7_75t_L g155 ( .A(n_6), .B(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_7), .A2(n_250), .B(n_251), .Y(n_249) );
INVx1_ASAP7_75t_L g110 ( .A(n_8), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_8), .B(n_41), .Y(n_128) );
INVx1_ASAP7_75t_L g482 ( .A(n_9), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_10), .B(n_188), .Y(n_470) );
INVx1_ASAP7_75t_L g190 ( .A(n_11), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_12), .B(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g152 ( .A(n_13), .Y(n_152) );
INVx1_ASAP7_75t_L g256 ( .A(n_14), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_15), .A2(n_191), .B(n_257), .C(n_491), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g132 ( .A1(n_16), .A2(n_133), .B1(n_134), .B2(n_135), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_16), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_17), .B(n_178), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_18), .B(n_201), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_19), .B(n_182), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_20), .B(n_524), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_21), .A2(n_158), .B(n_242), .C(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_22), .B(n_178), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_23), .B(n_188), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_24), .A2(n_254), .B(n_255), .C(n_257), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_25), .B(n_188), .Y(n_532) );
CKINVDCx16_ASAP7_75t_R g541 ( .A(n_26), .Y(n_541) );
INVx1_ASAP7_75t_L g531 ( .A(n_27), .Y(n_531) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_28), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_29), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_30), .B(n_188), .Y(n_275) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_31), .A2(n_66), .B1(n_738), .B2(n_739), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_31), .Y(n_739) );
INVx1_ASAP7_75t_L g520 ( .A(n_32), .Y(n_520) );
INVx1_ASAP7_75t_L g166 ( .A(n_33), .Y(n_166) );
INVx2_ASAP7_75t_L g160 ( .A(n_34), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_35), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_36), .A2(n_192), .B(n_242), .C(n_509), .Y(n_508) );
INVxp67_ASAP7_75t_L g521 ( .A(n_37), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_38), .A2(n_155), .B(n_167), .C(n_212), .Y(n_211) );
CKINVDCx14_ASAP7_75t_R g507 ( .A(n_39), .Y(n_507) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_40), .A2(n_167), .B(n_530), .C(n_534), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_41), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g164 ( .A(n_42), .Y(n_164) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_43), .A2(n_187), .B(n_217), .C(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_44), .B(n_188), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_45), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_46), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_47), .Y(n_517) );
INVx1_ASAP7_75t_L g497 ( .A(n_48), .Y(n_497) );
CKINVDCx16_ASAP7_75t_R g170 ( .A(n_49), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_50), .B(n_182), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g157 ( .A1(n_51), .A2(n_158), .B1(n_161), .B2(n_167), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_52), .Y(n_221) );
CKINVDCx16_ASAP7_75t_R g271 ( .A(n_53), .Y(n_271) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_54), .A2(n_187), .B(n_189), .C(n_192), .Y(n_186) );
CKINVDCx14_ASAP7_75t_R g479 ( .A(n_55), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g231 ( .A(n_56), .Y(n_231) );
INVx1_ASAP7_75t_L g184 ( .A(n_57), .Y(n_184) );
OAI22xp5_ASAP7_75t_SL g735 ( .A1(n_58), .A2(n_736), .B1(n_737), .B2(n_740), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_58), .Y(n_740) );
INVx1_ASAP7_75t_L g156 ( .A(n_59), .Y(n_156) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_60), .A2(n_104), .B1(n_115), .B2(n_742), .Y(n_103) );
OAI22xp5_ASAP7_75t_L g135 ( .A1(n_61), .A2(n_77), .B1(n_136), .B2(n_137), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_61), .Y(n_137) );
INVx1_ASAP7_75t_L g151 ( .A(n_62), .Y(n_151) );
INVx1_ASAP7_75t_SL g510 ( .A(n_63), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_64), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_65), .B(n_178), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_66), .Y(n_738) );
INVx1_ASAP7_75t_L g544 ( .A(n_67), .Y(n_544) );
A2O1A1Ixp33_ASAP7_75t_SL g200 ( .A1(n_68), .A2(n_192), .B(n_201), .C(n_202), .Y(n_200) );
INVxp67_ASAP7_75t_L g203 ( .A(n_69), .Y(n_203) );
INVx1_ASAP7_75t_L g114 ( .A(n_70), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_71), .A2(n_182), .B(n_478), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_72), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_73), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_74), .A2(n_182), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g224 ( .A(n_75), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_76), .A2(n_250), .B(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_77), .Y(n_136) );
INVx1_ASAP7_75t_L g489 ( .A(n_78), .Y(n_489) );
CKINVDCx16_ASAP7_75t_R g528 ( .A(n_79), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_80), .A2(n_155), .B(n_167), .C(n_226), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_81), .A2(n_182), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g492 ( .A(n_82), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_83), .B(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g149 ( .A(n_84), .Y(n_149) );
INVx1_ASAP7_75t_L g468 ( .A(n_85), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_86), .B(n_201), .Y(n_215) );
A2O1A1Ixp33_ASAP7_75t_L g272 ( .A1(n_87), .A2(n_155), .B(n_167), .C(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g124 ( .A(n_88), .B(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g455 ( .A(n_88), .Y(n_455) );
OR2x2_ASAP7_75t_L g723 ( .A(n_88), .B(n_126), .Y(n_723) );
A2O1A1Ixp33_ASAP7_75t_L g542 ( .A1(n_89), .A2(n_167), .B(n_543), .C(n_546), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_90), .B(n_195), .Y(n_194) );
AOI222xp33_ASAP7_75t_SL g130 ( .A1(n_91), .A2(n_131), .B1(n_132), .B2(n_138), .C1(n_724), .C2(n_728), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g278 ( .A(n_92), .Y(n_278) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_93), .A2(n_155), .B(n_167), .C(n_239), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g246 ( .A(n_94), .Y(n_246) );
INVx1_ASAP7_75t_L g199 ( .A(n_95), .Y(n_199) );
CKINVDCx16_ASAP7_75t_R g252 ( .A(n_96), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_97), .B(n_214), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_98), .B(n_180), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_99), .B(n_180), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_100), .B(n_114), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_101), .A2(n_182), .B(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g500 ( .A(n_102), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
CKINVDCx6p67_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_107), .Y(n_743) );
CKINVDCx9p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AOI22xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_130), .B1(n_731), .B2(n_732), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_118), .B(n_122), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_SL g731 ( .A(n_120), .Y(n_731) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g732 ( .A1(n_122), .A2(n_733), .B(n_741), .Y(n_732) );
NOR2xp33_ASAP7_75t_SL g122 ( .A(n_123), .B(n_129), .Y(n_122) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_124), .Y(n_741) );
NOR2x2_ASAP7_75t_L g730 ( .A(n_125), .B(n_455), .Y(n_730) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g454 ( .A(n_126), .B(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
CKINVDCx14_ASAP7_75t_R g134 ( .A(n_135), .Y(n_134) );
OAI22xp5_ASAP7_75t_SL g138 ( .A1(n_139), .A2(n_452), .B1(n_456), .B2(n_723), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OAI22xp5_ASAP7_75t_SL g724 ( .A1(n_140), .A2(n_452), .B1(n_725), .B2(n_726), .Y(n_724) );
AND3x1_ASAP7_75t_L g140 ( .A(n_141), .B(n_377), .C(n_426), .Y(n_140) );
NOR3xp33_ASAP7_75t_SL g141 ( .A(n_142), .B(n_284), .C(n_322), .Y(n_141) );
OAI222xp33_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_205), .B1(n_259), .B2(n_265), .C1(n_279), .C2(n_282), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_176), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_144), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_144), .B(n_327), .Y(n_418) );
BUFx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OR2x2_ASAP7_75t_L g295 ( .A(n_145), .B(n_196), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_145), .B(n_177), .Y(n_303) );
AND2x2_ASAP7_75t_L g338 ( .A(n_145), .B(n_315), .Y(n_338) );
OR2x2_ASAP7_75t_L g362 ( .A(n_145), .B(n_177), .Y(n_362) );
OR2x2_ASAP7_75t_L g370 ( .A(n_145), .B(n_269), .Y(n_370) );
AND2x2_ASAP7_75t_L g373 ( .A(n_145), .B(n_196), .Y(n_373) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
OR2x2_ASAP7_75t_L g267 ( .A(n_146), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g281 ( .A(n_146), .B(n_196), .Y(n_281) );
AND2x2_ASAP7_75t_L g331 ( .A(n_146), .B(n_269), .Y(n_331) );
AND2x2_ASAP7_75t_L g344 ( .A(n_146), .B(n_177), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_146), .B(n_430), .Y(n_451) );
AO21x2_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_153), .B(n_174), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_147), .B(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g219 ( .A(n_147), .Y(n_219) );
AO21x2_ASAP7_75t_L g269 ( .A1(n_147), .A2(n_270), .B(n_277), .Y(n_269) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_148), .Y(n_180) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
AND2x2_ASAP7_75t_SL g195 ( .A(n_149), .B(n_150), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
OAI22xp33_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_157), .B1(n_170), .B2(n_171), .Y(n_153) );
O2A1O1Ixp33_ASAP7_75t_L g183 ( .A1(n_154), .A2(n_184), .B(n_185), .C(n_186), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g198 ( .A1(n_154), .A2(n_185), .B(n_199), .C(n_200), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_L g251 ( .A1(n_154), .A2(n_185), .B(n_252), .C(n_253), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_SL g478 ( .A1(n_154), .A2(n_185), .B(n_479), .C(n_480), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_SL g488 ( .A1(n_154), .A2(n_185), .B(n_489), .C(n_490), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_SL g496 ( .A1(n_154), .A2(n_185), .B(n_497), .C(n_498), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_L g506 ( .A1(n_154), .A2(n_185), .B(n_507), .C(n_508), .Y(n_506) );
O2A1O1Ixp33_ASAP7_75t_SL g516 ( .A1(n_154), .A2(n_185), .B(n_517), .C(n_518), .Y(n_516) );
INVx1_ASAP7_75t_L g546 ( .A(n_154), .Y(n_546) );
INVx4_ASAP7_75t_SL g154 ( .A(n_155), .Y(n_154) );
NAND2x1p5_ASAP7_75t_L g171 ( .A(n_155), .B(n_172), .Y(n_171) );
AND2x4_ASAP7_75t_L g182 ( .A(n_155), .B(n_172), .Y(n_182) );
BUFx3_ASAP7_75t_L g534 ( .A(n_155), .Y(n_534) );
INVx2_ASAP7_75t_L g276 ( .A(n_158), .Y(n_276) );
INVx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g168 ( .A(n_160), .Y(n_168) );
INVx1_ASAP7_75t_L g173 ( .A(n_160), .Y(n_173) );
OAI22xp5_ASAP7_75t_SL g161 ( .A1(n_162), .A2(n_164), .B1(n_165), .B2(n_166), .Y(n_161) );
INVx2_ASAP7_75t_L g165 ( .A(n_162), .Y(n_165) );
INVx4_ASAP7_75t_L g254 ( .A(n_162), .Y(n_254) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g169 ( .A(n_163), .Y(n_169) );
AND2x2_ASAP7_75t_L g172 ( .A(n_163), .B(n_173), .Y(n_172) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_163), .Y(n_188) );
INVx3_ASAP7_75t_L g191 ( .A(n_163), .Y(n_191) );
INVx1_ASAP7_75t_L g201 ( .A(n_163), .Y(n_201) );
INVx2_ASAP7_75t_L g469 ( .A(n_165), .Y(n_469) );
INVx5_ASAP7_75t_L g185 ( .A(n_167), .Y(n_185) );
AND2x6_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_168), .Y(n_193) );
BUFx3_ASAP7_75t_L g218 ( .A(n_168), .Y(n_218) );
OAI21xp5_ASAP7_75t_L g223 ( .A1(n_171), .A2(n_224), .B(n_225), .Y(n_223) );
OAI21xp5_ASAP7_75t_L g270 ( .A1(n_171), .A2(n_271), .B(n_272), .Y(n_270) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_171), .A2(n_465), .B(n_466), .Y(n_464) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_171), .A2(n_195), .B(n_528), .C(n_529), .Y(n_527) );
OAI21xp5_ASAP7_75t_L g540 ( .A1(n_171), .A2(n_541), .B(n_542), .Y(n_540) );
INVx1_ASAP7_75t_L g522 ( .A(n_173), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_L g369 ( .A1(n_176), .A2(n_370), .B(n_371), .C(n_374), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_176), .B(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_176), .B(n_314), .Y(n_436) );
AND2x2_ASAP7_75t_L g176 ( .A(n_177), .B(n_196), .Y(n_176) );
AND2x2_ASAP7_75t_SL g280 ( .A(n_177), .B(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g294 ( .A(n_177), .Y(n_294) );
AND2x2_ASAP7_75t_L g321 ( .A(n_177), .B(n_315), .Y(n_321) );
INVx1_ASAP7_75t_SL g329 ( .A(n_177), .Y(n_329) );
AND2x2_ASAP7_75t_L g352 ( .A(n_177), .B(n_353), .Y(n_352) );
BUFx2_ASAP7_75t_L g430 ( .A(n_177), .Y(n_430) );
OA21x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_181), .B(n_194), .Y(n_177) );
INVx3_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_SL g220 ( .A(n_179), .B(n_221), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_179), .B(n_472), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_179), .B(n_536), .Y(n_535) );
AO21x2_ASAP7_75t_L g539 ( .A1(n_179), .A2(n_540), .B(n_547), .Y(n_539) );
INVx4_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
OA21x2_ASAP7_75t_L g196 ( .A1(n_180), .A2(n_197), .B(n_204), .Y(n_196) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_180), .Y(n_486) );
BUFx2_ASAP7_75t_L g250 ( .A(n_182), .Y(n_250) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx4_ASAP7_75t_L g242 ( .A(n_188), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_191), .B(n_203), .Y(n_202) );
INVx5_ASAP7_75t_L g214 ( .A(n_191), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_191), .B(n_482), .Y(n_481) );
INVx3_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_193), .Y(n_243) );
INVx1_ASAP7_75t_L g232 ( .A(n_195), .Y(n_232) );
INVx2_ASAP7_75t_L g236 ( .A(n_195), .Y(n_236) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_195), .A2(n_249), .B(n_258), .Y(n_248) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_195), .A2(n_477), .B(n_483), .Y(n_476) );
BUFx2_ASAP7_75t_L g266 ( .A(n_196), .Y(n_266) );
INVx1_ASAP7_75t_L g328 ( .A(n_196), .Y(n_328) );
INVx3_ASAP7_75t_L g353 ( .A(n_196), .Y(n_353) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_205), .B(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_233), .Y(n_205) );
INVx1_ASAP7_75t_L g349 ( .A(n_206), .Y(n_349) );
OAI32xp33_ASAP7_75t_L g355 ( .A1(n_206), .A2(n_294), .A3(n_356), .B1(n_357), .B2(n_358), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_206), .A2(n_360), .B1(n_363), .B2(n_368), .Y(n_359) );
INVx4_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g297 ( .A(n_207), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g375 ( .A(n_207), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g445 ( .A(n_207), .B(n_391), .Y(n_445) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_222), .Y(n_207) );
AND2x2_ASAP7_75t_L g260 ( .A(n_208), .B(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g290 ( .A(n_208), .Y(n_290) );
INVx1_ASAP7_75t_L g309 ( .A(n_208), .Y(n_309) );
OR2x2_ASAP7_75t_L g317 ( .A(n_208), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g324 ( .A(n_208), .B(n_298), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_208), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g345 ( .A(n_208), .B(n_263), .Y(n_345) );
INVx3_ASAP7_75t_L g367 ( .A(n_208), .Y(n_367) );
AND2x2_ASAP7_75t_L g392 ( .A(n_208), .B(n_264), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_208), .B(n_357), .Y(n_440) );
OR2x6_ASAP7_75t_L g208 ( .A(n_209), .B(n_220), .Y(n_208) );
AOI21xp5_ASAP7_75t_SL g209 ( .A1(n_210), .A2(n_211), .B(n_219), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_215), .B(n_216), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g273 ( .A1(n_214), .A2(n_274), .B(n_275), .C(n_276), .Y(n_273) );
OAI22xp33_ASAP7_75t_L g519 ( .A1(n_214), .A2(n_254), .B1(n_520), .B2(n_521), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_214), .A2(n_531), .B(n_532), .C(n_533), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_216), .A2(n_227), .B(n_228), .Y(n_226) );
O2A1O1Ixp5_ASAP7_75t_L g467 ( .A1(n_216), .A2(n_468), .B(n_469), .C(n_470), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_L g543 ( .A1(n_216), .A2(n_469), .B(n_544), .C(n_545), .Y(n_543) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g257 ( .A(n_218), .Y(n_257) );
INVx1_ASAP7_75t_L g229 ( .A(n_219), .Y(n_229) );
INVx2_ASAP7_75t_L g264 ( .A(n_222), .Y(n_264) );
AND2x2_ASAP7_75t_L g396 ( .A(n_222), .B(n_234), .Y(n_396) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_229), .B(n_230), .Y(n_222) );
INVx1_ASAP7_75t_L g514 ( .A(n_229), .Y(n_514) );
AO21x2_ASAP7_75t_L g566 ( .A1(n_229), .A2(n_567), .B(n_568), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_232), .B(n_246), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_232), .B(n_278), .Y(n_277) );
AO21x2_ASAP7_75t_L g463 ( .A1(n_232), .A2(n_464), .B(n_471), .Y(n_463) );
INVx2_ASAP7_75t_L g438 ( .A(n_233), .Y(n_438) );
OR2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_247), .Y(n_233) );
INVx1_ASAP7_75t_L g283 ( .A(n_234), .Y(n_283) );
AND2x2_ASAP7_75t_L g310 ( .A(n_234), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_234), .B(n_264), .Y(n_318) );
AND2x2_ASAP7_75t_L g376 ( .A(n_234), .B(n_299), .Y(n_376) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g262 ( .A(n_235), .Y(n_262) );
AND2x2_ASAP7_75t_L g289 ( .A(n_235), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g298 ( .A(n_235), .B(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_235), .B(n_264), .Y(n_364) );
AO21x2_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_245), .Y(n_235) );
INVx1_ASAP7_75t_L g524 ( .A(n_236), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_236), .B(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_244), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B(n_243), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_242), .B(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_247), .B(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g311 ( .A(n_247), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_247), .B(n_264), .Y(n_357) );
AND2x2_ASAP7_75t_L g366 ( .A(n_247), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g391 ( .A(n_247), .Y(n_391) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g263 ( .A(n_248), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g299 ( .A(n_248), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_254), .B(n_256), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_254), .B(n_492), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_254), .B(n_500), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_259), .A2(n_269), .B1(n_428), .B2(n_431), .Y(n_427) );
INVx1_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
OAI21xp5_ASAP7_75t_SL g450 ( .A1(n_261), .A2(n_372), .B(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_262), .B(n_367), .Y(n_384) );
INVx1_ASAP7_75t_L g409 ( .A(n_262), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_263), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g336 ( .A(n_263), .B(n_289), .Y(n_336) );
INVx2_ASAP7_75t_L g292 ( .A(n_264), .Y(n_292) );
INVx1_ASAP7_75t_L g342 ( .A(n_264), .Y(n_342) );
OAI221xp5_ASAP7_75t_L g433 ( .A1(n_265), .A2(n_417), .B1(n_434), .B2(n_437), .C(n_439), .Y(n_433) );
OR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx1_ASAP7_75t_L g304 ( .A(n_266), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_266), .B(n_315), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_267), .B(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g358 ( .A(n_267), .B(n_304), .Y(n_358) );
INVx3_ASAP7_75t_SL g399 ( .A(n_267), .Y(n_399) );
AND2x2_ASAP7_75t_L g343 ( .A(n_268), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g372 ( .A(n_268), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_268), .B(n_281), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_268), .B(n_327), .Y(n_413) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx3_ASAP7_75t_L g315 ( .A(n_269), .Y(n_315) );
OAI322xp33_ASAP7_75t_L g410 ( .A1(n_269), .A2(n_341), .A3(n_363), .B1(n_411), .B2(n_413), .C1(n_414), .C2(n_415), .Y(n_410) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AOI21xp33_ASAP7_75t_L g434 ( .A1(n_280), .A2(n_283), .B(n_435), .Y(n_434) );
NOR2xp33_ASAP7_75t_SL g360 ( .A(n_281), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g382 ( .A(n_281), .B(n_294), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_281), .B(n_321), .Y(n_397) );
INVxp67_ASAP7_75t_L g348 ( .A(n_283), .Y(n_348) );
AOI211xp5_ASAP7_75t_L g354 ( .A1(n_283), .A2(n_355), .B(n_359), .C(n_369), .Y(n_354) );
OAI221xp5_ASAP7_75t_SL g284 ( .A1(n_285), .A2(n_293), .B1(n_296), .B2(n_300), .C(n_305), .Y(n_284) );
INVxp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_291), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g308 ( .A(n_292), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g425 ( .A(n_292), .Y(n_425) );
OAI221xp5_ASAP7_75t_L g441 ( .A1(n_293), .A2(n_442), .B1(n_447), .B2(n_448), .C(n_450), .Y(n_441) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_294), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_SL g341 ( .A(n_294), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_294), .B(n_372), .Y(n_379) );
AND2x2_ASAP7_75t_L g421 ( .A(n_294), .B(n_399), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_295), .B(n_320), .Y(n_319) );
OAI22xp33_ASAP7_75t_L g416 ( .A1(n_295), .A2(n_307), .B1(n_417), .B2(n_418), .Y(n_416) );
OR2x2_ASAP7_75t_L g447 ( .A(n_295), .B(n_315), .Y(n_447) );
CKINVDCx16_ASAP7_75t_R g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g424 ( .A(n_298), .Y(n_424) );
AND2x2_ASAP7_75t_L g449 ( .A(n_298), .B(n_392), .Y(n_449) );
INVxp67_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NOR2xp33_ASAP7_75t_SL g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g313 ( .A(n_303), .B(n_314), .Y(n_313) );
AOI22xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_312), .B1(n_316), .B2(n_319), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .Y(n_307) );
INVx1_ASAP7_75t_L g380 ( .A(n_308), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_308), .B(n_348), .Y(n_415) );
AOI322xp5_ASAP7_75t_L g339 ( .A1(n_310), .A2(n_340), .A3(n_342), .B1(n_343), .B2(n_345), .C1(n_346), .C2(n_350), .Y(n_339) );
INVxp67_ASAP7_75t_L g333 ( .A(n_311), .Y(n_333) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_313), .A2(n_318), .B1(n_335), .B2(n_337), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_314), .B(n_327), .Y(n_414) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_315), .B(n_353), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_315), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g411 ( .A(n_317), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
NAND3xp33_ASAP7_75t_SL g322 ( .A(n_323), .B(n_339), .C(n_354), .Y(n_322) );
AOI221xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_325), .B1(n_330), .B2(n_332), .C(n_334), .Y(n_323) );
AND2x2_ASAP7_75t_L g330 ( .A(n_326), .B(n_331), .Y(n_330) );
INVx3_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
AND2x2_ASAP7_75t_L g340 ( .A(n_331), .B(n_341), .Y(n_340) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_333), .Y(n_412) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_338), .B(n_352), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_341), .B(n_399), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_342), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g417 ( .A(n_345), .Y(n_417) );
AND2x2_ASAP7_75t_L g432 ( .A(n_345), .B(n_409), .Y(n_432) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AOI211xp5_ASAP7_75t_L g426 ( .A1(n_356), .A2(n_427), .B(n_433), .C(n_441), .Y(n_426) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g395 ( .A(n_366), .B(n_396), .Y(n_395) );
NAND2x1_ASAP7_75t_SL g437 ( .A(n_367), .B(n_438), .Y(n_437) );
CKINVDCx16_ASAP7_75t_R g407 ( .A(n_370), .Y(n_407) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g402 ( .A(n_376), .Y(n_402) );
AND2x2_ASAP7_75t_L g406 ( .A(n_376), .B(n_392), .Y(n_406) );
NOR5xp2_ASAP7_75t_L g377 ( .A(n_378), .B(n_393), .C(n_410), .D(n_416), .E(n_419), .Y(n_377) );
OAI221xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B1(n_381), .B2(n_383), .C(n_385), .Y(n_378) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_382), .B(n_440), .Y(n_439) );
INVxp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_388), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g408 ( .A(n_392), .B(n_409), .Y(n_408) );
OAI221xp5_ASAP7_75t_SL g393 ( .A1(n_394), .A2(n_397), .B1(n_398), .B2(n_400), .C(n_403), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_406), .B1(n_407), .B2(n_408), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g446 ( .A(n_406), .Y(n_446) );
AOI211xp5_ASAP7_75t_SL g419 ( .A1(n_420), .A2(n_422), .B(n_424), .C(n_425), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVxp67_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_446), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
CKINVDCx14_ASAP7_75t_R g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g725 ( .A(n_456), .Y(n_725) );
XNOR2xp5_ASAP7_75t_L g734 ( .A(n_456), .B(n_735), .Y(n_734) );
OR2x2_ASAP7_75t_SL g456 ( .A(n_457), .B(n_678), .Y(n_456) );
NAND5xp2_ASAP7_75t_L g457 ( .A(n_458), .B(n_590), .C(n_628), .D(n_649), .E(n_666), .Y(n_457) );
NOR3xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_562), .C(n_583), .Y(n_458) );
OAI221xp5_ASAP7_75t_SL g459 ( .A1(n_460), .A2(n_502), .B1(n_525), .B2(n_549), .C(n_553), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_473), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_462), .B(n_551), .Y(n_570) );
OR2x2_ASAP7_75t_L g597 ( .A(n_462), .B(n_485), .Y(n_597) );
AND2x2_ASAP7_75t_L g611 ( .A(n_462), .B(n_485), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_462), .B(n_476), .Y(n_625) );
AND2x2_ASAP7_75t_L g663 ( .A(n_462), .B(n_627), .Y(n_663) );
AND2x2_ASAP7_75t_L g692 ( .A(n_462), .B(n_602), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_462), .B(n_574), .Y(n_709) );
INVx4_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g589 ( .A(n_463), .B(n_484), .Y(n_589) );
BUFx3_ASAP7_75t_L g614 ( .A(n_463), .Y(n_614) );
AND2x2_ASAP7_75t_L g643 ( .A(n_463), .B(n_485), .Y(n_643) );
AND3x2_ASAP7_75t_L g656 ( .A(n_463), .B(n_657), .C(n_658), .Y(n_656) );
INVx1_ASAP7_75t_L g579 ( .A(n_473), .Y(n_579) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_484), .Y(n_473) );
AOI32xp33_ASAP7_75t_L g634 ( .A1(n_474), .A2(n_586), .A3(n_635), .B1(n_638), .B2(n_639), .Y(n_634) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g561 ( .A(n_475), .B(n_484), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_475), .B(n_589), .Y(n_632) );
AND2x2_ASAP7_75t_L g639 ( .A(n_475), .B(n_611), .Y(n_639) );
OR2x2_ASAP7_75t_L g645 ( .A(n_475), .B(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_475), .B(n_600), .Y(n_670) );
OR2x2_ASAP7_75t_L g688 ( .A(n_475), .B(n_513), .Y(n_688) );
BUFx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g552 ( .A(n_476), .B(n_494), .Y(n_552) );
INVx2_ASAP7_75t_L g574 ( .A(n_476), .Y(n_574) );
OR2x2_ASAP7_75t_L g596 ( .A(n_476), .B(n_494), .Y(n_596) );
AND2x2_ASAP7_75t_L g601 ( .A(n_476), .B(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_476), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g657 ( .A(n_476), .B(n_551), .Y(n_657) );
INVx1_ASAP7_75t_SL g708 ( .A(n_484), .Y(n_708) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_494), .Y(n_484) );
INVx1_ASAP7_75t_SL g551 ( .A(n_485), .Y(n_551) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_485), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_485), .B(n_637), .Y(n_636) );
NAND3xp33_ASAP7_75t_L g703 ( .A(n_485), .B(n_574), .C(n_692), .Y(n_703) );
OA21x2_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_487), .B(n_493), .Y(n_485) );
OA21x2_ASAP7_75t_L g494 ( .A1(n_486), .A2(n_495), .B(n_501), .Y(n_494) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_486), .A2(n_505), .B(n_511), .Y(n_504) );
INVx2_ASAP7_75t_L g602 ( .A(n_494), .Y(n_602) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_494), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_512), .Y(n_502) );
INVx1_ASAP7_75t_L g638 ( .A(n_503), .Y(n_638) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g556 ( .A(n_504), .B(n_538), .Y(n_556) );
INVx2_ASAP7_75t_L g573 ( .A(n_504), .Y(n_573) );
AND2x2_ASAP7_75t_L g578 ( .A(n_504), .B(n_539), .Y(n_578) );
AND2x2_ASAP7_75t_L g593 ( .A(n_504), .B(n_526), .Y(n_593) );
AND2x2_ASAP7_75t_L g605 ( .A(n_504), .B(n_577), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_512), .B(n_621), .Y(n_620) );
NAND2x1p5_ASAP7_75t_L g677 ( .A(n_512), .B(n_578), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_512), .B(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_512), .B(n_572), .Y(n_700) );
BUFx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OR2x2_ASAP7_75t_L g537 ( .A(n_513), .B(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_513), .B(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g582 ( .A(n_513), .B(n_526), .Y(n_582) );
AND2x2_ASAP7_75t_L g608 ( .A(n_513), .B(n_538), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_513), .B(n_648), .Y(n_647) );
OA21x2_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B(n_523), .Y(n_513) );
INVx1_ASAP7_75t_L g567 ( .A(n_515), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_519), .B(n_522), .Y(n_518) );
INVx2_ASAP7_75t_L g533 ( .A(n_522), .Y(n_533) );
INVx1_ASAP7_75t_L g568 ( .A(n_523), .Y(n_568) );
OR2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_537), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_526), .B(n_559), .Y(n_558) );
AND2x4_ASAP7_75t_L g572 ( .A(n_526), .B(n_573), .Y(n_572) );
INVx3_ASAP7_75t_SL g577 ( .A(n_526), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_526), .B(n_564), .Y(n_630) );
OR2x2_ASAP7_75t_L g640 ( .A(n_526), .B(n_566), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_526), .B(n_608), .Y(n_668) );
OR2x2_ASAP7_75t_L g698 ( .A(n_526), .B(n_538), .Y(n_698) );
AND2x2_ASAP7_75t_L g702 ( .A(n_526), .B(n_539), .Y(n_702) );
NAND2xp5_ASAP7_75t_SL g715 ( .A(n_526), .B(n_578), .Y(n_715) );
AND2x2_ASAP7_75t_L g722 ( .A(n_526), .B(n_604), .Y(n_722) );
OR2x6_ASAP7_75t_L g526 ( .A(n_527), .B(n_535), .Y(n_526) );
INVx1_ASAP7_75t_SL g665 ( .A(n_537), .Y(n_665) );
AND2x2_ASAP7_75t_L g604 ( .A(n_538), .B(n_566), .Y(n_604) );
AND2x2_ASAP7_75t_L g618 ( .A(n_538), .B(n_573), .Y(n_618) );
AND2x2_ASAP7_75t_L g621 ( .A(n_538), .B(n_577), .Y(n_621) );
INVx1_ASAP7_75t_L g648 ( .A(n_538), .Y(n_648) );
INVx2_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
BUFx2_ASAP7_75t_L g560 ( .A(n_539), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
A2O1A1Ixp33_ASAP7_75t_L g719 ( .A1(n_550), .A2(n_596), .B(n_720), .C(n_721), .Y(n_719) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g626 ( .A(n_551), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_552), .B(n_569), .Y(n_584) );
AND2x2_ASAP7_75t_L g610 ( .A(n_552), .B(n_611), .Y(n_610) );
OAI21xp5_ASAP7_75t_SL g553 ( .A1(n_554), .A2(n_557), .B(n_561), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_555), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g581 ( .A(n_556), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_556), .B(n_577), .Y(n_622) );
AND2x2_ASAP7_75t_L g713 ( .A(n_556), .B(n_564), .Y(n_713) );
INVxp67_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g586 ( .A(n_560), .B(n_573), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_560), .B(n_571), .Y(n_587) );
OAI322xp33_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_570), .A3(n_571), .B1(n_574), .B2(n_575), .C1(n_579), .C2(n_580), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_569), .Y(n_563) );
AND2x2_ASAP7_75t_L g674 ( .A(n_564), .B(n_586), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_564), .B(n_638), .Y(n_720) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g617 ( .A(n_566), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g683 ( .A(n_570), .B(n_596), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_571), .B(n_665), .Y(n_664) );
INVx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_572), .B(n_604), .Y(n_661) );
AND2x2_ASAP7_75t_L g607 ( .A(n_573), .B(n_577), .Y(n_607) );
AND2x2_ASAP7_75t_L g615 ( .A(n_574), .B(n_616), .Y(n_615) );
A2O1A1Ixp33_ASAP7_75t_L g712 ( .A1(n_574), .A2(n_653), .B(n_713), .C(n_714), .Y(n_712) );
AOI21xp33_ASAP7_75t_L g685 ( .A1(n_575), .A2(n_588), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_577), .B(n_604), .Y(n_644) );
AND2x2_ASAP7_75t_L g650 ( .A(n_577), .B(n_618), .Y(n_650) );
AND2x2_ASAP7_75t_L g684 ( .A(n_577), .B(n_586), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_578), .B(n_593), .Y(n_592) );
INVx2_ASAP7_75t_SL g694 ( .A(n_578), .Y(n_694) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_582), .A2(n_610), .B1(n_612), .B2(n_617), .Y(n_609) );
OAI22xp5_ASAP7_75t_SL g583 ( .A1(n_584), .A2(n_585), .B1(n_587), .B2(n_588), .Y(n_583) );
OAI22xp33_ASAP7_75t_L g619 ( .A1(n_584), .A2(n_620), .B1(n_622), .B2(n_623), .Y(n_619) );
INVxp67_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_589), .A2(n_691), .B1(n_693), .B2(n_695), .C(n_699), .Y(n_690) );
AOI211xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_594), .B(n_598), .C(n_619), .Y(n_590) );
INVxp67_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
OR2x2_ASAP7_75t_L g660 ( .A(n_596), .B(n_613), .Y(n_660) );
INVx1_ASAP7_75t_L g711 ( .A(n_596), .Y(n_711) );
OAI221xp5_ASAP7_75t_L g598 ( .A1(n_597), .A2(n_599), .B1(n_603), .B2(n_606), .C(n_609), .Y(n_598) );
INVx2_ASAP7_75t_SL g653 ( .A(n_597), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g718 ( .A(n_600), .Y(n_718) );
AND2x2_ASAP7_75t_L g642 ( .A(n_601), .B(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g627 ( .A(n_602), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVx1_ASAP7_75t_L g689 ( .A(n_605), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_613), .B(n_715), .Y(n_714) );
CKINVDCx16_ASAP7_75t_R g613 ( .A(n_614), .Y(n_613) );
INVxp67_ASAP7_75t_L g658 ( .A(n_616), .Y(n_658) );
O2A1O1Ixp33_ASAP7_75t_L g628 ( .A1(n_617), .A2(n_629), .B(n_631), .C(n_633), .Y(n_628) );
INVx1_ASAP7_75t_L g706 ( .A(n_620), .Y(n_706) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_624), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
INVx2_ASAP7_75t_L g637 ( .A(n_627), .Y(n_637) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OAI222xp33_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_640), .B1(n_641), .B2(n_644), .C1(n_645), .C2(n_647), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_SL g673 ( .A(n_637), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_640), .B(n_694), .Y(n_693) );
NAND2xp33_ASAP7_75t_SL g671 ( .A(n_641), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_SL g646 ( .A(n_643), .Y(n_646) );
AND2x2_ASAP7_75t_L g710 ( .A(n_643), .B(n_711), .Y(n_710) );
OR2x2_ASAP7_75t_L g676 ( .A(n_646), .B(n_673), .Y(n_676) );
INVx1_ASAP7_75t_L g705 ( .A(n_647), .Y(n_705) );
AOI211xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_651), .B(n_654), .C(n_659), .Y(n_649) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_653), .B(n_673), .Y(n_672) );
INVx2_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
AOI322xp5_ASAP7_75t_L g704 ( .A1(n_656), .A2(n_684), .A3(n_689), .B1(n_705), .B2(n_706), .C1(n_707), .C2(n_710), .Y(n_704) );
AND2x2_ASAP7_75t_L g691 ( .A(n_657), .B(n_692), .Y(n_691) );
OAI22xp33_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_661), .B1(n_662), .B2(n_664), .Y(n_659) );
INVxp33_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AOI221xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_669), .B1(n_671), .B2(n_674), .C(n_675), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
NAND5xp2_ASAP7_75t_L g678 ( .A(n_679), .B(n_690), .C(n_704), .D(n_712), .E(n_716), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_684), .B(n_685), .Y(n_679) );
INVxp67_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVxp33_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
A2O1A1Ixp33_ASAP7_75t_L g716 ( .A1(n_692), .A2(n_717), .B(n_718), .C(n_719), .Y(n_716) );
AOI31xp33_ASAP7_75t_L g699 ( .A1(n_694), .A2(n_700), .A3(n_701), .B(n_703), .Y(n_699) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
INVx1_ASAP7_75t_L g717 ( .A(n_715), .Y(n_717) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g727 ( .A(n_723), .Y(n_727) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_737), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_743), .Y(n_742) );
endmodule