module fake_jpeg_16126_n_33 (n_3, n_2, n_1, n_0, n_4, n_5, n_33);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_33;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx6_ASAP7_75t_SL g6 ( 
.A(n_2),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_4),
.B(n_5),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_SL g8 ( 
.A(n_5),
.B(n_3),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_4),
.B(n_3),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_8),
.B(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_6),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_15)
);

OAI32xp33_ASAP7_75t_L g19 ( 
.A1(n_15),
.A2(n_16),
.A3(n_17),
.B1(n_7),
.B2(n_11),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_0),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_6),
.A2(n_1),
.B1(n_2),
.B2(n_11),
.Y(n_17)
);

OAI21xp33_ASAP7_75t_SL g23 ( 
.A1(n_19),
.A2(n_17),
.B(n_16),
.Y(n_23)
);

AND2x6_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_1),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_13),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_25),
.B(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_24),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_18),
.A2(n_11),
.B1(n_7),
.B2(n_10),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_11),
.C(n_10),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_29),
.C(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_27),
.B(n_24),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_31),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_22),
.Y(n_33)
);


endmodule