module real_jpeg_22998_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_35;
wire n_33;
wire n_38;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_23;
wire n_11;
wire n_14;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_40;
wire n_36;
wire n_39;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_2),
.A2(n_19),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

AO21x1_ASAP7_75t_SL g41 ( 
.A1(n_2),
.A2(n_17),
.B(n_20),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_3),
.B(n_11),
.Y(n_35)
);

OR2x2_ASAP7_75t_SL g39 ( 
.A(n_3),
.B(n_11),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_4),
.B(n_15),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_4),
.B(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_5),
.B(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_5),
.B(n_18),
.Y(n_20)
);

NOR3xp33_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_33),
.C(n_40),
.Y(n_6)
);

OAI22xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_12),
.B1(n_28),
.B2(n_29),
.Y(n_7)
);

INVx1_ASAP7_75t_SL g8 ( 
.A(n_9),
.Y(n_8)
);

AND2x2_ASAP7_75t_SL g9 ( 
.A(n_10),
.B(n_11),
.Y(n_9)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_11),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_21),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_23),
.Y(n_32)
);

OA21x2_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_19),
.B(n_20),
.Y(n_16)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_27),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_20),
.Y(n_27)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_24),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_23),
.B(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_23),
.B(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_24),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);


endmodule