module fake_jpeg_24728_n_179 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_14),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_16),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_38),
.Y(n_45)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_43),
.Y(n_46)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_41),
.Y(n_61)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_1),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_23),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_28),
.B1(n_18),
.B2(n_20),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_41),
.B1(n_24),
.B2(n_23),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_20),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_54),
.Y(n_70)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_59),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_32),
.B1(n_40),
.B2(n_37),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_58),
.A2(n_22),
.B1(n_18),
.B2(n_21),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_26),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_43),
.B1(n_35),
.B2(n_22),
.Y(n_62)
);

AO22x1_ASAP7_75t_SL g102 ( 
.A1(n_62),
.A2(n_73),
.B1(n_42),
.B2(n_31),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_54),
.A2(n_20),
.B1(n_18),
.B2(n_32),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_72),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_66),
.B(n_67),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_45),
.B(n_39),
.Y(n_68)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_71),
.A2(n_21),
.B(n_30),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_41),
.B1(n_22),
.B2(n_42),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_22),
.B1(n_15),
.B2(n_24),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_76),
.Y(n_92)
);

BUFx4f_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_80),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_16),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_79),
.B(n_83),
.Y(n_90)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_47),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_17),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_17),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_86),
.B(n_26),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_42),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_95),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_94),
.B(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_67),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_79),
.B(n_25),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_99),
.A2(n_102),
.B1(n_80),
.B2(n_75),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g100 ( 
.A1(n_67),
.A2(n_2),
.B(n_3),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_106),
.B(n_29),
.C(n_72),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_71),
.B(n_30),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_105),
.B(n_13),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_73),
.A2(n_29),
.B(n_25),
.Y(n_106)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_115),
.Y(n_126)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_109),
.Y(n_127)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_77),
.Y(n_110)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_63),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_111),
.B(n_114),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_121),
.B1(n_96),
.B2(n_84),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_78),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_73),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_102),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_123),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_119),
.A2(n_95),
.B(n_90),
.Y(n_132)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_122),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_73),
.B1(n_84),
.B2(n_75),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_104),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_91),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_132),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_101),
.Y(n_129)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_134),
.B(n_135),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_108),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_96),
.B(n_106),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_137),
.A2(n_119),
.B(n_115),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_101),
.C(n_105),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_120),
.C(n_90),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_85),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_117),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_141),
.B(n_143),
.C(n_147),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_145),
.A2(n_146),
.B(n_149),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_137),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_118),
.C(n_121),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_113),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_150),
.B(n_138),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_141),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_153),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_155),
.Y(n_159)
);

A2O1A1O1Ixp25_ASAP7_75t_L g153 ( 
.A1(n_146),
.A2(n_130),
.B(n_132),
.C(n_126),
.D(n_131),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_127),
.C(n_136),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_69),
.Y(n_156)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_156),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_148),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_158),
.B(n_98),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_157),
.A2(n_147),
.B1(n_144),
.B2(n_142),
.Y(n_161)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_161),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_69),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_154),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_153),
.C(n_69),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_151),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_165),
.B(n_168),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_167),
.A2(n_169),
.B1(n_159),
.B2(n_2),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_91),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_166),
.A2(n_164),
.B1(n_162),
.B2(n_104),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_171),
.A2(n_173),
.B(n_7),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_8),
.C(n_9),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_L g173 ( 
.A1(n_167),
.A2(n_6),
.B(n_7),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_174),
.B(n_175),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_176),
.B(n_170),
.Y(n_177)
);

AO21x1_ASAP7_75t_L g178 ( 
.A1(n_177),
.A2(n_172),
.B(n_14),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_2),
.Y(n_179)
);


endmodule