module fake_netlist_1_3508_n_529 (n_117, n_44, n_133, n_149, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_125, n_9, n_161, n_10, n_130, n_103, n_19, n_87, n_137, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_165, n_146, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_46, n_31, n_58, n_122, n_138, n_126, n_118, n_32, n_0, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_162, n_75, n_163, n_105, n_159, n_72, n_136, n_43, n_76, n_89, n_68, n_144, n_27, n_53, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_15, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_529);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_125;
input n_9;
input n_161;
input n_10;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_165;
input n_146;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_118;
input n_32;
input n_0;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_162;
input n_75;
input n_163;
input n_105;
input n_159;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_68;
input n_144;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_15;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_529;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_431;
wire n_484;
wire n_496;
wire n_177;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_202;
wire n_386;
wire n_432;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_205;
wire n_330;
wire n_387;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_517;
wire n_479;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_259;
wire n_308;
wire n_412;
wire n_207;
wire n_224;
wire n_219;
wire n_475;
wire n_214;
wire n_204;
wire n_430;
wire n_450;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_379;
wire n_527;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_217;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_260;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_178;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_524;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_335;
wire n_272;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_198;
wire n_169;
wire n_424;
wire n_297;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_187;
wire n_375;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_421;
wire n_175;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_153), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_101), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_141), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_138), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_48), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_76), .Y(n_171) );
BUFx3_ASAP7_75t_L g172 ( .A(n_20), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_6), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_0), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_115), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_49), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_67), .Y(n_177) );
BUFx10_ASAP7_75t_L g178 ( .A(n_71), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_126), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_152), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_13), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_64), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_129), .Y(n_183) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_140), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_95), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_62), .Y(n_186) );
INVx1_ASAP7_75t_SL g187 ( .A(n_40), .Y(n_187) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_142), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_100), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_41), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_25), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_103), .Y(n_192) );
BUFx3_ASAP7_75t_L g193 ( .A(n_92), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_79), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_119), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_135), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_117), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_57), .Y(n_198) );
CKINVDCx16_ASAP7_75t_R g199 ( .A(n_50), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_31), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_131), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_125), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_91), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_56), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_111), .Y(n_205) );
OR2x2_ASAP7_75t_L g206 ( .A(n_38), .B(n_61), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_63), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_134), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_99), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_108), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_123), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_4), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_53), .Y(n_213) );
INVx2_ASAP7_75t_SL g214 ( .A(n_106), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_74), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_151), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_116), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_154), .Y(n_218) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_14), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_148), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_77), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_35), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_65), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_69), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_124), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_113), .Y(n_226) );
INVx1_ASAP7_75t_SL g227 ( .A(n_96), .Y(n_227) );
CKINVDCx16_ASAP7_75t_R g228 ( .A(n_144), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_16), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_145), .Y(n_230) );
BUFx3_ASAP7_75t_L g231 ( .A(n_155), .Y(n_231) );
INVx2_ASAP7_75t_SL g232 ( .A(n_30), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_83), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_143), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_137), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_84), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_80), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_133), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_122), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_27), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_36), .Y(n_241) );
BUFx2_ASAP7_75t_L g242 ( .A(n_120), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_118), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_156), .Y(n_244) );
BUFx3_ASAP7_75t_L g245 ( .A(n_146), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_105), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_128), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_121), .Y(n_248) );
INVx2_ASAP7_75t_SL g249 ( .A(n_158), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_44), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g251 ( .A(n_130), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g252 ( .A(n_110), .Y(n_252) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_139), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_9), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_164), .Y(n_255) );
BUFx2_ASAP7_75t_L g256 ( .A(n_132), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_160), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_149), .Y(n_258) );
INVx1_ASAP7_75t_SL g259 ( .A(n_85), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g260 ( .A(n_58), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_136), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_15), .Y(n_262) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_127), .Y(n_263) );
BUFx10_ASAP7_75t_L g264 ( .A(n_55), .Y(n_264) );
BUFx2_ASAP7_75t_L g265 ( .A(n_159), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_2), .Y(n_266) );
CKINVDCx14_ASAP7_75t_R g267 ( .A(n_68), .Y(n_267) );
NOR2xp67_ASAP7_75t_L g268 ( .A(n_161), .B(n_73), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_24), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_5), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_214), .Y(n_271) );
OAI21x1_ASAP7_75t_L g272 ( .A1(n_168), .A2(n_90), .B(n_163), .Y(n_272) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_170), .A2(n_89), .B(n_162), .Y(n_273) );
BUFx12f_ASAP7_75t_L g274 ( .A(n_178), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_253), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_242), .B(n_0), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_182), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_256), .B(n_1), .Y(n_278) );
OA21x2_ASAP7_75t_L g279 ( .A1(n_167), .A2(n_93), .B(n_157), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_176), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_181), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_265), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_232), .B(n_1), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_249), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_173), .B(n_2), .Y(n_285) );
NAND2xp33_ASAP7_75t_L g286 ( .A(n_206), .B(n_11), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_183), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_211), .Y(n_288) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_184), .Y(n_289) );
BUFx3_ASAP7_75t_L g290 ( .A(n_172), .Y(n_290) );
BUFx3_ASAP7_75t_L g291 ( .A(n_193), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_174), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_254), .B(n_3), .Y(n_293) );
INVx1_ASAP7_75t_SL g294 ( .A(n_280), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_271), .B(n_238), .Y(n_295) );
INVxp67_ASAP7_75t_SL g296 ( .A(n_292), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_293), .Y(n_297) );
INVx2_ASAP7_75t_SL g298 ( .A(n_274), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_290), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_275), .B(n_270), .Y(n_300) );
INVx2_ASAP7_75t_SL g301 ( .A(n_290), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_289), .Y(n_302) );
NAND3xp33_ASAP7_75t_L g303 ( .A(n_278), .B(n_266), .C(n_212), .Y(n_303) );
INVx2_ASAP7_75t_SL g304 ( .A(n_291), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_291), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_284), .B(n_246), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_277), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_286), .A2(n_177), .B1(n_180), .B2(n_171), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_296), .B(n_276), .Y(n_309) );
INVxp67_ASAP7_75t_SL g310 ( .A(n_296), .Y(n_310) );
INVx8_ASAP7_75t_L g311 ( .A(n_298), .Y(n_311) );
INVx4_ASAP7_75t_L g312 ( .A(n_299), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_305), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_297), .B(n_282), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_308), .B(n_199), .Y(n_315) );
NAND2xp5_ASAP7_75t_SL g316 ( .A(n_308), .B(n_228), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_307), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_301), .Y(n_318) );
INVxp67_ASAP7_75t_SL g319 ( .A(n_295), .Y(n_319) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_303), .B(n_278), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_294), .B(n_281), .Y(n_321) );
AO22x1_ASAP7_75t_L g322 ( .A1(n_295), .A2(n_285), .B1(n_283), .B2(n_169), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_319), .B(n_304), .Y(n_323) );
OAI21xp5_ASAP7_75t_L g324 ( .A1(n_320), .A2(n_273), .B(n_272), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_309), .A2(n_286), .B(n_279), .Y(n_325) );
A2O1A1Ixp33_ASAP7_75t_L g326 ( .A1(n_314), .A2(n_283), .B(n_300), .C(n_306), .Y(n_326) );
O2A1O1Ixp33_ASAP7_75t_L g327 ( .A1(n_315), .A2(n_285), .B(n_306), .C(n_288), .Y(n_327) );
BUFx2_ASAP7_75t_L g328 ( .A(n_311), .Y(n_328) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_311), .Y(n_329) );
O2A1O1Ixp5_ASAP7_75t_L g330 ( .A1(n_322), .A2(n_277), .B(n_248), .C(n_287), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_310), .A2(n_279), .B(n_189), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_316), .B(n_188), .Y(n_332) );
OAI321xp33_ASAP7_75t_L g333 ( .A1(n_321), .A2(n_224), .A3(n_194), .B1(n_195), .B2(n_186), .C(n_190), .Y(n_333) );
NAND2xp5_ASAP7_75t_SL g334 ( .A(n_318), .B(n_166), .Y(n_334) );
AO32x2_ASAP7_75t_L g335 ( .A1(n_312), .A2(n_279), .A3(n_268), .B1(n_289), .B2(n_263), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_312), .B(n_191), .Y(n_336) );
NAND2x1p5_ASAP7_75t_L g337 ( .A(n_317), .B(n_187), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_328), .Y(n_338) );
AOI21xp5_ASAP7_75t_L g339 ( .A1(n_325), .A2(n_313), .B(n_196), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_323), .Y(n_340) );
AO31x2_ASAP7_75t_L g341 ( .A1(n_331), .A2(n_192), .A3(n_200), .B(n_197), .Y(n_341) );
AOI21xp5_ASAP7_75t_L g342 ( .A1(n_324), .A2(n_205), .B(n_204), .Y(n_342) );
BUFx2_ASAP7_75t_R g343 ( .A(n_336), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_326), .B(n_233), .Y(n_344) );
A2O1A1Ixp33_ASAP7_75t_L g345 ( .A1(n_327), .A2(n_244), .B(n_221), .C(n_222), .Y(n_345) );
AOI221xp5_ASAP7_75t_SL g346 ( .A1(n_332), .A2(n_239), .B1(n_208), .B2(n_209), .C(n_210), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_323), .Y(n_347) );
OAI21x1_ASAP7_75t_L g348 ( .A1(n_330), .A2(n_213), .B(n_207), .Y(n_348) );
BUFx4_ASAP7_75t_SL g349 ( .A(n_329), .Y(n_349) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_334), .A2(n_216), .B(n_215), .Y(n_350) );
AOI21xp5_ASAP7_75t_L g351 ( .A1(n_333), .A2(n_218), .B(n_217), .Y(n_351) );
OAI21x1_ASAP7_75t_L g352 ( .A1(n_337), .A2(n_223), .B(n_220), .Y(n_352) );
OAI21xp5_ASAP7_75t_L g353 ( .A1(n_335), .A2(n_226), .B(n_225), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_335), .Y(n_354) );
AOI21xp5_ASAP7_75t_L g355 ( .A1(n_325), .A2(n_235), .B(n_230), .Y(n_355) );
OA21x2_ASAP7_75t_L g356 ( .A1(n_331), .A2(n_240), .B(n_237), .Y(n_356) );
OAI21x1_ASAP7_75t_SL g357 ( .A1(n_353), .A2(n_354), .B(n_355), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_344), .A2(n_178), .B1(n_264), .B2(n_251), .Y(n_358) );
OAI21x1_ASAP7_75t_L g359 ( .A1(n_339), .A2(n_243), .B(n_241), .Y(n_359) );
AND2x4_ASAP7_75t_L g360 ( .A(n_340), .B(n_252), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_347), .Y(n_361) );
INVx6_ASAP7_75t_L g362 ( .A(n_349), .Y(n_362) );
BUFx2_ASAP7_75t_SL g363 ( .A(n_338), .Y(n_363) );
AO21x2_ASAP7_75t_L g364 ( .A1(n_342), .A2(n_250), .B(n_247), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_343), .B(n_260), .Y(n_365) );
OAI21x1_ASAP7_75t_L g366 ( .A1(n_348), .A2(n_258), .B(n_255), .Y(n_366) );
OA21x2_ASAP7_75t_L g367 ( .A1(n_346), .A2(n_262), .B(n_261), .Y(n_367) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_352), .Y(n_368) );
OA21x2_ASAP7_75t_L g369 ( .A1(n_345), .A2(n_302), .B(n_227), .Y(n_369) );
AO21x2_ASAP7_75t_L g370 ( .A1(n_351), .A2(n_302), .B(n_289), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_341), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_350), .B(n_267), .Y(n_372) );
AO31x2_ASAP7_75t_L g373 ( .A1(n_356), .A2(n_289), .A3(n_184), .B(n_263), .Y(n_373) );
AOI22x1_ASAP7_75t_L g374 ( .A1(n_341), .A2(n_227), .B1(n_187), .B2(n_259), .Y(n_374) );
O2A1O1Ixp33_ASAP7_75t_L g375 ( .A1(n_356), .A2(n_259), .B(n_245), .C(n_231), .Y(n_375) );
OA21x2_ASAP7_75t_L g376 ( .A1(n_354), .A2(n_179), .B(n_175), .Y(n_376) );
OA21x2_ASAP7_75t_L g377 ( .A1(n_354), .A2(n_198), .B(n_185), .Y(n_377) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_349), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_344), .B(n_264), .Y(n_379) );
AO21x2_ASAP7_75t_L g380 ( .A1(n_353), .A2(n_263), .B(n_184), .Y(n_380) );
AOI21x1_ASAP7_75t_L g381 ( .A1(n_354), .A2(n_17), .B(n_12), .Y(n_381) );
INVx6_ASAP7_75t_L g382 ( .A(n_349), .Y(n_382) );
AO31x2_ASAP7_75t_L g383 ( .A1(n_354), .A2(n_3), .A3(n_4), .B(n_5), .Y(n_383) );
OR2x6_ASAP7_75t_L g384 ( .A(n_349), .B(n_6), .Y(n_384) );
OA21x2_ASAP7_75t_L g385 ( .A1(n_354), .A2(n_269), .B(n_257), .Y(n_385) );
OAI21x1_ASAP7_75t_L g386 ( .A1(n_339), .A2(n_107), .B(n_165), .Y(n_386) );
OA21x2_ASAP7_75t_L g387 ( .A1(n_354), .A2(n_236), .B(n_234), .Y(n_387) );
OA21x2_ASAP7_75t_L g388 ( .A1(n_354), .A2(n_229), .B(n_219), .Y(n_388) );
OAI21x1_ASAP7_75t_L g389 ( .A1(n_339), .A2(n_104), .B(n_150), .Y(n_389) );
OAI21x1_ASAP7_75t_L g390 ( .A1(n_339), .A2(n_102), .B(n_147), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_361), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_360), .B(n_7), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_360), .B(n_8), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_368), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_383), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_379), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_367), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_363), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_374), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_384), .A2(n_382), .B1(n_362), .B2(n_364), .Y(n_400) );
AO21x2_ASAP7_75t_L g401 ( .A1(n_357), .A2(n_9), .B(n_10), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_369), .B(n_201), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_378), .B(n_202), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_359), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_366), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_365), .B(n_358), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_372), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_369), .B(n_203), .Y(n_408) );
NAND2x1p5_ASAP7_75t_L g409 ( .A(n_386), .B(n_18), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_373), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_381), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_376), .B(n_19), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_380), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_389), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_390), .Y(n_415) );
OAI21xp5_ASAP7_75t_L g416 ( .A1(n_375), .A2(n_21), .B(n_22), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_377), .Y(n_417) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_377), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_385), .B(n_23), .Y(n_419) );
OAI21x1_ASAP7_75t_L g420 ( .A1(n_385), .A2(n_26), .B(n_28), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_387), .A2(n_29), .B1(n_32), .B2(n_33), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_387), .B(n_34), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_388), .Y(n_423) );
OAI21x1_ASAP7_75t_L g424 ( .A1(n_370), .A2(n_37), .B(n_39), .Y(n_424) );
OR2x6_ASAP7_75t_L g425 ( .A(n_362), .B(n_42), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_371), .B(n_43), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_361), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_360), .B(n_45), .Y(n_428) );
BUFx4f_ASAP7_75t_SL g429 ( .A(n_362), .Y(n_429) );
OAI22xp33_ASAP7_75t_L g430 ( .A1(n_384), .A2(n_46), .B1(n_47), .B2(n_51), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_373), .Y(n_431) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_394), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_396), .B(n_52), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_392), .B(n_393), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_394), .Y(n_435) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_398), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_427), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_391), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_428), .B(n_54), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_407), .B(n_59), .Y(n_440) );
AND2x4_ASAP7_75t_SL g441 ( .A(n_425), .B(n_60), .Y(n_441) );
BUFx3_ASAP7_75t_L g442 ( .A(n_429), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_395), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_400), .B(n_66), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_401), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_397), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_406), .B(n_70), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_403), .B(n_72), .Y(n_448) );
NAND3xp33_ASAP7_75t_L g449 ( .A(n_399), .B(n_75), .C(n_78), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_426), .Y(n_450) );
BUFx2_ASAP7_75t_L g451 ( .A(n_429), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_405), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_426), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_404), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_402), .B(n_81), .Y(n_455) );
INVxp67_ASAP7_75t_SL g456 ( .A(n_418), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_402), .B(n_82), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_417), .Y(n_458) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_431), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_408), .Y(n_460) );
AND2x4_ASAP7_75t_L g461 ( .A(n_423), .B(n_86), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_408), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_412), .B(n_87), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_430), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_419), .B(n_88), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_434), .B(n_415), .Y(n_466) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_432), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_438), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_437), .B(n_431), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_460), .B(n_410), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_432), .B(n_430), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_435), .B(n_413), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_436), .B(n_416), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_462), .B(n_411), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_436), .B(n_422), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_458), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_436), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_443), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_464), .B(n_414), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_446), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_454), .Y(n_481) );
BUFx3_ASAP7_75t_L g482 ( .A(n_451), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_447), .B(n_409), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_461), .B(n_421), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_456), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_450), .B(n_409), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_441), .B(n_420), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_453), .B(n_424), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_481), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_466), .B(n_445), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_468), .B(n_444), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_485), .Y(n_492) );
AND2x4_ASAP7_75t_L g493 ( .A(n_472), .B(n_459), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_467), .B(n_452), .Y(n_494) );
INVxp67_ASAP7_75t_L g495 ( .A(n_482), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_481), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_478), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_476), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_498), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_498), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_489), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_490), .B(n_480), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_495), .B(n_482), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_493), .B(n_477), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_493), .B(n_475), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_497), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_499), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_503), .A2(n_471), .B1(n_484), .B2(n_483), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_500), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_502), .B(n_492), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_505), .B(n_496), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_506), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_508), .A2(n_504), .B1(n_491), .B2(n_487), .Y(n_513) );
OAI21xp33_ASAP7_75t_SL g514 ( .A1(n_511), .A2(n_484), .B(n_501), .Y(n_514) );
AOI221xp5_ASAP7_75t_L g515 ( .A1(n_514), .A2(n_512), .B1(n_509), .B2(n_507), .C(n_510), .Y(n_515) );
NAND4xp25_ASAP7_75t_L g516 ( .A(n_513), .B(n_442), .C(n_448), .D(n_487), .Y(n_516) );
OAI221xp5_ASAP7_75t_L g517 ( .A1(n_515), .A2(n_501), .B1(n_486), .B2(n_470), .C(n_457), .Y(n_517) );
NOR4xp25_ASAP7_75t_L g518 ( .A(n_516), .B(n_433), .C(n_440), .D(n_457), .Y(n_518) );
CKINVDCx12_ASAP7_75t_R g519 ( .A(n_518), .Y(n_519) );
NOR3xp33_ASAP7_75t_L g520 ( .A(n_517), .B(n_455), .C(n_449), .Y(n_520) );
OAI221xp5_ASAP7_75t_SL g521 ( .A1(n_519), .A2(n_439), .B1(n_473), .B2(n_494), .C(n_474), .Y(n_521) );
INVx2_ASAP7_75t_SL g522 ( .A(n_521), .Y(n_522) );
AOI211xp5_ASAP7_75t_L g523 ( .A1(n_522), .A2(n_520), .B(n_463), .C(n_465), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_523), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_524), .A2(n_488), .B1(n_469), .B2(n_479), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_525), .B(n_94), .Y(n_526) );
AOI21xp33_ASAP7_75t_L g527 ( .A1(n_526), .A2(n_97), .B(n_98), .Y(n_527) );
INVxp67_ASAP7_75t_L g528 ( .A(n_527), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_528), .A2(n_109), .B1(n_112), .B2(n_114), .Y(n_529) );
endmodule