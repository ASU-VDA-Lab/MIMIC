module real_aes_7106_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_119;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_756;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_728;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g488 ( .A1(n_0), .A2(n_170), .B(n_489), .C(n_492), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_1), .B(n_483), .Y(n_494) );
INVx1_ASAP7_75t_L g440 ( .A(n_2), .Y(n_440) );
NAND3xp33_ASAP7_75t_SL g767 ( .A(n_2), .B(n_748), .C(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g219 ( .A(n_3), .Y(n_219) );
OAI211xp5_ASAP7_75t_L g111 ( .A1(n_4), .A2(n_112), .B(n_442), .C(n_445), .Y(n_111) );
OAI211xp5_ASAP7_75t_L g442 ( .A1(n_4), .A2(n_114), .B(n_433), .C(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_5), .B(n_158), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_6), .A2(n_467), .B(n_537), .Y(n_536) );
OAI22xp5_ASAP7_75t_SL g429 ( .A1(n_7), .A2(n_11), .B1(n_430), .B2(n_431), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_7), .Y(n_430) );
AO21x2_ASAP7_75t_L g545 ( .A1(n_8), .A2(n_175), .B(n_546), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g169 ( .A1(n_9), .A2(n_39), .B1(n_131), .B2(n_143), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_10), .B(n_175), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_11), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_11), .A2(n_116), .B1(n_431), .B2(n_432), .Y(n_450) );
AND2x6_ASAP7_75t_L g146 ( .A(n_12), .B(n_147), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g558 ( .A1(n_13), .A2(n_146), .B(n_470), .C(n_559), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_14), .B(n_40), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_14), .B(n_40), .Y(n_766) );
INVx1_ASAP7_75t_L g127 ( .A(n_15), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_16), .B(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g213 ( .A(n_17), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_18), .B(n_158), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_19), .B(n_173), .Y(n_191) );
AO32x2_ASAP7_75t_L g167 ( .A1(n_20), .A2(n_168), .A3(n_172), .B1(n_174), .B2(n_175), .Y(n_167) );
OAI22xp5_ASAP7_75t_L g753 ( .A1(n_21), .A2(n_58), .B1(n_754), .B2(n_755), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_21), .Y(n_755) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_22), .B(n_131), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_23), .B(n_173), .Y(n_221) );
AOI22xp33_ASAP7_75t_L g171 ( .A1(n_24), .A2(n_56), .B1(n_131), .B2(n_143), .Y(n_171) );
AOI22xp33_ASAP7_75t_SL g184 ( .A1(n_25), .A2(n_83), .B1(n_131), .B2(n_135), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_26), .B(n_131), .Y(n_161) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_27), .A2(n_174), .B(n_470), .C(n_472), .Y(n_469) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_28), .A2(n_174), .B(n_470), .C(n_549), .Y(n_548) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_29), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_30), .B(n_123), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_31), .A2(n_105), .B1(n_763), .B2(n_771), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_32), .A2(n_467), .B(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_33), .B(n_123), .Y(n_165) );
INVx2_ASAP7_75t_L g133 ( .A(n_34), .Y(n_133) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_35), .A2(n_501), .B(n_502), .C(n_506), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_36), .B(n_131), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_37), .B(n_123), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_38), .B(n_138), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_41), .B(n_466), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g563 ( .A(n_42), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_43), .B(n_158), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_44), .B(n_467), .Y(n_547) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_45), .A2(n_501), .B(n_506), .C(n_528), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_46), .A2(n_751), .B1(n_752), .B2(n_753), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_46), .Y(n_751) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_47), .B(n_131), .Y(n_201) );
INVx1_ASAP7_75t_L g490 ( .A(n_48), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g182 ( .A1(n_49), .A2(n_92), .B1(n_143), .B2(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g529 ( .A(n_50), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_51), .B(n_131), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_52), .B(n_131), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_53), .B(n_436), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_54), .B(n_467), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_55), .B(n_206), .Y(n_205) );
AOI22xp33_ASAP7_75t_SL g195 ( .A1(n_57), .A2(n_62), .B1(n_131), .B2(n_135), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_58), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_59), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g130 ( .A(n_60), .B(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_61), .B(n_131), .Y(n_232) );
INVx1_ASAP7_75t_L g147 ( .A(n_63), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_64), .B(n_467), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_65), .B(n_483), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g539 ( .A1(n_66), .A2(n_206), .B(n_216), .C(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_67), .B(n_131), .Y(n_220) );
INVx1_ASAP7_75t_L g126 ( .A(n_68), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_69), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_70), .B(n_158), .Y(n_504) );
AO32x2_ASAP7_75t_L g180 ( .A1(n_71), .A2(n_174), .A3(n_175), .B1(n_181), .B2(n_185), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_72), .B(n_159), .Y(n_560) );
INVx1_ASAP7_75t_L g231 ( .A(n_73), .Y(n_231) );
INVx1_ASAP7_75t_L g156 ( .A(n_74), .Y(n_156) );
CKINVDCx16_ASAP7_75t_R g486 ( .A(n_75), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_76), .B(n_474), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_77), .B(n_115), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_77), .Y(n_434) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_78), .A2(n_470), .B(n_506), .C(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_79), .B(n_135), .Y(n_157) );
CKINVDCx16_ASAP7_75t_R g538 ( .A(n_80), .Y(n_538) );
INVx1_ASAP7_75t_L g770 ( .A(n_81), .Y(n_770) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_82), .B(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_84), .B(n_143), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_85), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_86), .B(n_135), .Y(n_162) );
AOI222xp33_ASAP7_75t_L g447 ( .A1(n_87), .A2(n_448), .B1(n_749), .B2(n_750), .C1(n_756), .C2(n_758), .Y(n_447) );
INVx2_ASAP7_75t_L g124 ( .A(n_88), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_89), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_90), .B(n_145), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_91), .B(n_135), .Y(n_202) );
OR2x2_ASAP7_75t_L g437 ( .A(n_93), .B(n_438), .Y(n_437) );
OR2x2_ASAP7_75t_L g453 ( .A(n_93), .B(n_439), .Y(n_453) );
INVx2_ASAP7_75t_L g748 ( .A(n_93), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_94), .A2(n_103), .B1(n_135), .B2(n_136), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_95), .B(n_467), .Y(n_499) );
INVx1_ASAP7_75t_L g503 ( .A(n_96), .Y(n_503) );
INVxp67_ASAP7_75t_L g541 ( .A(n_97), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_98), .B(n_135), .Y(n_229) );
INVx1_ASAP7_75t_L g516 ( .A(n_99), .Y(n_516) );
INVx1_ASAP7_75t_L g556 ( .A(n_100), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_101), .B(n_770), .Y(n_769) );
AND2x2_ASAP7_75t_L g531 ( .A(n_102), .B(n_123), .Y(n_531) );
OA21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_111), .B(n_446), .Y(n_105) );
BUFx2_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_SL g762 ( .A(n_109), .Y(n_762) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
NOR3xp33_ASAP7_75t_L g113 ( .A(n_114), .B(n_433), .C(n_436), .Y(n_113) );
INVx1_ASAP7_75t_L g435 ( .A(n_115), .Y(n_435) );
OAI22xp5_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_428), .B1(n_429), .B2(n_432), .Y(n_115) );
INVx1_ASAP7_75t_L g432 ( .A(n_116), .Y(n_432) );
OR2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_350), .Y(n_116) );
NAND5xp2_ASAP7_75t_L g117 ( .A(n_118), .B(n_269), .C(n_284), .D(n_310), .E(n_332), .Y(n_117) );
NOR2xp33_ASAP7_75t_SL g118 ( .A(n_119), .B(n_249), .Y(n_118) );
OAI221xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_186), .B1(n_222), .B2(n_238), .C(n_239), .Y(n_119) );
NOR2xp33_ASAP7_75t_SL g120 ( .A(n_121), .B(n_176), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_121), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_SL g426 ( .A(n_121), .Y(n_426) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_149), .Y(n_121) );
INVx1_ASAP7_75t_L g266 ( .A(n_122), .Y(n_266) );
AND2x2_ASAP7_75t_L g268 ( .A(n_122), .B(n_167), .Y(n_268) );
AND2x2_ASAP7_75t_L g278 ( .A(n_122), .B(n_166), .Y(n_278) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_122), .Y(n_296) );
INVx1_ASAP7_75t_L g306 ( .A(n_122), .Y(n_306) );
OR2x2_ASAP7_75t_L g344 ( .A(n_122), .B(n_243), .Y(n_344) );
INVx2_ASAP7_75t_L g394 ( .A(n_122), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_122), .B(n_242), .Y(n_411) );
OA21x2_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_128), .B(n_148), .Y(n_122) );
OA21x2_ASAP7_75t_L g152 ( .A1(n_123), .A2(n_153), .B(n_165), .Y(n_152) );
INVx2_ASAP7_75t_L g185 ( .A(n_123), .Y(n_185) );
INVx1_ASAP7_75t_L g480 ( .A(n_123), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_123), .A2(n_499), .B(n_500), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_123), .A2(n_526), .B(n_527), .Y(n_525) );
AND2x2_ASAP7_75t_SL g123 ( .A(n_124), .B(n_125), .Y(n_123) );
AND2x2_ASAP7_75t_L g173 ( .A(n_124), .B(n_125), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
OAI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_140), .B(n_146), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_134), .B(n_137), .Y(n_129) );
INVx3_ASAP7_75t_L g155 ( .A(n_131), .Y(n_155) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_131), .Y(n_518) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g143 ( .A(n_132), .Y(n_143) );
BUFx3_ASAP7_75t_L g183 ( .A(n_132), .Y(n_183) );
AND2x6_ASAP7_75t_L g470 ( .A(n_132), .B(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g136 ( .A(n_133), .Y(n_136) );
INVx1_ASAP7_75t_L g207 ( .A(n_133), .Y(n_207) );
INVx2_ASAP7_75t_L g214 ( .A(n_135), .Y(n_214) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_139), .Y(n_145) );
INVx3_ASAP7_75t_L g159 ( .A(n_139), .Y(n_159) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_139), .Y(n_164) );
AND2x2_ASAP7_75t_L g468 ( .A(n_139), .B(n_207), .Y(n_468) );
INVx1_ASAP7_75t_L g471 ( .A(n_139), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_142), .B(n_144), .Y(n_140) );
O2A1O1Ixp5_ASAP7_75t_L g230 ( .A1(n_144), .A2(n_218), .B(n_231), .C(n_232), .Y(n_230) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OAI22xp5_ASAP7_75t_L g168 ( .A1(n_145), .A2(n_169), .B1(n_170), .B2(n_171), .Y(n_168) );
OAI22xp5_ASAP7_75t_SL g181 ( .A1(n_145), .A2(n_159), .B1(n_182), .B2(n_184), .Y(n_181) );
OAI22xp5_ASAP7_75t_L g193 ( .A1(n_145), .A2(n_170), .B1(n_194), .B2(n_195), .Y(n_193) );
INVx4_ASAP7_75t_L g491 ( .A(n_145), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g153 ( .A1(n_146), .A2(n_154), .B(n_160), .Y(n_153) );
BUFx3_ASAP7_75t_L g174 ( .A(n_146), .Y(n_174) );
OAI21xp5_ASAP7_75t_L g199 ( .A1(n_146), .A2(n_200), .B(n_203), .Y(n_199) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_146), .A2(n_212), .B(n_217), .Y(n_211) );
AND2x4_ASAP7_75t_L g467 ( .A(n_146), .B(n_468), .Y(n_467) );
INVx4_ASAP7_75t_SL g493 ( .A(n_146), .Y(n_493) );
NAND2x1p5_ASAP7_75t_L g557 ( .A(n_146), .B(n_468), .Y(n_557) );
NOR2xp67_ASAP7_75t_L g149 ( .A(n_150), .B(n_166), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_151), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_151), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_SL g326 ( .A(n_151), .B(n_266), .Y(n_326) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
HB1xp67_ASAP7_75t_L g178 ( .A(n_152), .Y(n_178) );
INVx2_ASAP7_75t_L g243 ( .A(n_152), .Y(n_243) );
OR2x2_ASAP7_75t_L g305 ( .A(n_152), .B(n_306), .Y(n_305) );
O2A1O1Ixp5_ASAP7_75t_SL g154 ( .A1(n_155), .A2(n_156), .B(n_157), .C(n_158), .Y(n_154) );
INVx2_ASAP7_75t_L g170 ( .A(n_158), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_158), .A2(n_201), .B(n_202), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_158), .A2(n_228), .B(n_229), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_158), .B(n_541), .Y(n_540) );
INVx5_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_162), .B(n_163), .Y(n_160) );
INVx1_ASAP7_75t_L g216 ( .A(n_163), .Y(n_216) );
INVx4_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g474 ( .A(n_164), .Y(n_474) );
AND2x2_ASAP7_75t_L g244 ( .A(n_166), .B(n_180), .Y(n_244) );
AND2x2_ASAP7_75t_L g261 ( .A(n_166), .B(n_241), .Y(n_261) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_L g179 ( .A(n_167), .B(n_180), .Y(n_179) );
BUFx2_ASAP7_75t_L g264 ( .A(n_167), .Y(n_264) );
AND2x2_ASAP7_75t_L g393 ( .A(n_167), .B(n_394), .Y(n_393) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_170), .A2(n_204), .B(n_205), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_170), .A2(n_218), .B(n_219), .C(n_220), .Y(n_217) );
INVx2_ASAP7_75t_L g210 ( .A(n_172), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_172), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_173), .Y(n_175) );
NAND3xp33_ASAP7_75t_L g192 ( .A(n_174), .B(n_193), .C(n_196), .Y(n_192) );
OAI21xp5_ASAP7_75t_L g226 ( .A1(n_174), .A2(n_227), .B(n_230), .Y(n_226) );
INVx4_ASAP7_75t_L g196 ( .A(n_175), .Y(n_196) );
OA21x2_ASAP7_75t_L g198 ( .A1(n_175), .A2(n_199), .B(n_208), .Y(n_198) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_175), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_175), .A2(n_547), .B(n_548), .Y(n_546) );
INVx1_ASAP7_75t_L g238 ( .A(n_176), .Y(n_238) );
AND2x2_ASAP7_75t_L g176 ( .A(n_177), .B(n_179), .Y(n_176) );
AND2x2_ASAP7_75t_L g356 ( .A(n_177), .B(n_244), .Y(n_356) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g357 ( .A(n_178), .B(n_268), .Y(n_357) );
O2A1O1Ixp33_ASAP7_75t_L g324 ( .A1(n_179), .A2(n_325), .B(n_327), .C(n_329), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_179), .B(n_325), .Y(n_334) );
AOI221xp5_ASAP7_75t_L g397 ( .A1(n_179), .A2(n_255), .B1(n_398), .B2(n_399), .C(n_401), .Y(n_397) );
INVx1_ASAP7_75t_L g241 ( .A(n_180), .Y(n_241) );
INVx1_ASAP7_75t_L g277 ( .A(n_180), .Y(n_277) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_180), .Y(n_286) );
INVx2_ASAP7_75t_L g492 ( .A(n_183), .Y(n_492) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_183), .Y(n_505) );
INVx1_ASAP7_75t_L g477 ( .A(n_185), .Y(n_477) );
INVx1_ASAP7_75t_SL g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_197), .Y(n_187) );
AND2x2_ASAP7_75t_L g303 ( .A(n_188), .B(n_248), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_188), .B(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_189), .B(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g395 ( .A(n_189), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g427 ( .A(n_189), .Y(n_427) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx3_ASAP7_75t_L g257 ( .A(n_190), .Y(n_257) );
AND2x2_ASAP7_75t_L g283 ( .A(n_190), .B(n_237), .Y(n_283) );
NOR2x1_ASAP7_75t_L g292 ( .A(n_190), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g299 ( .A(n_190), .B(n_300), .Y(n_299) );
AND2x4_ASAP7_75t_L g190 ( .A(n_191), .B(n_192), .Y(n_190) );
INVx1_ASAP7_75t_L g235 ( .A(n_191), .Y(n_235) );
AO21x1_ASAP7_75t_L g234 ( .A1(n_193), .A2(n_196), .B(n_235), .Y(n_234) );
INVx3_ASAP7_75t_L g483 ( .A(n_196), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_196), .B(n_508), .Y(n_507) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_196), .A2(n_513), .B(n_520), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_196), .B(n_521), .Y(n_520) );
AO21x2_ASAP7_75t_L g554 ( .A1(n_196), .A2(n_555), .B(n_562), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_197), .B(n_339), .Y(n_374) );
INVx1_ASAP7_75t_SL g378 ( .A(n_197), .Y(n_378) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_209), .Y(n_197) );
INVx3_ASAP7_75t_L g237 ( .A(n_198), .Y(n_237) );
AND2x2_ASAP7_75t_L g248 ( .A(n_198), .B(n_225), .Y(n_248) );
AND2x2_ASAP7_75t_L g270 ( .A(n_198), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g315 ( .A(n_198), .B(n_309), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_198), .B(n_247), .Y(n_396) );
INVx2_ASAP7_75t_L g218 ( .A(n_206), .Y(n_218) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g236 ( .A(n_209), .B(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g247 ( .A(n_209), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_209), .B(n_225), .Y(n_272) );
AND2x2_ASAP7_75t_L g308 ( .A(n_209), .B(n_309), .Y(n_308) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_221), .Y(n_209) );
OA21x2_ASAP7_75t_L g225 ( .A1(n_210), .A2(n_226), .B(n_233), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_215), .C(n_216), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_214), .A2(n_550), .B(n_551), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_214), .A2(n_560), .B(n_561), .Y(n_559) );
O2A1O1Ixp33_ASAP7_75t_L g515 ( .A1(n_216), .A2(n_516), .B(n_517), .C(n_518), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_218), .A2(n_473), .B(n_475), .Y(n_472) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_236), .Y(n_223) );
INVx1_ASAP7_75t_L g288 ( .A(n_224), .Y(n_288) );
AND2x2_ASAP7_75t_L g330 ( .A(n_224), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g336 ( .A(n_224), .B(n_251), .Y(n_336) );
AOI21xp5_ASAP7_75t_SL g410 ( .A1(n_224), .A2(n_242), .B(n_265), .Y(n_410) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_234), .Y(n_224) );
OR2x2_ASAP7_75t_L g253 ( .A(n_225), .B(n_234), .Y(n_253) );
AND2x2_ASAP7_75t_L g300 ( .A(n_225), .B(n_237), .Y(n_300) );
INVx2_ASAP7_75t_L g309 ( .A(n_225), .Y(n_309) );
INVx1_ASAP7_75t_L g415 ( .A(n_225), .Y(n_415) );
AND2x2_ASAP7_75t_L g339 ( .A(n_234), .B(n_309), .Y(n_339) );
INVx1_ASAP7_75t_L g364 ( .A(n_234), .Y(n_364) );
AND2x2_ASAP7_75t_L g273 ( .A(n_236), .B(n_257), .Y(n_273) );
AND2x2_ASAP7_75t_L g285 ( .A(n_236), .B(n_286), .Y(n_285) );
INVx2_ASAP7_75t_SL g403 ( .A(n_236), .Y(n_403) );
INVx2_ASAP7_75t_L g293 ( .A(n_237), .Y(n_293) );
AND2x2_ASAP7_75t_L g331 ( .A(n_237), .B(n_247), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_237), .B(n_415), .Y(n_414) );
OAI21xp33_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_244), .B(n_245), .Y(n_239) );
AND2x2_ASAP7_75t_L g346 ( .A(n_240), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g400 ( .A(n_240), .Y(n_400) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
INVx1_ASAP7_75t_L g320 ( .A(n_241), .Y(n_320) );
BUFx2_ASAP7_75t_L g419 ( .A(n_241), .Y(n_419) );
BUFx2_ASAP7_75t_L g290 ( .A(n_242), .Y(n_290) );
AND2x2_ASAP7_75t_L g392 ( .A(n_242), .B(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g375 ( .A(n_243), .Y(n_375) );
AND2x4_ASAP7_75t_L g302 ( .A(n_244), .B(n_265), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g338 ( .A(n_244), .B(n_326), .Y(n_338) );
AOI32xp33_ASAP7_75t_L g262 ( .A1(n_245), .A2(n_263), .A3(n_265), .B1(n_267), .B2(n_268), .Y(n_262) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_248), .Y(n_245) );
INVx3_ASAP7_75t_L g251 ( .A(n_246), .Y(n_251) );
OR2x2_ASAP7_75t_L g387 ( .A(n_246), .B(n_343), .Y(n_387) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g256 ( .A(n_247), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g363 ( .A(n_247), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g255 ( .A(n_248), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g267 ( .A(n_248), .B(n_257), .Y(n_267) );
INVx1_ASAP7_75t_L g388 ( .A(n_248), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_248), .B(n_363), .Y(n_421) );
A2O1A1Ixp33_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_254), .B(n_258), .C(n_262), .Y(n_249) );
OAI322xp33_ASAP7_75t_L g358 ( .A1(n_250), .A2(n_295), .A3(n_359), .B1(n_361), .B2(n_365), .C1(n_366), .C2(n_370), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
INVxp67_ASAP7_75t_L g323 ( .A(n_251), .Y(n_323) );
INVx1_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g377 ( .A(n_253), .B(n_378), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_253), .B(n_293), .Y(n_424) );
INVxp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g316 ( .A(n_256), .Y(n_316) );
OR2x2_ASAP7_75t_L g402 ( .A(n_257), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_260), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g311 ( .A(n_261), .B(n_290), .Y(n_311) );
AND2x2_ASAP7_75t_L g382 ( .A(n_261), .B(n_295), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_261), .B(n_369), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g269 ( .A1(n_263), .A2(n_270), .B1(n_273), .B2(n_274), .C(n_279), .Y(n_269) );
OR2x2_ASAP7_75t_L g280 ( .A(n_263), .B(n_276), .Y(n_280) );
AND2x2_ASAP7_75t_L g368 ( .A(n_263), .B(n_369), .Y(n_368) );
AOI32xp33_ASAP7_75t_L g407 ( .A1(n_263), .A2(n_293), .A3(n_408), .B1(n_409), .B2(n_412), .Y(n_407) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND3xp33_ASAP7_75t_L g341 ( .A(n_264), .B(n_300), .C(n_323), .Y(n_341) );
AND2x2_ASAP7_75t_L g367 ( .A(n_264), .B(n_360), .Y(n_367) );
INVxp67_ASAP7_75t_L g347 ( .A(n_265), .Y(n_347) );
BUFx3_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g376 ( .A(n_268), .B(n_320), .Y(n_376) );
INVx2_ASAP7_75t_L g386 ( .A(n_268), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_268), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g355 ( .A(n_271), .Y(n_355) );
OR2x2_ASAP7_75t_L g281 ( .A(n_272), .B(n_282), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_274), .B(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_278), .Y(n_274) );
INVx1_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_277), .Y(n_360) );
AND2x2_ASAP7_75t_L g319 ( .A(n_278), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g365 ( .A(n_278), .Y(n_365) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_278), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
AOI21xp33_ASAP7_75t_SL g304 ( .A1(n_280), .A2(n_305), .B(n_307), .Y(n_304) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g398 ( .A(n_283), .B(n_308), .Y(n_398) );
AOI211xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_287), .B(n_297), .C(n_304), .Y(n_284) );
AND2x2_ASAP7_75t_L g328 ( .A(n_286), .B(n_296), .Y(n_328) );
INVx2_ASAP7_75t_L g343 ( .A(n_286), .Y(n_343) );
OR2x2_ASAP7_75t_L g381 ( .A(n_286), .B(n_344), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_286), .B(n_424), .Y(n_423) );
AOI211xp5_ASAP7_75t_SL g287 ( .A1(n_288), .A2(n_289), .B(n_291), .C(n_294), .Y(n_287) );
INVxp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_290), .B(n_328), .Y(n_327) );
OAI211xp5_ASAP7_75t_L g409 ( .A1(n_291), .A2(n_386), .B(n_410), .C(n_411), .Y(n_409) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2x1p5_ASAP7_75t_L g307 ( .A(n_292), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g349 ( .A(n_293), .B(n_339), .Y(n_349) );
INVx1_ASAP7_75t_L g354 ( .A(n_293), .Y(n_354) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_298), .B(n_301), .Y(n_297) );
INVxp33_ASAP7_75t_L g405 ( .A(n_299), .Y(n_405) );
AND2x2_ASAP7_75t_L g384 ( .A(n_300), .B(n_363), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g366 ( .A1(n_305), .A2(n_367), .B(n_368), .Y(n_366) );
OAI322xp33_ASAP7_75t_L g385 ( .A1(n_307), .A2(n_386), .A3(n_387), .B1(n_388), .B2(n_389), .C1(n_391), .C2(n_395), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_312), .B1(n_317), .B2(n_321), .C(n_324), .Y(n_310) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g362 ( .A(n_315), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g406 ( .A(n_319), .Y(n_406) );
INVxp67_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_322), .B(n_342), .Y(n_408) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g371 ( .A(n_331), .B(n_339), .Y(n_371) );
AOI221xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_335), .B1(n_337), .B2(n_339), .C(n_340), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AOI221xp5_ASAP7_75t_L g351 ( .A1(n_335), .A2(n_352), .B1(n_356), .B2(n_357), .C(n_358), .Y(n_351) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVxp67_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_339), .B(n_354), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_342), .B1(n_345), .B2(n_348), .Y(n_340) );
OR2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx2_ASAP7_75t_SL g369 ( .A(n_344), .Y(n_369) );
INVxp67_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND5xp2_ASAP7_75t_L g350 ( .A(n_351), .B(n_372), .C(n_397), .D(n_407), .E(n_417), .Y(n_350) );
NAND2xp5_ASAP7_75t_SL g352 ( .A(n_353), .B(n_355), .Y(n_352) );
NOR4xp25_ASAP7_75t_L g425 ( .A(n_354), .B(n_360), .C(n_426), .D(n_427), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g417 ( .A1(n_357), .A2(n_418), .B1(n_420), .B2(n_422), .C(n_425), .Y(n_417) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g416 ( .A(n_363), .Y(n_416) );
OAI322xp33_ASAP7_75t_L g373 ( .A1(n_367), .A2(n_374), .A3(n_375), .B1(n_376), .B2(n_377), .C1(n_379), .C2(n_383), .Y(n_373) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_373), .B(n_385), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g418 ( .A(n_393), .B(n_419), .Y(n_418) );
OAI22xp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_404), .B1(n_405), .B2(n_406), .Y(n_401) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_416), .Y(n_413) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVxp67_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
INVx1_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g444 ( .A(n_437), .Y(n_444) );
NOR2x2_ASAP7_75t_L g760 ( .A(n_438), .B(n_748), .Y(n_760) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OR2x2_ASAP7_75t_L g747 ( .A(n_439), .B(n_748), .Y(n_747) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NAND3xp33_ASAP7_75t_L g446 ( .A(n_445), .B(n_447), .C(n_761), .Y(n_446) );
OAI22x1_ASAP7_75t_SL g448 ( .A1(n_449), .A2(n_451), .B1(n_454), .B2(n_745), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OAI22xp5_ASAP7_75t_SL g756 ( .A1(n_450), .A2(n_455), .B1(n_745), .B2(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g757 ( .A(n_452), .Y(n_757) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_SL g455 ( .A(n_456), .B(n_700), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_635), .Y(n_456) );
NAND4xp25_ASAP7_75t_SL g457 ( .A(n_458), .B(n_580), .C(n_604), .D(n_627), .Y(n_457) );
AOI221xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_522), .B1(n_552), .B2(n_564), .C(n_567), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_495), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_461), .A2(n_481), .B1(n_523), .B2(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_461), .B(n_496), .Y(n_638) );
AND2x2_ASAP7_75t_L g657 ( .A(n_461), .B(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_461), .B(n_641), .Y(n_727) );
AND2x4_ASAP7_75t_L g461 ( .A(n_462), .B(n_481), .Y(n_461) );
AND2x2_ASAP7_75t_L g595 ( .A(n_462), .B(n_496), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_462), .B(n_610), .Y(n_609) );
OR2x2_ASAP7_75t_L g618 ( .A(n_462), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g623 ( .A(n_462), .B(n_482), .Y(n_623) );
INVx2_ASAP7_75t_L g655 ( .A(n_462), .Y(n_655) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_462), .Y(n_699) );
AND2x2_ASAP7_75t_L g716 ( .A(n_462), .B(n_593), .Y(n_716) );
INVx5_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g634 ( .A(n_463), .B(n_593), .Y(n_634) );
AND2x4_ASAP7_75t_L g648 ( .A(n_463), .B(n_481), .Y(n_648) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_463), .Y(n_652) );
AND2x2_ASAP7_75t_L g672 ( .A(n_463), .B(n_587), .Y(n_672) );
AND2x2_ASAP7_75t_L g722 ( .A(n_463), .B(n_497), .Y(n_722) );
AND2x2_ASAP7_75t_L g732 ( .A(n_463), .B(n_482), .Y(n_732) );
OR2x6_ASAP7_75t_L g463 ( .A(n_464), .B(n_478), .Y(n_463) );
AOI21xp5_ASAP7_75t_SL g464 ( .A1(n_465), .A2(n_469), .B(n_477), .Y(n_464) );
BUFx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx5_ASAP7_75t_L g487 ( .A(n_470), .Y(n_487) );
INVx2_ASAP7_75t_L g476 ( .A(n_474), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g502 ( .A1(n_476), .A2(n_503), .B(n_504), .C(n_505), .Y(n_502) );
O2A1O1Ixp33_ASAP7_75t_L g528 ( .A1(n_476), .A2(n_505), .B(n_529), .C(n_530), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
AND2x2_ASAP7_75t_L g588 ( .A(n_481), .B(n_496), .Y(n_588) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_481), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_481), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g678 ( .A(n_481), .Y(n_678) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g566 ( .A(n_482), .B(n_511), .Y(n_566) );
AND2x2_ASAP7_75t_L g593 ( .A(n_482), .B(n_512), .Y(n_593) );
OA21x2_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B(n_494), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_SL g485 ( .A1(n_486), .A2(n_487), .B(n_488), .C(n_493), .Y(n_485) );
INVx2_ASAP7_75t_L g501 ( .A(n_487), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_L g537 ( .A1(n_487), .A2(n_493), .B(n_538), .C(n_539), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
INVx1_ASAP7_75t_L g506 ( .A(n_493), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_495), .B(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_509), .Y(n_495) );
OR2x2_ASAP7_75t_L g619 ( .A(n_496), .B(n_510), .Y(n_619) );
AND2x2_ASAP7_75t_L g656 ( .A(n_496), .B(n_566), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_496), .B(n_587), .Y(n_667) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_496), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_496), .B(n_623), .Y(n_740) );
INVx5_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx2_ASAP7_75t_L g565 ( .A(n_497), .Y(n_565) );
AND2x2_ASAP7_75t_L g574 ( .A(n_497), .B(n_510), .Y(n_574) );
AND2x2_ASAP7_75t_L g690 ( .A(n_497), .B(n_585), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_497), .B(n_623), .Y(n_712) );
OR2x6_ASAP7_75t_L g497 ( .A(n_498), .B(n_507), .Y(n_497) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_510), .Y(n_658) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_511), .Y(n_610) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx2_ASAP7_75t_L g587 ( .A(n_512), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_519), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_523), .B(n_532), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_523), .B(n_600), .Y(n_719) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_524), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g571 ( .A(n_524), .B(n_572), .Y(n_571) );
INVx5_ASAP7_75t_SL g579 ( .A(n_524), .Y(n_579) );
OR2x2_ASAP7_75t_L g602 ( .A(n_524), .B(n_572), .Y(n_602) );
OR2x2_ASAP7_75t_L g612 ( .A(n_524), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g675 ( .A(n_524), .B(n_534), .Y(n_675) );
AND2x2_ASAP7_75t_SL g713 ( .A(n_524), .B(n_533), .Y(n_713) );
NOR4xp25_ASAP7_75t_L g734 ( .A(n_524), .B(n_655), .C(n_735), .D(n_736), .Y(n_734) );
AND2x2_ASAP7_75t_L g744 ( .A(n_524), .B(n_576), .Y(n_744) );
OR2x6_ASAP7_75t_L g524 ( .A(n_525), .B(n_531), .Y(n_524) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g569 ( .A(n_533), .B(n_565), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_533), .B(n_571), .Y(n_738) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_543), .Y(n_533) );
OR2x2_ASAP7_75t_L g578 ( .A(n_534), .B(n_579), .Y(n_578) );
INVx3_ASAP7_75t_L g585 ( .A(n_534), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_534), .B(n_554), .Y(n_597) );
INVxp67_ASAP7_75t_L g600 ( .A(n_534), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_534), .B(n_572), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_534), .B(n_544), .Y(n_666) );
AND2x2_ASAP7_75t_L g681 ( .A(n_534), .B(n_576), .Y(n_681) );
OR2x2_ASAP7_75t_L g710 ( .A(n_534), .B(n_544), .Y(n_710) );
OA21x2_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_536), .B(n_542), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_543), .B(n_615), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_543), .B(n_579), .Y(n_718) );
OR2x2_ASAP7_75t_L g739 ( .A(n_543), .B(n_616), .Y(n_739) );
INVx1_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
OR2x2_ASAP7_75t_L g553 ( .A(n_544), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g576 ( .A(n_544), .B(n_572), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_544), .B(n_554), .Y(n_591) );
AND2x2_ASAP7_75t_L g661 ( .A(n_544), .B(n_585), .Y(n_661) );
AND2x2_ASAP7_75t_L g695 ( .A(n_544), .B(n_579), .Y(n_695) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_545), .B(n_579), .Y(n_598) );
AND2x2_ASAP7_75t_L g626 ( .A(n_545), .B(n_554), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_552), .B(n_634), .Y(n_633) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_553), .A2(n_641), .B1(n_677), .B2(n_694), .C(n_696), .Y(n_693) );
INVx5_ASAP7_75t_SL g572 ( .A(n_554), .Y(n_572) );
OAI21xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B(n_558), .Y(n_555) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
OAI33xp33_ASAP7_75t_L g592 ( .A1(n_565), .A2(n_593), .A3(n_594), .B1(n_596), .B2(n_599), .B3(n_603), .Y(n_592) );
OR2x2_ASAP7_75t_L g608 ( .A(n_565), .B(n_609), .Y(n_608) );
AOI322xp5_ASAP7_75t_L g717 ( .A1(n_565), .A2(n_634), .A3(n_641), .B1(n_718), .B2(n_719), .C1(n_720), .C2(n_723), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_565), .B(n_593), .Y(n_735) );
A2O1A1Ixp33_ASAP7_75t_SL g741 ( .A1(n_565), .A2(n_593), .B(n_742), .C(n_744), .Y(n_741) );
AOI221xp5_ASAP7_75t_L g580 ( .A1(n_566), .A2(n_581), .B1(n_586), .B2(n_589), .C(n_592), .Y(n_580) );
INVx1_ASAP7_75t_L g673 ( .A(n_566), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_566), .B(n_722), .Y(n_721) );
OAI22xp33_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_570), .B1(n_573), .B2(n_575), .Y(n_567) );
INVx1_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g650 ( .A(n_571), .B(n_585), .Y(n_650) );
AND2x2_ASAP7_75t_L g708 ( .A(n_571), .B(n_709), .Y(n_708) );
OR2x2_ASAP7_75t_L g616 ( .A(n_572), .B(n_579), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_572), .B(n_585), .Y(n_644) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_574), .B(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_574), .B(n_652), .Y(n_706) );
OAI321xp33_ASAP7_75t_L g725 ( .A1(n_574), .A2(n_647), .A3(n_726), .B1(n_727), .B2(n_728), .C(n_729), .Y(n_725) );
INVx1_ASAP7_75t_L g692 ( .A(n_575), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_576), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g631 ( .A(n_576), .B(n_579), .Y(n_631) );
AOI321xp33_ASAP7_75t_L g689 ( .A1(n_576), .A2(n_593), .A3(n_690), .B1(n_691), .B2(n_692), .C(n_693), .Y(n_689) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g606 ( .A(n_578), .B(n_591), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_579), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_579), .B(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_579), .B(n_665), .Y(n_702) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x4_ASAP7_75t_L g625 ( .A(n_583), .B(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g590 ( .A(n_584), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g698 ( .A(n_585), .Y(n_698) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_588), .B(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g621 ( .A(n_593), .Y(n_621) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_595), .B(n_630), .Y(n_679) );
OR2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
OR2x2_ASAP7_75t_L g643 ( .A(n_598), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_SL g688 ( .A(n_598), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_599), .A2(n_646), .B1(n_649), .B2(n_651), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx1_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g743 ( .A(n_602), .B(n_666), .Y(n_743) );
AOI221xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_607), .B1(n_611), .B2(n_617), .C(n_620), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
BUFx2_ASAP7_75t_L g641 ( .A(n_610), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
INVx1_ASAP7_75t_SL g687 ( .A(n_613), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_615), .B(n_665), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_615), .A2(n_683), .B(n_685), .Y(n_682) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OR2x2_ASAP7_75t_L g728 ( .A(n_616), .B(n_710), .Y(n_728) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_SL g630 ( .A(n_619), .Y(n_630) );
AOI21xp33_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_622), .B(n_624), .Y(n_620) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g674 ( .A(n_626), .B(n_675), .Y(n_674) );
INVxp67_ASAP7_75t_L g736 ( .A(n_626), .Y(n_736) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_631), .B(n_632), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_630), .B(n_648), .Y(n_684) );
INVxp67_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g705 ( .A(n_634), .Y(n_705) );
NAND5xp2_ASAP7_75t_L g635 ( .A(n_636), .B(n_653), .C(n_662), .D(n_682), .E(n_689), .Y(n_635) );
O2A1O1Ixp33_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_639), .B(n_642), .C(n_645), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g677 ( .A(n_641), .Y(n_677) );
CKINVDCx16_ASAP7_75t_R g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_649), .B(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g691 ( .A(n_651), .Y(n_691) );
OAI21xp5_ASAP7_75t_SL g653 ( .A1(n_654), .A2(n_657), .B(n_659), .Y(n_653) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_654), .A2(n_708), .B1(n_711), .B2(n_713), .C(n_714), .Y(n_707) );
AND2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
AOI321xp33_ASAP7_75t_L g662 ( .A1(n_655), .A2(n_663), .A3(n_667), .B1(n_668), .B2(n_674), .C(n_676), .Y(n_662) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g733 ( .A(n_667), .Y(n_733) );
NAND2xp5_ASAP7_75t_SL g668 ( .A(n_669), .B(n_673), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g685 ( .A(n_670), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
NOR2xp67_ASAP7_75t_SL g697 ( .A(n_671), .B(n_678), .Y(n_697) );
AOI321xp33_ASAP7_75t_SL g729 ( .A1(n_674), .A2(n_730), .A3(n_731), .B1(n_732), .B2(n_733), .C(n_734), .Y(n_729) );
O2A1O1Ixp33_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_678), .B(n_679), .C(n_680), .Y(n_676) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_687), .B(n_695), .Y(n_724) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
NAND3xp33_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .C(n_699), .Y(n_696) );
NOR3xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_725), .C(n_737), .Y(n_700) );
OAI211xp5_ASAP7_75t_SL g701 ( .A1(n_702), .A2(n_703), .B(n_707), .C(n_717), .Y(n_701) );
INVxp67_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_705), .B(n_706), .Y(n_704) );
OAI221xp5_ASAP7_75t_L g737 ( .A1(n_706), .A2(n_738), .B1(n_739), .B2(n_740), .C(n_741), .Y(n_737) );
INVx1_ASAP7_75t_L g726 ( .A(n_708), .Y(n_726) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g730 ( .A(n_728), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
CKINVDCx14_ASAP7_75t_R g742 ( .A(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
INVx3_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_SL g771 ( .A(n_765), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
INVx1_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
endmodule