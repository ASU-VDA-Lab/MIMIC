module fake_jpeg_5281_n_214 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_214);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_214;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_2),
.B(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_36),
.Y(n_53)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

AND2x2_ASAP7_75t_SL g34 ( 
.A(n_27),
.B(n_6),
.Y(n_34)
);

NAND2x1p5_ASAP7_75t_L g84 ( 
.A(n_34),
.B(n_13),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_42),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_39),
.A2(n_40),
.B1(n_24),
.B2(n_7),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_21),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_41),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_5),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_17),
.B(n_5),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_46),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_22),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_34),
.A2(n_21),
.B1(n_20),
.B2(n_25),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_49),
.A2(n_83),
.B(n_76),
.C(n_75),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_20),
.B1(n_28),
.B2(n_25),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_51),
.A2(n_56),
.B1(n_61),
.B2(n_78),
.Y(n_100)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_52),
.B(n_55),
.Y(n_112)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_32),
.A2(n_28),
.B1(n_16),
.B2(n_18),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_65),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_48),
.A2(n_18),
.B1(n_29),
.B2(n_30),
.Y(n_61)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_67),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_69),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_29),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_36),
.B(n_15),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_71),
.Y(n_108)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_15),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_73),
.Y(n_88)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_31),
.B(n_30),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_80),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_44),
.A2(n_24),
.B(n_17),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_10),
.C(n_12),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_41),
.A2(n_26),
.B1(n_23),
.B2(n_13),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_23),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_79),
.B(n_86),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_26),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_83),
.B1(n_76),
.B2(n_75),
.Y(n_102)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_82),
.A2(n_83),
.B1(n_87),
.B2(n_63),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_45),
.A2(n_13),
.B1(n_27),
.B2(n_0),
.Y(n_83)
);

OR2x2_ASAP7_75t_SL g99 ( 
.A(n_84),
.B(n_83),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_43),
.B(n_7),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_34),
.A2(n_22),
.B1(n_8),
.B2(n_9),
.Y(n_87)
);

AND2x6_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_9),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_109),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_84),
.A2(n_10),
.B1(n_12),
.B2(n_0),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_93),
.A2(n_101),
.B1(n_102),
.B2(n_110),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_94),
.B(n_99),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_12),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_77),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_59),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_104),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_53),
.B(n_60),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_58),
.B(n_66),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_105),
.B(n_85),
.Y(n_122)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_66),
.B(n_82),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_63),
.A2(n_71),
.B1(n_62),
.B2(n_54),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_111),
.A2(n_50),
.B1(n_54),
.B2(n_62),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_58),
.B(n_52),
.C(n_67),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_73),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_112),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_115),
.Y(n_143)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_108),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_118),
.Y(n_145)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_125),
.Y(n_153)
);

AOI21xp33_ASAP7_75t_L g120 ( 
.A1(n_97),
.A2(n_67),
.B(n_73),
.Y(n_120)
);

AOI21xp33_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_131),
.B(n_109),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_121),
.A2(n_124),
.B1(n_100),
.B2(n_109),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_113),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_90),
.A2(n_50),
.B1(n_85),
.B2(n_73),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_67),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_126),
.B(n_128),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_103),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_92),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_133),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_96),
.B(n_92),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_91),
.Y(n_134)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_91),
.Y(n_136)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_94),
.B(n_104),
.Y(n_137)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_107),
.Y(n_138)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_99),
.B1(n_102),
.B2(n_101),
.Y(n_140)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_138),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_144),
.Y(n_170)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_148),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_159),
.B(n_126),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_129),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_140),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_150),
.B(n_155),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_116),
.B(n_105),
.Y(n_152)
);

NAND3xp33_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_135),
.C(n_127),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_107),
.Y(n_154)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_103),
.Y(n_157)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_157),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_130),
.B(n_133),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_157),
.Y(n_163)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_166),
.B(n_168),
.Y(n_175)
);

AO21x1_ASAP7_75t_L g181 ( 
.A1(n_167),
.A2(n_173),
.B(n_151),
.Y(n_181)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_169),
.A2(n_171),
.B1(n_141),
.B2(n_142),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_146),
.A2(n_125),
.B1(n_115),
.B2(n_118),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_150),
.A2(n_119),
.B(n_137),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_172),
.A2(n_148),
.B(n_159),
.Y(n_177)
);

NAND2xp67_ASAP7_75t_SL g173 ( 
.A(n_139),
.B(n_135),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_123),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_155),
.C(n_152),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_178),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_177),
.A2(n_182),
.B(n_185),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_168),
.B(n_128),
.Y(n_179)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_179),
.Y(n_191)
);

AOI31xp67_ASAP7_75t_L g190 ( 
.A1(n_181),
.A2(n_173),
.A3(n_165),
.B(n_166),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_160),
.C(n_151),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_160),
.A2(n_149),
.B1(n_132),
.B2(n_153),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_183),
.A2(n_184),
.B1(n_139),
.B2(n_124),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_123),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_170),
.B(n_141),
.Y(n_186)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_186),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_187),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_180),
.A2(n_170),
.B1(n_144),
.B2(n_158),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_189),
.A2(n_190),
.B(n_145),
.Y(n_200)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_142),
.Y(n_197)
);

INVxp33_ASAP7_75t_L g195 ( 
.A(n_190),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_195),
.A2(n_197),
.B(n_200),
.Y(n_203)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_198),
.B(n_162),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_176),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_178),
.Y(n_204)
);

OAI31xp33_ASAP7_75t_L g201 ( 
.A1(n_195),
.A2(n_181),
.A3(n_177),
.B(n_183),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_202),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_196),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_205),
.Y(n_208)
);

AOI322xp5_ASAP7_75t_L g206 ( 
.A1(n_203),
.A2(n_199),
.A3(n_194),
.B1(n_185),
.B2(n_162),
.C1(n_182),
.C2(n_191),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_161),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_201),
.A2(n_161),
.B(n_143),
.C(n_192),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_207),
.A2(n_158),
.B1(n_143),
.B2(n_122),
.Y(n_212)
);

AOI211xp5_ASAP7_75t_L g213 ( 
.A1(n_210),
.A2(n_212),
.B(n_206),
.C(n_208),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_209),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_213),
.B(n_211),
.Y(n_214)
);


endmodule