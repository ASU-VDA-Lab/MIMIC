module fake_jpeg_37_n_596 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_596);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_596;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_8),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_12),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g173 ( 
.A(n_60),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_23),
.B(n_18),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_61),
.B(n_74),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_62),
.Y(n_152)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_19),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_64),
.B(n_72),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_65),
.Y(n_161)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_66),
.Y(n_147)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_40),
.Y(n_67)
);

INVx5_ASAP7_75t_SL g134 ( 
.A(n_67),
.Y(n_134)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_68),
.Y(n_139)
);

BUFx16f_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_70),
.Y(n_162)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_26),
.B(n_18),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_28),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_73),
.B(n_93),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_26),
.B(n_18),
.Y(n_74)
);

BUFx16f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_75),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_76),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_24),
.Y(n_77)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_79),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_29),
.B(n_1),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_80),
.B(n_82),
.Y(n_148)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_1),
.Y(n_82)
);

BUFx10_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_84),
.Y(n_193)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_44),
.B(n_2),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_86),
.B(n_91),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_87),
.Y(n_167)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_88),
.Y(n_178)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_29),
.B(n_2),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_92),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_47),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_95),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_32),
.B(n_3),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_96),
.B(n_103),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_97),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_98),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_99),
.Y(n_172)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_39),
.Y(n_102)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_102),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_33),
.B(n_3),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_104),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_34),
.Y(n_105)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_106),
.Y(n_169)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_36),
.Y(n_107)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_107),
.Y(n_179)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_108),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_47),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_112),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_111),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_57),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_114),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_57),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_120),
.Y(n_164)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_32),
.Y(n_116)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_116),
.Y(n_182)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_48),
.Y(n_117)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_117),
.Y(n_183)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_32),
.Y(n_118)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_118),
.Y(n_194)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_49),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_34),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_58),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_36),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_121),
.B(n_122),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_37),
.B(n_3),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_123),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_96),
.A2(n_51),
.B1(n_49),
.B2(n_58),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_125),
.A2(n_146),
.B1(n_170),
.B2(n_167),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_82),
.A2(n_51),
.B1(n_49),
.B2(n_58),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_133),
.A2(n_138),
.B1(n_141),
.B2(n_145),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_86),
.A2(n_51),
.B1(n_58),
.B2(n_45),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_67),
.A2(n_34),
.B1(n_45),
.B2(n_43),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_143),
.B(n_136),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_117),
.A2(n_34),
.B1(n_41),
.B2(n_38),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_89),
.A2(n_27),
.B1(n_56),
.B2(n_55),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_77),
.A2(n_43),
.B1(n_41),
.B2(n_38),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_154),
.A2(n_156),
.B1(n_158),
.B2(n_159),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_95),
.A2(n_70),
.B1(n_92),
.B2(n_62),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_72),
.A2(n_37),
.B1(n_56),
.B2(n_55),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_105),
.A2(n_20),
.B1(n_53),
.B2(n_50),
.Y(n_159)
);

OA22x2_ASAP7_75t_L g165 ( 
.A1(n_116),
.A2(n_52),
.B1(n_59),
.B2(n_21),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_165),
.B(n_186),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_65),
.A2(n_20),
.B1(n_53),
.B2(n_50),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_69),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_181),
.B(n_185),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_122),
.B(n_59),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_66),
.B(n_46),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_118),
.B(n_46),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_187),
.B(n_191),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_119),
.B(n_42),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_78),
.A2(n_85),
.B1(n_90),
.B2(n_42),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_192),
.B(n_156),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_76),
.A2(n_35),
.B1(n_27),
.B2(n_25),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_196),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_81),
.A2(n_35),
.B1(n_25),
.B2(n_21),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_197),
.A2(n_198),
.B1(n_88),
.B2(n_71),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_108),
.A2(n_52),
.B1(n_5),
.B2(n_6),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_60),
.B(n_4),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_200),
.B(n_201),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_60),
.B(n_4),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_94),
.B(n_16),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_202),
.B(n_9),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_203),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_84),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_204),
.B(n_205),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_126),
.B(n_99),
.Y(n_205)
);

INVx11_ASAP7_75t_L g206 ( 
.A(n_134),
.Y(n_206)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_206),
.Y(n_332)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_147),
.Y(n_207)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_207),
.Y(n_280)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_208),
.Y(n_299)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

INVx3_ASAP7_75t_SL g304 ( 
.A(n_209),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_186),
.A2(n_69),
.B(n_75),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_211),
.A2(n_244),
.B(n_145),
.Y(n_282)
);

BUFx5_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

INVx4_ASAP7_75t_SL g283 ( 
.A(n_212),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_149),
.B(n_97),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_213),
.B(n_223),
.Y(n_312)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_128),
.Y(n_214)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_214),
.Y(n_298)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_215),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_168),
.B(n_114),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_216),
.B(n_234),
.Y(n_324)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_129),
.Y(n_217)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_217),
.Y(n_277)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_157),
.Y(n_218)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_218),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_155),
.A2(n_102),
.B1(n_79),
.B2(n_68),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_219),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_125),
.A2(n_113),
.B1(n_111),
.B2(n_104),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_220),
.A2(n_272),
.B1(n_274),
.B2(n_195),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_150),
.B(n_75),
.C(n_83),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_221),
.B(n_261),
.C(n_180),
.Y(n_288)
);

AND2x4_ASAP7_75t_L g222 ( 
.A(n_143),
.B(n_83),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_222),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_169),
.B(n_94),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_132),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_225),
.B(n_230),
.Y(n_278)
);

BUFx12f_ASAP7_75t_L g226 ( 
.A(n_153),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_226),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_184),
.A2(n_102),
.B1(n_87),
.B2(n_123),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_227),
.Y(n_331)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_130),
.Y(n_228)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_228),
.Y(n_305)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_182),
.Y(n_229)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_229),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_142),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_135),
.Y(n_231)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_231),
.Y(n_285)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_194),
.Y(n_232)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_232),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_148),
.B(n_5),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_164),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_235),
.B(n_255),
.Y(n_286)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_140),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_237),
.B(n_239),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_179),
.B(n_8),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_238),
.B(n_247),
.Y(n_302)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_151),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_131),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_240),
.B(n_241),
.Y(n_292)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_131),
.Y(n_241)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_139),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_242),
.B(n_243),
.Y(n_294)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_160),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_159),
.A2(n_109),
.B(n_98),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_163),
.B(n_8),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_245),
.B(n_256),
.Y(n_281)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_139),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_246),
.B(n_251),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_249),
.A2(n_253),
.B1(n_167),
.B2(n_175),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_127),
.B(n_9),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_250),
.B(n_252),
.Y(n_314)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_172),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_137),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_133),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_253)
);

A2O1A1Ixp33_ASAP7_75t_L g254 ( 
.A1(n_165),
.A2(n_10),
.B(n_13),
.C(n_15),
.Y(n_254)
);

A2O1A1Ixp33_ASAP7_75t_L g279 ( 
.A1(n_254),
.A2(n_262),
.B(n_198),
.C(n_141),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_146),
.B(n_170),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_165),
.B(n_10),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_176),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_257),
.Y(n_276)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_124),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_258),
.B(n_267),
.Y(n_319)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_137),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_259),
.Y(n_295)
);

AND2x2_ASAP7_75t_SL g261 ( 
.A(n_183),
.B(n_13),
.Y(n_261)
);

A2O1A1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_197),
.A2(n_15),
.B(n_16),
.C(n_196),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_176),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_263),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_154),
.B(n_15),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_264),
.B(n_270),
.Y(n_321)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_136),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_265),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_152),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_266),
.Y(n_317)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_152),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_134),
.B(n_135),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_268),
.A2(n_269),
.B1(n_144),
.B2(n_180),
.Y(n_301)
);

BUFx8_ASAP7_75t_L g269 ( 
.A(n_173),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_161),
.Y(n_270)
);

AND2x2_ASAP7_75t_SL g309 ( 
.A(n_271),
.B(n_178),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_188),
.B(n_174),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_166),
.Y(n_284)
);

AO21x1_ASAP7_75t_L g356 ( 
.A1(n_279),
.A2(n_282),
.B(n_307),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_284),
.B(n_242),
.Y(n_345)
);

NAND3xp33_ASAP7_75t_L g364 ( 
.A(n_288),
.B(n_269),
.C(n_212),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_297),
.A2(n_308),
.B1(n_316),
.B2(n_320),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_216),
.B(n_199),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_300),
.B(n_311),
.C(n_226),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_301),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_244),
.A2(n_199),
.B(n_124),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_303),
.A2(n_322),
.B(n_330),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_256),
.A2(n_178),
.B1(n_162),
.B2(n_166),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_248),
.A2(n_195),
.B1(n_162),
.B2(n_175),
.Y(n_308)
);

CKINVDCx14_ASAP7_75t_R g360 ( 
.A(n_309),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_214),
.B(n_173),
.C(n_161),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_210),
.A2(n_274),
.B1(n_272),
.B2(n_233),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_313),
.A2(n_315),
.B1(n_318),
.B2(n_325),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_210),
.A2(n_173),
.B1(n_190),
.B2(n_260),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_264),
.A2(n_261),
.B1(n_253),
.B2(n_245),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_236),
.A2(n_190),
.B1(n_234),
.B2(n_254),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_262),
.A2(n_211),
.B(n_271),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_261),
.A2(n_271),
.B1(n_207),
.B2(n_249),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_222),
.A2(n_229),
.B1(n_232),
.B2(n_252),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_327),
.A2(n_334),
.B1(n_208),
.B2(n_226),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_259),
.A2(n_263),
.B1(n_267),
.B2(n_270),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_328),
.A2(n_266),
.B1(n_246),
.B2(n_215),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_221),
.A2(n_222),
.B(n_251),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_222),
.A2(n_217),
.B1(n_218),
.B2(n_209),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_280),
.Y(n_335)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_335),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_287),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_336),
.B(n_350),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_282),
.A2(n_322),
.B(n_303),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_337),
.A2(n_362),
.B(n_381),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_324),
.B(n_225),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_338),
.B(n_339),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_324),
.B(n_243),
.Y(n_339)
);

AO22x1_ASAP7_75t_L g340 ( 
.A1(n_313),
.A2(n_206),
.B1(n_241),
.B2(n_258),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_340),
.B(n_359),
.Y(n_418)
);

BUFx5_ASAP7_75t_L g341 ( 
.A(n_277),
.Y(n_341)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_341),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_300),
.B(n_224),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_343),
.B(n_354),
.C(n_311),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_281),
.B(n_239),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_344),
.B(n_345),
.Y(n_391)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_280),
.Y(n_346)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_346),
.Y(n_389)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_298),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_347),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_310),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_348),
.A2(n_283),
.B1(n_332),
.B2(n_317),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_287),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_281),
.B(n_237),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_351),
.B(n_352),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_284),
.B(n_228),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_298),
.Y(n_353)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_353),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_288),
.B(n_240),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_289),
.B(n_265),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_355),
.B(n_365),
.Y(n_384)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_304),
.Y(n_358)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_358),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_361),
.A2(n_379),
.B1(n_334),
.B2(n_319),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_291),
.A2(n_269),
.B(n_231),
.Y(n_362)
);

OAI21xp33_ASAP7_75t_L g400 ( 
.A1(n_364),
.A2(n_306),
.B(n_299),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_292),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_278),
.B(n_226),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_366),
.B(n_369),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_310),
.Y(n_367)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_367),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_368),
.B(n_326),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_286),
.B(n_312),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_326),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_370),
.B(n_380),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_318),
.B(n_296),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_371),
.B(n_374),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_325),
.A2(n_308),
.B1(n_321),
.B2(n_279),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_372),
.A2(n_373),
.B1(n_376),
.B2(n_309),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_321),
.A2(n_297),
.B1(n_275),
.B2(n_330),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_296),
.B(n_276),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_323),
.Y(n_375)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_375),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_275),
.A2(n_307),
.B1(n_331),
.B2(n_314),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_323),
.Y(n_377)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_377),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_276),
.B(n_333),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_378),
.B(n_295),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_327),
.A2(n_331),
.B1(n_309),
.B2(n_293),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_289),
.B(n_312),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_293),
.A2(n_319),
.B(n_332),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_383),
.A2(n_388),
.B1(n_398),
.B2(n_403),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_374),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_385),
.B(n_407),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_390),
.B(n_340),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_L g436 ( 
.A1(n_393),
.A2(n_283),
.B1(n_370),
.B2(n_363),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_338),
.B(n_302),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_395),
.B(n_404),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_349),
.A2(n_301),
.B1(n_317),
.B2(n_333),
.Y(n_398)
);

OAI32xp33_ASAP7_75t_L g399 ( 
.A1(n_371),
.A2(n_351),
.A3(n_344),
.B1(n_339),
.B2(n_349),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_399),
.B(n_411),
.Y(n_428)
);

OAI21xp33_ASAP7_75t_L g429 ( 
.A1(n_400),
.A2(n_381),
.B(n_379),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_372),
.A2(n_295),
.B1(n_306),
.B2(n_294),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_354),
.B(n_292),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_343),
.B(n_292),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_410),
.B(n_415),
.C(n_416),
.Y(n_432)
);

OAI32xp33_ASAP7_75t_L g412 ( 
.A1(n_363),
.A2(n_305),
.A3(n_294),
.B1(n_326),
.B2(n_287),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_412),
.B(n_417),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_378),
.B(n_329),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_413),
.B(n_304),
.Y(n_426)
);

FAx1_ASAP7_75t_SL g414 ( 
.A(n_337),
.B(n_328),
.CI(n_294),
.CON(n_414),
.SN(n_414)
);

FAx1_ASAP7_75t_SL g433 ( 
.A(n_414),
.B(n_360),
.CI(n_362),
.CON(n_433),
.SN(n_433)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_368),
.B(n_342),
.C(n_352),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_336),
.B(n_305),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_350),
.B(n_347),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_419),
.B(n_353),
.Y(n_424)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_335),
.Y(n_421)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_421),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_402),
.A2(n_342),
.B(n_356),
.Y(n_422)
);

AO21x1_ASAP7_75t_L g465 ( 
.A1(n_422),
.A2(n_433),
.B(n_437),
.Y(n_465)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_424),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_426),
.B(n_429),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_427),
.B(n_438),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_407),
.A2(n_373),
.B1(n_357),
.B2(n_376),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_430),
.A2(n_449),
.B1(n_450),
.B2(n_418),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_431),
.B(n_441),
.C(n_443),
.Y(n_459)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_411),
.Y(n_435)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_435),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_436),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_402),
.A2(n_356),
.B(n_340),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_409),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_382),
.A2(n_346),
.B(n_375),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_439),
.A2(n_420),
.B(n_405),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_397),
.B(n_285),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g477 ( 
.A(n_440),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_416),
.B(n_377),
.C(n_361),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_390),
.B(n_410),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_442),
.B(n_401),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_415),
.B(n_299),
.C(n_277),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_409),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_444),
.B(n_448),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_404),
.B(n_395),
.C(n_386),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_445),
.B(n_447),
.C(n_454),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_408),
.B(n_285),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_446),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_386),
.B(n_399),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_391),
.B(n_358),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_383),
.A2(n_359),
.B1(n_348),
.B2(n_367),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_418),
.A2(n_394),
.B1(n_391),
.B2(n_388),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_387),
.B(n_290),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_451),
.B(n_455),
.Y(n_481)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_406),
.Y(n_453)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_453),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_394),
.B(n_290),
.C(n_283),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_417),
.B(n_304),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_384),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_456),
.B(n_479),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_430),
.A2(n_398),
.B1(n_403),
.B2(n_419),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_457),
.A2(n_460),
.B1(n_462),
.B2(n_467),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_434),
.A2(n_418),
.B1(n_414),
.B2(n_412),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_434),
.A2(n_414),
.B1(n_421),
.B2(n_406),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_452),
.A2(n_392),
.B1(n_389),
.B2(n_396),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_469),
.B(n_455),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_432),
.B(n_431),
.C(n_443),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_471),
.B(n_476),
.C(n_441),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_439),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_474),
.B(n_475),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_424),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_451),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_478),
.B(n_483),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_432),
.B(n_401),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_450),
.A2(n_405),
.B1(n_420),
.B2(n_348),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_480),
.A2(n_485),
.B1(n_444),
.B2(n_438),
.Y(n_486)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_482),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_422),
.A2(n_310),
.B(n_341),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_445),
.B(n_425),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_484),
.B(n_476),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_452),
.A2(n_435),
.B1(n_428),
.B2(n_449),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_486),
.A2(n_493),
.B1(n_470),
.B2(n_504),
.Y(n_526)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_487),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_488),
.B(n_494),
.C(n_502),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_479),
.B(n_447),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_490),
.B(n_510),
.Y(n_523)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_468),
.Y(n_491)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_491),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_456),
.B(n_448),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_492),
.B(n_464),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_462),
.A2(n_428),
.B1(n_437),
.B2(n_433),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_471),
.B(n_425),
.C(n_454),
.Y(n_494)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_470),
.Y(n_496)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_496),
.Y(n_519)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_468),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_498),
.B(n_503),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_458),
.B(n_426),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_499),
.Y(n_514)
);

FAx1_ASAP7_75t_SL g500 ( 
.A(n_465),
.B(n_433),
.CI(n_423),
.CON(n_500),
.SN(n_500)
);

FAx1_ASAP7_75t_SL g518 ( 
.A(n_500),
.B(n_509),
.CI(n_511),
.CON(n_518),
.SN(n_518)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_459),
.B(n_423),
.C(n_453),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_461),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_505),
.B(n_506),
.C(n_509),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_459),
.B(n_463),
.C(n_484),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_458),
.B(n_469),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_507),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_461),
.B(n_482),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_508),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_463),
.B(n_466),
.C(n_467),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_481),
.B(n_466),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_460),
.B(n_485),
.C(n_483),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_511),
.B(n_490),
.C(n_494),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_489),
.A2(n_465),
.B(n_472),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g548 ( 
.A1(n_513),
.A2(n_524),
.B(n_514),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_493),
.A2(n_473),
.B1(n_457),
.B2(n_477),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_517),
.B(n_526),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_518),
.B(n_532),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_507),
.A2(n_473),
.B1(n_480),
.B2(n_481),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_521),
.A2(n_527),
.B1(n_510),
.B2(n_496),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_525),
.B(n_529),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_491),
.A2(n_498),
.B1(n_487),
.B2(n_503),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_502),
.B(n_488),
.C(n_506),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_530),
.B(n_528),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_497),
.Y(n_531)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_531),
.Y(n_543)
);

AO22x1_ASAP7_75t_L g532 ( 
.A1(n_486),
.A2(n_489),
.B1(n_501),
.B2(n_500),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_508),
.Y(n_533)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_533),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_526),
.B(n_505),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_534),
.B(n_535),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_529),
.B(n_495),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_530),
.B(n_520),
.C(n_528),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_536),
.B(n_538),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_515),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_SL g539 ( 
.A(n_531),
.B(n_499),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_539),
.B(n_542),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_540),
.A2(n_549),
.B1(n_522),
.B2(n_516),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_523),
.B(n_520),
.Y(n_542)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_519),
.Y(n_546)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_546),
.B(n_547),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_513),
.A2(n_500),
.B(n_495),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_548),
.B(n_550),
.Y(n_557)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_519),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_540),
.A2(n_517),
.B1(n_514),
.B2(n_524),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_551),
.B(n_555),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_541),
.A2(n_522),
.B1(n_516),
.B2(n_512),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_545),
.B(n_532),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_558),
.B(n_560),
.Y(n_566)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_559),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_534),
.B(n_532),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_541),
.A2(n_527),
.B1(n_521),
.B2(n_512),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_561),
.A2(n_544),
.B1(n_546),
.B2(n_549),
.Y(n_569)
);

INVx6_ASAP7_75t_L g562 ( 
.A(n_536),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_562),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_543),
.A2(n_533),
.B1(n_515),
.B2(n_518),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_563),
.B(n_564),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_SL g564 ( 
.A1(n_548),
.A2(n_518),
.B(n_547),
.Y(n_564)
);

NAND3xp33_ASAP7_75t_L g567 ( 
.A(n_553),
.B(n_552),
.C(n_562),
.Y(n_567)
);

NAND3xp33_ASAP7_75t_L g581 ( 
.A(n_567),
.B(n_556),
.C(n_551),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_569),
.B(n_572),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_557),
.B(n_543),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_557),
.B(n_537),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_573),
.B(n_574),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_554),
.B(n_535),
.C(n_537),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_554),
.B(n_544),
.C(n_560),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_575),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_568),
.B(n_558),
.Y(n_576)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_576),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_SL g577 ( 
.A(n_571),
.B(n_555),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_577),
.B(n_579),
.Y(n_585)
);

OAI21xp5_ASAP7_75t_SL g579 ( 
.A1(n_570),
.A2(n_556),
.B(n_561),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g587 ( 
.A(n_581),
.Y(n_587)
);

OAI211xp5_ASAP7_75t_L g583 ( 
.A1(n_565),
.A2(n_566),
.B(n_575),
.C(n_574),
.Y(n_583)
);

INVxp67_ASAP7_75t_SL g588 ( 
.A(n_583),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_578),
.B(n_566),
.C(n_565),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_L g591 ( 
.A1(n_584),
.A2(n_569),
.B(n_588),
.Y(n_591)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_586),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_589),
.B(n_590),
.Y(n_592)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_587),
.A2(n_582),
.B(n_580),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_591),
.B(n_588),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_593),
.Y(n_594)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_594),
.B(n_585),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_595),
.B(n_592),
.Y(n_596)
);


endmodule