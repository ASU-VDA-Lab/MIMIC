module fake_jpeg_8820_n_63 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_63);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_63;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_55;
wire n_27;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

INVx2_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_9),
.B(n_10),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_13),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_25),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_35),
.B1(n_32),
.B2(n_33),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_1),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_37),
.C(n_3),
.Y(n_40)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_26),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_5),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_21),
.B1(n_17),
.B2(n_18),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_2),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_4),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_40),
.B(n_41),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_36),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_48),
.B(n_49),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_32),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

AND2x6_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_19),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_54),
.B(n_44),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_51),
.Y(n_57)
);

MAJx2_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_57),
.C(n_52),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_55),
.B(n_50),
.Y(n_60)
);

AOI322xp5_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_50),
.A3(n_51),
.B1(n_53),
.B2(n_42),
.C1(n_45),
.C2(n_27),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_46),
.C(n_7),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_SL g63 ( 
.A1(n_62),
.A2(n_6),
.B(n_14),
.C(n_15),
.Y(n_63)
);


endmodule