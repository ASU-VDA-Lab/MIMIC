module fake_jpeg_18322_n_269 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_269);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_269;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_21;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_11),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_11),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_35),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_34),
.Y(n_46)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_40),
.B(n_31),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_22),
.Y(n_42)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_48),
.A2(n_56),
.B1(n_64),
.B2(n_46),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_34),
.C(n_27),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_54),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_30),
.B(n_33),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_SL g72 ( 
.A(n_52),
.B(n_58),
.C(n_44),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_28),
.B1(n_35),
.B2(n_20),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_39),
.B1(n_36),
.B2(n_46),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_30),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_55),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_20),
.B1(n_35),
.B2(n_19),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_20),
.B1(n_28),
.B2(n_15),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_62),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_37),
.B(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_63),
.Y(n_79)
);

OAI32xp33_ASAP7_75t_L g63 ( 
.A1(n_37),
.A2(n_17),
.A3(n_12),
.B1(n_13),
.B2(n_24),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_23),
.B1(n_19),
.B2(n_17),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_23),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_22),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_72),
.A2(n_75),
.B1(n_56),
.B2(n_65),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_39),
.B1(n_36),
.B2(n_44),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_73),
.A2(n_52),
.B1(n_59),
.B2(n_50),
.Y(n_101)
);

BUFx4f_ASAP7_75t_SL g74 ( 
.A(n_59),
.Y(n_74)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_39),
.B1(n_36),
.B2(n_46),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_76),
.A2(n_82),
.B1(n_83),
.B2(n_57),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_13),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_68),
.Y(n_86)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_47),
.B1(n_44),
.B2(n_33),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_65),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_79),
.B(n_51),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_97),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_92),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_55),
.B(n_54),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_89),
.A2(n_95),
.B(n_77),
.Y(n_106)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_99),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_91),
.A2(n_77),
.B1(n_58),
.B2(n_72),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_61),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_51),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_96),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_L g95 ( 
.A1(n_68),
.A2(n_54),
.B(n_55),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_51),
.Y(n_97)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_101),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_104),
.A2(n_106),
.B(n_116),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_86),
.B(n_93),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_109),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_98),
.A2(n_75),
.B1(n_49),
.B2(n_71),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_123),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_96),
.B(n_84),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_71),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_122),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_55),
.B(n_54),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_115),
.A2(n_106),
.B(n_112),
.Y(n_129)
);

NAND2xp33_ASAP7_75t_SL g116 ( 
.A(n_94),
.B(n_58),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_49),
.C(n_73),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_47),
.C(n_99),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_53),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_101),
.A2(n_64),
.B1(n_65),
.B2(n_48),
.Y(n_123)
);

AO21x2_ASAP7_75t_L g124 ( 
.A1(n_87),
.A2(n_67),
.B(n_45),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_102),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_119),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_126),
.B(n_128),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_107),
.A2(n_87),
.B1(n_102),
.B2(n_90),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_135),
.B(n_115),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_88),
.Y(n_130)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_131),
.A2(n_45),
.B1(n_67),
.B2(n_17),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_88),
.Y(n_132)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_100),
.B(n_78),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_113),
.C(n_124),
.Y(n_153)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_147),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_22),
.Y(n_139)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_139),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_74),
.Y(n_140)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_124),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_142),
.B(n_146),
.Y(n_150)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_32),
.Y(n_144)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_32),
.Y(n_145)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_74),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_104),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_125),
.B(n_114),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_152),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_160),
.C(n_166),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_124),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_154),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_137),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_155),
.B(n_158),
.Y(n_189)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_124),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_45),
.C(n_32),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_74),
.Y(n_164)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_164),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_78),
.Y(n_165)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_45),
.C(n_27),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_137),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_168),
.B(n_149),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_134),
.A2(n_0),
.B(n_1),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_169),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_48),
.B1(n_24),
.B2(n_12),
.Y(n_170)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_171),
.A2(n_128),
.B1(n_141),
.B2(n_146),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_133),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_174),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_161),
.A2(n_127),
.B1(n_142),
.B2(n_131),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_178),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_133),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_147),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_175),
.B(n_134),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_158),
.A2(n_127),
.B1(n_130),
.B2(n_145),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_133),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_180),
.B(n_139),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_181),
.A2(n_191),
.B1(n_163),
.B2(n_149),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_148),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_183),
.B(n_184),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_150),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_156),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_186),
.B(n_156),
.Y(n_206)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_190),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_154),
.A2(n_144),
.B1(n_132),
.B2(n_126),
.Y(n_191)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_192),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_189),
.Y(n_195)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_195),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_207),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_182),
.A2(n_135),
.B(n_169),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_198),
.A2(n_171),
.B(n_138),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_159),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_200),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_159),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_201),
.A2(n_173),
.B1(n_154),
.B2(n_157),
.Y(n_217)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_202),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_176),
.Y(n_204)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_206),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_175),
.B(n_166),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_160),
.C(n_157),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_209),
.C(n_180),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_203),
.A2(n_163),
.B1(n_179),
.B2(n_181),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_213),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_197),
.A2(n_177),
.B1(n_188),
.B2(n_185),
.Y(n_213)
);

INVxp67_ASAP7_75t_SL g214 ( 
.A(n_194),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_214),
.Y(n_232)
);

AO221x1_ASAP7_75t_L g215 ( 
.A1(n_205),
.A2(n_178),
.B1(n_141),
.B2(n_138),
.C(n_177),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_215),
.A2(n_217),
.B(n_210),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_196),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_219),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_222),
.A2(n_223),
.B(n_12),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_195),
.A2(n_7),
.B(n_10),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_208),
.C(n_193),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_226),
.C(n_234),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_207),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_225),
.B(n_233),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_193),
.C(n_209),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_228),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_220),
.B(n_16),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_230),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_235),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_212),
.A2(n_221),
.B(n_214),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_227),
.A2(n_21),
.B1(n_14),
.B2(n_10),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_240),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_230),
.A2(n_9),
.B1(n_7),
.B2(n_2),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_224),
.B(n_9),
.Y(n_241)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_241),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_9),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_3),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_225),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_2),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_237),
.A2(n_234),
.B(n_226),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_236),
.C(n_245),
.Y(n_254)
);

AOI21x1_ASAP7_75t_L g248 ( 
.A1(n_243),
.A2(n_0),
.B(n_2),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_248),
.B(n_252),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_251),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_3),
.B(n_4),
.Y(n_251)
);

NOR2xp67_ASAP7_75t_SL g253 ( 
.A(n_236),
.B(n_16),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_16),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_255),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_239),
.C(n_14),
.Y(n_255)
);

OAI21x1_ASAP7_75t_L g262 ( 
.A1(n_257),
.A2(n_259),
.B(n_21),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_14),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_258),
.A2(n_256),
.B(n_21),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_260),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_262),
.A2(n_256),
.B1(n_261),
.B2(n_21),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_264),
.A2(n_4),
.B(n_5),
.Y(n_265)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_265),
.B(n_263),
.C(n_5),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_266),
.A2(n_5),
.B(n_6),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_267),
.B(n_5),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_268),
.A2(n_6),
.B(n_249),
.Y(n_269)
);


endmodule