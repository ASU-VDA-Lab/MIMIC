module fake_jpeg_11827_n_565 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_565);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_565;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx3_ASAP7_75t_SL g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_5),
.B(n_3),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_7),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_61),
.B(n_64),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_63),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_66),
.B(n_74),
.Y(n_145)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_67),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_68),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_69),
.Y(n_176)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_70),
.Y(n_149)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_71),
.Y(n_188)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_72),
.Y(n_150)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_43),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_17),
.B(n_7),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_75),
.B(n_76),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_25),
.B(n_7),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_77),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_35),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_78),
.B(n_83),
.Y(n_172)
);

INVx11_ASAP7_75t_SL g79 ( 
.A(n_35),
.Y(n_79)
);

INVx4_ASAP7_75t_SL g163 ( 
.A(n_79),
.Y(n_163)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_80),
.Y(n_195)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_82),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_6),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_17),
.B(n_8),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_84),
.B(n_85),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_35),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_86),
.Y(n_158)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_87),
.Y(n_175)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_88),
.Y(n_151)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_89),
.Y(n_162)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_90),
.Y(n_161)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_91),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_94),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_96),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_31),
.B(n_16),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_97),
.B(n_98),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_31),
.B(n_5),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_99),
.Y(n_190)
);

BUFx12_ASAP7_75t_L g100 ( 
.A(n_21),
.Y(n_100)
);

INVx6_ASAP7_75t_SL g191 ( 
.A(n_100),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_34),
.B(n_4),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_101),
.B(n_109),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_34),
.B(n_39),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_117),
.Y(n_128)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_21),
.Y(n_103)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_45),
.B(n_4),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_104),
.B(n_122),
.Y(n_186)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_32),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_107),
.Y(n_179)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_39),
.B(n_4),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_20),
.Y(n_111)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_111),
.Y(n_194)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_40),
.Y(n_112)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_112),
.Y(n_184)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_22),
.Y(n_113)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_51),
.Y(n_114)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_32),
.Y(n_115)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_115),
.Y(n_170)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_22),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_20),
.Y(n_118)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_53),
.Y(n_119)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_119),
.Y(n_196)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_120),
.Y(n_197)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_38),
.Y(n_121)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_20),
.B(n_10),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_41),
.B(n_3),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_14),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_100),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_126),
.B(n_56),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_104),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_133),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g202 ( 
.A(n_135),
.Y(n_202)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_152),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_61),
.A2(n_57),
.B1(n_54),
.B2(n_32),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_153),
.A2(n_166),
.B1(n_169),
.B2(n_26),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_155),
.B(n_171),
.Y(n_216)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_95),
.Y(n_165)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_71),
.A2(n_54),
.B1(n_42),
.B2(n_41),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_73),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_167),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_69),
.A2(n_54),
.B1(n_55),
.B2(n_38),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_122),
.B(n_43),
.Y(n_171)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_110),
.Y(n_173)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_173),
.Y(n_262)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_111),
.Y(n_174)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_174),
.Y(n_256)
);

INVx11_ASAP7_75t_L g178 ( 
.A(n_63),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g253 ( 
.A(n_178),
.Y(n_253)
);

BUFx12f_ASAP7_75t_L g180 ( 
.A(n_73),
.Y(n_180)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_180),
.Y(n_214)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_181),
.Y(n_269)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_110),
.Y(n_182)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_79),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_183),
.B(n_48),
.Y(n_225)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_80),
.Y(n_185)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_87),
.Y(n_187)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g193 ( 
.A(n_67),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g265 ( 
.A(n_193),
.Y(n_265)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_93),
.Y(n_198)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_198),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_114),
.B(n_56),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_48),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_162),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_203),
.B(n_222),
.Y(n_282)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_211),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_176),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_212),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_55),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_215),
.B(n_223),
.Y(n_324)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_143),
.Y(n_217)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_217),
.Y(n_288)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_139),
.Y(n_218)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_218),
.Y(n_299)
);

OR2x2_ASAP7_75t_SL g219 ( 
.A(n_186),
.B(n_138),
.Y(n_219)
);

NAND2xp33_ASAP7_75t_SL g314 ( 
.A(n_219),
.B(n_252),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_169),
.A2(n_91),
.B1(n_105),
.B2(n_68),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_220),
.A2(n_242),
.B1(n_190),
.B2(n_154),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_128),
.B(n_51),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_221),
.B(n_224),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_50),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_172),
.B(n_50),
.Y(n_224)
);

INVxp67_ASAP7_75t_SL g283 ( 
.A(n_225),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_172),
.B(n_42),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_226),
.B(n_227),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_159),
.B(n_56),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_127),
.Y(n_228)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_228),
.Y(n_274)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_131),
.Y(n_229)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_229),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_168),
.B(n_138),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_230),
.B(n_239),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_168),
.B(n_28),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_231),
.B(n_243),
.Y(n_301)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_176),
.Y(n_232)
);

INVx3_ASAP7_75t_SL g290 ( 
.A(n_232),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_189),
.Y(n_233)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_233),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_234),
.B(n_260),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_150),
.A2(n_60),
.B1(n_62),
.B2(n_82),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_235),
.A2(n_244),
.B1(n_246),
.B2(n_254),
.Y(n_312)
);

CKINVDCx12_ASAP7_75t_R g236 ( 
.A(n_163),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_236),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_189),
.Y(n_237)
);

INVx3_ASAP7_75t_SL g303 ( 
.A(n_237),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_186),
.B(n_56),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_238),
.B(n_156),
.C(n_157),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_145),
.B(n_49),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_145),
.B(n_49),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_240),
.B(n_245),
.Y(n_291)
);

A2O1A1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_201),
.A2(n_100),
.B(n_28),
.C(n_26),
.Y(n_241)
);

OAI32xp33_ASAP7_75t_L g300 ( 
.A1(n_241),
.A2(n_129),
.A3(n_164),
.B1(n_194),
.B2(n_175),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_201),
.B(n_23),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_158),
.A2(n_115),
.B1(n_106),
.B2(n_99),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_161),
.B(n_23),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_179),
.A2(n_96),
.B1(n_92),
.B2(n_77),
.Y(n_246)
);

CKINVDCx12_ASAP7_75t_R g247 ( 
.A(n_163),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_247),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_184),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_248),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_160),
.A2(n_37),
.B1(n_52),
.B2(n_38),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_249),
.A2(n_257),
.B1(n_266),
.B2(n_129),
.Y(n_308)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_146),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_250),
.Y(n_285)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_146),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_251),
.Y(n_297)
);

INVx13_ASAP7_75t_L g252 ( 
.A(n_183),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_196),
.A2(n_37),
.B1(n_44),
.B2(n_52),
.Y(n_254)
);

INVx8_ASAP7_75t_L g255 ( 
.A(n_125),
.Y(n_255)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_255),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_160),
.A2(n_44),
.B1(n_11),
.B2(n_3),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_125),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_258),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_197),
.A2(n_44),
.B1(n_11),
.B2(n_13),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_259),
.A2(n_261),
.B1(n_205),
.B2(n_255),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_149),
.B(n_11),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_192),
.A2(n_13),
.B1(n_14),
.B2(n_2),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_144),
.B(n_0),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_263),
.B(n_2),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_124),
.B(n_0),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_264),
.B(n_267),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_167),
.B(n_180),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_134),
.B(n_0),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_137),
.B(n_1),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_268),
.B(n_2),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_200),
.A2(n_151),
.B1(n_177),
.B2(n_170),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_270),
.A2(n_136),
.B(n_141),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_230),
.B(n_148),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_273),
.B(n_278),
.Y(n_350)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_229),
.Y(n_279)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_279),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_SL g280 ( 
.A(n_219),
.B(n_140),
.C(n_132),
.Y(n_280)
);

NOR2x1_ASAP7_75t_L g329 ( 
.A(n_280),
.B(n_234),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_281),
.B(n_292),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_242),
.A2(n_190),
.B1(n_130),
.B2(n_147),
.Y(n_287)
);

OAI22xp33_ASAP7_75t_L g325 ( 
.A1(n_287),
.A2(n_232),
.B1(n_258),
.B2(n_237),
.Y(n_325)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_210),
.Y(n_289)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_289),
.Y(n_342)
);

OAI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_221),
.A2(n_188),
.B1(n_195),
.B2(n_142),
.Y(n_293)
);

OA22x2_ASAP7_75t_L g359 ( 
.A1(n_293),
.A2(n_296),
.B1(n_320),
.B2(n_323),
.Y(n_359)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_210),
.Y(n_295)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_295),
.Y(n_344)
);

OA22x2_ASAP7_75t_L g296 ( 
.A1(n_241),
.A2(n_130),
.B1(n_147),
.B2(n_195),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_239),
.A2(n_175),
.B1(n_188),
.B2(n_154),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g347 ( 
.A1(n_298),
.A2(n_311),
.B1(n_250),
.B2(n_251),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_300),
.B(n_296),
.Y(n_346)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_213),
.Y(n_305)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_305),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_306),
.B(n_315),
.Y(n_339)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_213),
.Y(n_307)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_307),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_308),
.Y(n_336)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_217),
.Y(n_310)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_310),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_240),
.A2(n_2),
.B1(n_164),
.B2(n_245),
.Y(n_311)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_228),
.Y(n_317)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_317),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_270),
.A2(n_234),
.B(n_238),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_318),
.A2(n_214),
.B(n_262),
.Y(n_354)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_256),
.Y(n_319)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_319),
.Y(n_365)
);

OAI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_205),
.A2(n_211),
.B1(n_218),
.B2(n_207),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_269),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_322),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g398 ( 
.A1(n_325),
.A2(n_284),
.B1(n_302),
.B2(n_277),
.Y(n_398)
);

INVx6_ASAP7_75t_SL g326 ( 
.A(n_309),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_326),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_216),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_327),
.B(n_328),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_208),
.Y(n_328)
);

OAI21xp33_ASAP7_75t_SL g366 ( 
.A1(n_329),
.A2(n_346),
.B(n_347),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_321),
.Y(n_330)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_330),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_299),
.Y(n_331)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_331),
.Y(n_392)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_274),
.Y(n_332)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_332),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_312),
.A2(n_264),
.B1(n_267),
.B2(n_233),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_333),
.A2(n_345),
.B1(n_298),
.B2(n_311),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_299),
.Y(n_334)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_334),
.Y(n_382)
);

O2A1O1Ixp33_ASAP7_75t_L g335 ( 
.A1(n_278),
.A2(n_252),
.B(n_238),
.C(n_253),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_335),
.B(n_354),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_282),
.B(n_209),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_337),
.B(n_341),
.Y(n_386)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_276),
.Y(n_340)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_340),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_294),
.B(n_209),
.Y(n_341)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_274),
.Y(n_343)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_343),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_312),
.A2(n_212),
.B1(n_207),
.B2(n_253),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_285),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_349),
.B(n_358),
.Y(n_393)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_317),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_356),
.B(n_360),
.Y(n_371)
);

INVx13_ASAP7_75t_L g357 ( 
.A(n_309),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_357),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_297),
.Y(n_358)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_276),
.Y(n_360)
);

A2O1A1Ixp33_ASAP7_75t_L g361 ( 
.A1(n_271),
.A2(n_202),
.B(n_262),
.C(n_208),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_361),
.B(n_364),
.Y(n_372)
);

INVx13_ASAP7_75t_L g363 ( 
.A(n_275),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_363),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_304),
.B(n_204),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_367),
.B(n_375),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_350),
.A2(n_300),
.B1(n_296),
.B2(n_272),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_368),
.A2(n_387),
.B1(n_390),
.B2(n_399),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_350),
.B(n_273),
.C(n_314),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_370),
.B(n_377),
.C(n_378),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_364),
.B(n_304),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_350),
.B(n_271),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_329),
.B(n_292),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_352),
.B(n_280),
.C(n_272),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_381),
.B(n_389),
.C(n_395),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_346),
.A2(n_323),
.B1(n_296),
.B2(n_318),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_383),
.A2(n_388),
.B1(n_339),
.B2(n_359),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_352),
.A2(n_272),
.B1(n_283),
.B2(n_291),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_336),
.A2(n_286),
.B1(n_291),
.B2(n_306),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_329),
.B(n_301),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_352),
.A2(n_315),
.B1(n_277),
.B2(n_290),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_333),
.B(n_315),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_391),
.B(n_353),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_354),
.B(n_322),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_336),
.B(n_319),
.C(n_279),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_396),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_362),
.B(n_289),
.C(n_295),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_397),
.B(n_349),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_398),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_345),
.A2(n_290),
.B1(n_303),
.B2(n_321),
.Y(n_399)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_393),
.Y(n_401)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_401),
.Y(n_441)
);

BUFx12_ASAP7_75t_L g402 ( 
.A(n_380),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_402),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_368),
.A2(n_359),
.B1(n_335),
.B2(n_362),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_403),
.A2(n_429),
.B1(n_390),
.B2(n_392),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_404),
.B(n_410),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_374),
.B(n_358),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_406),
.B(n_411),
.Y(n_451)
);

INVx4_ASAP7_75t_L g407 ( 
.A(n_376),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_407),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_385),
.A2(n_361),
.B(n_326),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_408),
.Y(n_439)
);

AND2x6_ASAP7_75t_L g409 ( 
.A(n_366),
.B(n_359),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_409),
.B(n_417),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_369),
.B(n_355),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_385),
.A2(n_359),
.B(n_284),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_412),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_385),
.A2(n_355),
.B(n_356),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_413),
.A2(n_310),
.B(n_288),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_384),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_414),
.Y(n_447)
);

OAI32xp33_ASAP7_75t_L g417 ( 
.A1(n_372),
.A2(n_332),
.A3(n_343),
.B1(n_365),
.B2(n_339),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_386),
.B(n_365),
.Y(n_419)
);

NOR3xp33_ASAP7_75t_L g435 ( 
.A(n_419),
.B(n_391),
.C(n_381),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_420),
.B(n_422),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_397),
.B(n_348),
.Y(n_421)
);

NAND3xp33_ASAP7_75t_L g445 ( 
.A(n_421),
.B(n_357),
.C(n_363),
.Y(n_445)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_371),
.Y(n_422)
);

INVx13_ASAP7_75t_L g423 ( 
.A(n_371),
.Y(n_423)
);

INVx8_ASAP7_75t_L g449 ( 
.A(n_423),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_372),
.A2(n_342),
.B(n_338),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_424),
.A2(n_396),
.B(n_388),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_375),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_426),
.B(n_427),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_392),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_383),
.A2(n_325),
.B1(n_351),
.B2(n_342),
.Y(n_428)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_428),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_367),
.A2(n_338),
.B1(n_353),
.B2(n_351),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_379),
.B(n_394),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_430),
.B(n_307),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_435),
.B(n_436),
.Y(n_469)
);

A2O1A1Ixp33_ASAP7_75t_L g436 ( 
.A1(n_412),
.A2(n_377),
.B(n_370),
.C(n_395),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_437),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g438 ( 
.A(n_418),
.B(n_378),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_438),
.B(n_450),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_440),
.A2(n_443),
.B1(n_444),
.B2(n_400),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_403),
.A2(n_387),
.B1(n_389),
.B2(n_373),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_405),
.A2(n_382),
.B1(n_373),
.B2(n_399),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_445),
.B(n_454),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_418),
.B(n_344),
.C(n_348),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_446),
.B(n_452),
.C(n_410),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_425),
.B(n_344),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_425),
.B(n_305),
.Y(n_452)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_453),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_408),
.A2(n_360),
.B(n_340),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_413),
.B(n_406),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_455),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_456),
.B(n_427),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_448),
.A2(n_405),
.B1(n_416),
.B2(n_429),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_460),
.A2(n_472),
.B1(n_443),
.B2(n_440),
.Y(n_488)
);

FAx1_ASAP7_75t_SL g461 ( 
.A(n_436),
.B(n_426),
.CI(n_420),
.CON(n_461),
.SN(n_461)
);

FAx1_ASAP7_75t_SL g492 ( 
.A(n_461),
.B(n_467),
.CI(n_469),
.CON(n_492),
.SN(n_492)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_462),
.B(n_473),
.C(n_474),
.Y(n_486)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_442),
.Y(n_463)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_463),
.Y(n_484)
);

BUFx5_ASAP7_75t_L g464 ( 
.A(n_434),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_464),
.B(n_466),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_SL g467 ( 
.A(n_431),
.B(n_421),
.C(n_416),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_432),
.B(n_419),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_468),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_450),
.B(n_404),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_470),
.B(n_478),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_457),
.B(n_422),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_471),
.B(n_477),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_448),
.A2(n_415),
.B1(n_401),
.B2(n_409),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_446),
.B(n_424),
.C(n_430),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_438),
.B(n_411),
.C(n_428),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_432),
.B(n_407),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_475),
.A2(n_476),
.B1(n_463),
.B2(n_459),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_441),
.B(n_407),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_441),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_447),
.B(n_417),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_479),
.A2(n_458),
.B1(n_456),
.B2(n_423),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_452),
.B(n_414),
.C(n_400),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_482),
.B(n_455),
.C(n_439),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_485),
.B(n_487),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_469),
.A2(n_431),
.B(n_439),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_488),
.A2(n_489),
.B1(n_490),
.B2(n_493),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_460),
.A2(n_433),
.B1(n_437),
.B2(n_444),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_465),
.A2(n_451),
.B1(n_449),
.B2(n_447),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_491),
.B(n_503),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_492),
.B(n_494),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_472),
.A2(n_458),
.B1(n_409),
.B2(n_451),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_462),
.B(n_455),
.C(n_454),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_495),
.B(n_502),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_479),
.A2(n_449),
.B1(n_434),
.B2(n_423),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_496),
.B(n_501),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_478),
.A2(n_330),
.B1(n_402),
.B2(n_303),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_473),
.B(n_474),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_481),
.B(n_470),
.C(n_482),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_494),
.A2(n_467),
.B(n_483),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_504),
.A2(n_510),
.B(n_491),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_486),
.B(n_481),
.C(n_483),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_505),
.B(n_507),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_497),
.B(n_459),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_506),
.B(n_519),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_492),
.B(n_461),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_486),
.B(n_480),
.C(n_471),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_509),
.B(n_510),
.C(n_517),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_502),
.B(n_477),
.C(n_461),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_489),
.A2(n_402),
.B1(n_330),
.B2(n_464),
.Y(n_514)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_514),
.Y(n_525)
);

O2A1O1Ixp33_ASAP7_75t_L g515 ( 
.A1(n_500),
.A2(n_402),
.B(n_253),
.C(n_265),
.Y(n_515)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_515),
.Y(n_532)
);

A2O1A1Ixp33_ASAP7_75t_SL g517 ( 
.A1(n_487),
.A2(n_402),
.B(n_265),
.C(n_214),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_500),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_508),
.B(n_492),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_520),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_513),
.A2(n_493),
.B1(n_488),
.B2(n_484),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_521),
.B(n_523),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_511),
.B(n_503),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_522),
.B(n_529),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_SL g523 ( 
.A1(n_517),
.A2(n_484),
.B1(n_499),
.B2(n_501),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_518),
.B(n_498),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_528),
.B(n_531),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_511),
.B(n_498),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_530),
.B(n_516),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_509),
.A2(n_496),
.B1(n_495),
.B2(n_316),
.Y(n_531)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_535),
.B(n_539),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_524),
.B(n_512),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_536),
.B(n_538),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_521),
.B(n_512),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_529),
.B(n_505),
.C(n_514),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_526),
.B(n_316),
.Y(n_540)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_540),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_522),
.B(n_515),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_541),
.B(n_526),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_543),
.B(n_517),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_539),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_544),
.A2(n_549),
.B1(n_550),
.B2(n_547),
.Y(n_552)
);

NOR2x1_ASAP7_75t_SL g545 ( 
.A(n_537),
.B(n_520),
.Y(n_545)
);

A2O1A1Ixp33_ASAP7_75t_L g551 ( 
.A1(n_545),
.A2(n_532),
.B(n_517),
.C(n_533),
.Y(n_551)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_542),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_534),
.A2(n_527),
.B1(n_525),
.B2(n_531),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_551),
.B(n_552),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_548),
.B(n_533),
.C(n_535),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_553),
.B(n_554),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_546),
.B(n_530),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_555),
.B(n_543),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_556),
.B(n_288),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_557),
.B(n_554),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_559),
.B(n_560),
.C(n_558),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_561),
.B(n_204),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_562),
.A2(n_206),
.B1(n_202),
.B2(n_265),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_563),
.B(n_202),
.Y(n_564)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_564),
.B(n_206),
.Y(n_565)
);


endmodule