module fake_jpeg_28478_n_157 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_157);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_157;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_40),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_23),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_41),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_25),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_8),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_33),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_1),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_64),
.Y(n_76)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_1),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_69),
.Y(n_77)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_66),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_83),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_51),
.B1(n_54),
.B2(n_60),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_59),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_75),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_42),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_42),
.Y(n_78)
);

FAx1_ASAP7_75t_SL g88 ( 
.A(n_78),
.B(n_48),
.CI(n_61),
.CON(n_88),
.SN(n_88)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_62),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_82),
.A2(n_79),
.B1(n_56),
.B2(n_73),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_52),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_88),
.Y(n_113)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_58),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_94),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_61),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_95),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_55),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_72),
.A2(n_45),
.B1(n_53),
.B2(n_43),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_3),
.Y(n_103)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_72),
.A2(n_54),
.B1(n_51),
.B2(n_26),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_99),
.B1(n_5),
.B2(n_6),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_103),
.A2(n_6),
.B(n_7),
.Y(n_123)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_105),
.A2(n_12),
.B1(n_14),
.B2(n_16),
.Y(n_129)
);

MAJx2_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_27),
.C(n_37),
.Y(n_108)
);

NAND3xp33_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_39),
.C(n_18),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_88),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_115),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_24),
.C(n_36),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_118),
.Y(n_132)
);

INVxp67_ASAP7_75t_SL g111 ( 
.A(n_85),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_111),
.Y(n_126)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_21),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_94),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_101),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_119),
.B(n_123),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_100),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_125),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_125)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_130),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_111),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_109),
.A2(n_28),
.B(n_30),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_134),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_31),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_107),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_135),
.Y(n_141)
);

AOI221xp5_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_107),
.B1(n_113),
.B2(n_103),
.C(n_102),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_144),
.Y(n_148)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_143),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_146),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_128),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_149),
.A2(n_147),
.B(n_131),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_125),
.B(n_136),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_140),
.B(n_137),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_152),
.A2(n_142),
.B(n_138),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_153),
.B(n_126),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_120),
.C(n_148),
.Y(n_155)
);

OAI221xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_127),
.B1(n_132),
.B2(n_130),
.C(n_34),
.Y(n_156)
);

BUFx24_ASAP7_75t_SL g157 ( 
.A(n_156),
.Y(n_157)
);


endmodule