module fake_netlist_5_2035_n_3172 (n_137, n_676, n_294, n_431, n_318, n_380, n_419, n_653, n_611, n_444, n_642, n_469, n_615, n_851, n_82, n_194, n_316, n_785, n_389, n_843, n_549, n_684, n_850, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_705, n_619, n_408, n_61, n_678, n_664, n_376, n_697, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_776, n_667, n_515, n_790, n_57, n_353, n_351, n_367, n_620, n_643, n_452, n_397, n_493, n_111, n_525, n_703, n_698, n_483, n_544, n_683, n_155, n_780, n_649, n_552, n_547, n_43, n_721, n_116, n_841, n_22, n_467, n_564, n_802, n_423, n_840, n_284, n_46, n_245, n_21, n_501, n_823, n_725, n_139, n_38, n_105, n_280, n_744, n_590, n_629, n_672, n_4, n_378, n_551, n_762, n_17, n_581, n_688, n_382, n_554, n_800, n_254, n_690, n_33, n_23, n_583, n_671, n_718, n_819, n_302, n_265, n_526, n_719, n_293, n_372, n_443, n_244, n_677, n_47, n_173, n_821, n_198, n_714, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_625, n_621, n_753, n_100, n_455, n_674, n_417, n_612, n_212, n_385, n_498, n_516, n_788, n_507, n_119, n_497, n_689, n_738, n_606, n_559, n_275, n_640, n_252, n_624, n_825, n_26, n_295, n_133, n_330, n_508, n_739, n_506, n_2, n_737, n_610, n_692, n_755, n_6, n_509, n_568, n_39, n_147, n_373, n_820, n_757, n_67, n_307, n_633, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_758, n_668, n_733, n_375, n_301, n_828, n_779, n_576, n_68, n_804, n_93, n_186, n_537, n_134, n_191, n_587, n_659, n_51, n_63, n_492, n_792, n_563, n_171, n_153, n_756, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_741, n_548, n_543, n_260, n_812, n_842, n_298, n_650, n_320, n_694, n_518, n_505, n_286, n_122, n_282, n_752, n_331, n_10, n_24, n_406, n_519, n_470, n_782, n_325, n_449, n_132, n_90, n_724, n_546, n_101, n_760, n_658, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_731, n_31, n_456, n_13, n_371, n_481, n_535, n_709, n_152, n_540, n_317, n_618, n_9, n_323, n_569, n_769, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_831, n_826, n_335, n_123, n_654, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_833, n_297, n_156, n_5, n_853, n_603, n_225, n_377, n_751, n_484, n_775, n_219, n_442, n_157, n_814, n_131, n_192, n_636, n_786, n_600, n_660, n_223, n_392, n_158, n_655, n_704, n_787, n_138, n_264, n_109, n_669, n_472, n_742, n_750, n_454, n_387, n_771, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_635, n_347, n_763, n_169, n_59, n_522, n_550, n_255, n_696, n_215, n_350, n_196, n_798, n_662, n_459, n_646, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_622, n_723, n_386, n_578, n_287, n_344, n_848, n_555, n_783, n_473, n_422, n_475, n_777, n_72, n_661, n_104, n_41, n_682, n_415, n_56, n_141, n_485, n_496, n_355, n_849, n_486, n_670, n_15, n_816, n_336, n_584, n_681, n_591, n_145, n_48, n_521, n_614, n_663, n_845, n_50, n_337, n_430, n_313, n_631, n_673, n_837, n_88, n_479, n_528, n_510, n_216, n_680, n_168, n_395, n_164, n_432, n_553, n_727, n_839, n_311, n_813, n_830, n_773, n_208, n_142, n_743, n_214, n_328, n_140, n_801, n_299, n_303, n_369, n_675, n_296, n_613, n_241, n_637, n_357, n_598, n_685, n_608, n_184, n_446, n_445, n_65, n_78, n_749, n_829, n_144, n_114, n_96, n_772, n_691, n_717, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_789, n_363, n_402, n_413, n_734, n_638, n_700, n_197, n_796, n_107, n_573, n_69, n_236, n_388, n_761, n_1, n_249, n_740, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_693, n_309, n_30, n_512, n_14, n_836, n_84, n_462, n_130, n_322, n_567, n_258, n_652, n_778, n_29, n_79, n_151, n_25, n_306, n_722, n_458, n_288, n_770, n_188, n_190, n_844, n_201, n_263, n_471, n_609, n_852, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_711, n_781, n_834, n_474, n_112, n_765, n_542, n_85, n_463, n_488, n_595, n_736, n_502, n_239, n_466, n_420, n_630, n_489, n_632, n_699, n_55, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_748, n_586, n_846, n_465, n_838, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_745, n_627, n_767, n_172, n_206, n_217, n_440, n_726, n_478, n_793, n_545, n_441, n_450, n_648, n_312, n_476, n_818, n_429, n_534, n_345, n_210, n_494, n_641, n_628, n_365, n_774, n_91, n_729, n_730, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_647, n_237, n_425, n_513, n_407, n_527, n_679, n_707, n_710, n_795, n_695, n_832, n_180, n_560, n_656, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_665, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_720, n_0, n_58, n_623, n_405, n_824, n_18, n_359, n_490, n_805, n_117, n_326, n_794, n_768, n_233, n_404, n_686, n_205, n_366, n_572, n_113, n_712, n_754, n_847, n_815, n_246, n_596, n_179, n_125, n_410, n_558, n_708, n_269, n_529, n_128, n_735, n_702, n_285, n_822, n_412, n_120, n_232, n_327, n_135, n_657, n_126, n_644, n_728, n_202, n_266, n_272, n_491, n_427, n_791, n_732, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_808, n_409, n_797, n_589, n_716, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_651, n_435, n_809, n_159, n_334, n_599, n_766, n_811, n_541, n_807, n_391, n_701, n_434, n_645, n_539, n_835, n_175, n_538, n_666, n_262, n_803, n_238, n_639, n_799, n_99, n_687, n_715, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_817, n_360, n_36, n_594, n_764, n_200, n_162, n_64, n_759, n_222, n_28, n_89, n_438, n_806, n_115, n_713, n_324, n_810, n_634, n_416, n_199, n_827, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_626, n_11, n_424, n_7, n_706, n_746, n_256, n_305, n_533, n_747, n_52, n_278, n_784, n_110, n_3172);

input n_137;
input n_676;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_653;
input n_611;
input n_444;
input n_642;
input n_469;
input n_615;
input n_851;
input n_82;
input n_194;
input n_316;
input n_785;
input n_389;
input n_843;
input n_549;
input n_684;
input n_850;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_705;
input n_619;
input n_408;
input n_61;
input n_678;
input n_664;
input n_376;
input n_697;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_776;
input n_667;
input n_515;
input n_790;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_643;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_703;
input n_698;
input n_483;
input n_544;
input n_683;
input n_155;
input n_780;
input n_649;
input n_552;
input n_547;
input n_43;
input n_721;
input n_116;
input n_841;
input n_22;
input n_467;
input n_564;
input n_802;
input n_423;
input n_840;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_823;
input n_725;
input n_139;
input n_38;
input n_105;
input n_280;
input n_744;
input n_590;
input n_629;
input n_672;
input n_4;
input n_378;
input n_551;
input n_762;
input n_17;
input n_581;
input n_688;
input n_382;
input n_554;
input n_800;
input n_254;
input n_690;
input n_33;
input n_23;
input n_583;
input n_671;
input n_718;
input n_819;
input n_302;
input n_265;
input n_526;
input n_719;
input n_293;
input n_372;
input n_443;
input n_244;
input n_677;
input n_47;
input n_173;
input n_821;
input n_198;
input n_714;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_625;
input n_621;
input n_753;
input n_100;
input n_455;
input n_674;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_788;
input n_507;
input n_119;
input n_497;
input n_689;
input n_738;
input n_606;
input n_559;
input n_275;
input n_640;
input n_252;
input n_624;
input n_825;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_739;
input n_506;
input n_2;
input n_737;
input n_610;
input n_692;
input n_755;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_820;
input n_757;
input n_67;
input n_307;
input n_633;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_758;
input n_668;
input n_733;
input n_375;
input n_301;
input n_828;
input n_779;
input n_576;
input n_68;
input n_804;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_659;
input n_51;
input n_63;
input n_492;
input n_792;
input n_563;
input n_171;
input n_153;
input n_756;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_741;
input n_548;
input n_543;
input n_260;
input n_812;
input n_842;
input n_298;
input n_650;
input n_320;
input n_694;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_752;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_782;
input n_325;
input n_449;
input n_132;
input n_90;
input n_724;
input n_546;
input n_101;
input n_760;
input n_658;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_731;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_709;
input n_152;
input n_540;
input n_317;
input n_618;
input n_9;
input n_323;
input n_569;
input n_769;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_831;
input n_826;
input n_335;
input n_123;
input n_654;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_833;
input n_297;
input n_156;
input n_5;
input n_853;
input n_603;
input n_225;
input n_377;
input n_751;
input n_484;
input n_775;
input n_219;
input n_442;
input n_157;
input n_814;
input n_131;
input n_192;
input n_636;
input n_786;
input n_600;
input n_660;
input n_223;
input n_392;
input n_158;
input n_655;
input n_704;
input n_787;
input n_138;
input n_264;
input n_109;
input n_669;
input n_472;
input n_742;
input n_750;
input n_454;
input n_387;
input n_771;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_635;
input n_347;
input n_763;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_696;
input n_215;
input n_350;
input n_196;
input n_798;
input n_662;
input n_459;
input n_646;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_723;
input n_386;
input n_578;
input n_287;
input n_344;
input n_848;
input n_555;
input n_783;
input n_473;
input n_422;
input n_475;
input n_777;
input n_72;
input n_661;
input n_104;
input n_41;
input n_682;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_849;
input n_486;
input n_670;
input n_15;
input n_816;
input n_336;
input n_584;
input n_681;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_663;
input n_845;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_673;
input n_837;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_680;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_727;
input n_839;
input n_311;
input n_813;
input n_830;
input n_773;
input n_208;
input n_142;
input n_743;
input n_214;
input n_328;
input n_140;
input n_801;
input n_299;
input n_303;
input n_369;
input n_675;
input n_296;
input n_613;
input n_241;
input n_637;
input n_357;
input n_598;
input n_685;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_749;
input n_829;
input n_144;
input n_114;
input n_96;
input n_772;
input n_691;
input n_717;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_789;
input n_363;
input n_402;
input n_413;
input n_734;
input n_638;
input n_700;
input n_197;
input n_796;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_761;
input n_1;
input n_249;
input n_740;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_693;
input n_309;
input n_30;
input n_512;
input n_14;
input n_836;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_652;
input n_778;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_722;
input n_458;
input n_288;
input n_770;
input n_188;
input n_190;
input n_844;
input n_201;
input n_263;
input n_471;
input n_609;
input n_852;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_711;
input n_781;
input n_834;
input n_474;
input n_112;
input n_765;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_736;
input n_502;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_632;
input n_699;
input n_55;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_748;
input n_586;
input n_846;
input n_465;
input n_838;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_745;
input n_627;
input n_767;
input n_172;
input n_206;
input n_217;
input n_440;
input n_726;
input n_478;
input n_793;
input n_545;
input n_441;
input n_450;
input n_648;
input n_312;
input n_476;
input n_818;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_641;
input n_628;
input n_365;
input n_774;
input n_91;
input n_729;
input n_730;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_647;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_679;
input n_707;
input n_710;
input n_795;
input n_695;
input n_832;
input n_180;
input n_560;
input n_656;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_665;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_720;
input n_0;
input n_58;
input n_623;
input n_405;
input n_824;
input n_18;
input n_359;
input n_490;
input n_805;
input n_117;
input n_326;
input n_794;
input n_768;
input n_233;
input n_404;
input n_686;
input n_205;
input n_366;
input n_572;
input n_113;
input n_712;
input n_754;
input n_847;
input n_815;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_708;
input n_269;
input n_529;
input n_128;
input n_735;
input n_702;
input n_285;
input n_822;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_657;
input n_126;
input n_644;
input n_728;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_791;
input n_732;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_808;
input n_409;
input n_797;
input n_589;
input n_716;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_651;
input n_435;
input n_809;
input n_159;
input n_334;
input n_599;
input n_766;
input n_811;
input n_541;
input n_807;
input n_391;
input n_701;
input n_434;
input n_645;
input n_539;
input n_835;
input n_175;
input n_538;
input n_666;
input n_262;
input n_803;
input n_238;
input n_639;
input n_799;
input n_99;
input n_687;
input n_715;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_817;
input n_360;
input n_36;
input n_594;
input n_764;
input n_200;
input n_162;
input n_64;
input n_759;
input n_222;
input n_28;
input n_89;
input n_438;
input n_806;
input n_115;
input n_713;
input n_324;
input n_810;
input n_634;
input n_416;
input n_199;
input n_827;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_626;
input n_11;
input n_424;
input n_7;
input n_706;
input n_746;
input n_256;
input n_305;
input n_533;
input n_747;
input n_52;
input n_278;
input n_784;
input n_110;

output n_3172;

wire n_924;
wire n_1263;
wire n_1378;
wire n_977;
wire n_2253;
wire n_2417;
wire n_2756;
wire n_1423;
wire n_1126;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_2617;
wire n_2200;
wire n_3006;
wire n_1161;
wire n_3027;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_3127;
wire n_1780;
wire n_1488;
wire n_2899;
wire n_2955;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_3086;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1360;
wire n_1198;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_3064;
wire n_2391;
wire n_3088;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_2143;
wire n_2853;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_3019;
wire n_3039;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_3163;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1728;
wire n_1107;
wire n_2076;
wire n_2031;
wire n_3036;
wire n_2482;
wire n_2677;
wire n_1230;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_3010;
wire n_2770;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_3107;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2963;
wire n_2142;
wire n_3082;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_3048;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1243;
wire n_1016;
wire n_2959;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_2761;
wire n_1483;
wire n_2888;
wire n_1314;
wire n_1512;
wire n_3157;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_2983;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_3022;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_2715;
wire n_3087;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_2936;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_3060;
wire n_2651;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_3013;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_3049;
wire n_1723;
wire n_955;
wire n_1850;
wire n_3028;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_3156;
wire n_3101;
wire n_897;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_1414;
wire n_1216;
wire n_2693;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_2976;
wire n_926;
wire n_2249;
wire n_2180;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_3089;
wire n_1547;
wire n_1070;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_1561;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_1513;
wire n_2908;
wire n_2970;
wire n_1600;
wire n_2235;
wire n_1862;
wire n_1239;
wire n_2915;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_1587;
wire n_1473;
wire n_2682;
wire n_901;
wire n_2432;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_2934;
wire n_1672;
wire n_2506;
wire n_2699;
wire n_888;
wire n_1880;
wire n_2769;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_2615;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_2985;
wire n_1151;
wire n_2944;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_2932;
wire n_2753;
wire n_2980;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_3136;
wire n_1836;
wire n_2868;
wire n_1450;
wire n_3141;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_3164;
wire n_2738;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_2968;
wire n_1700;
wire n_2833;
wire n_1585;
wire n_2712;
wire n_2684;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_2855;
wire n_2713;
wire n_2644;
wire n_2700;
wire n_1211;
wire n_1197;
wire n_2951;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_3008;
wire n_1447;
wire n_907;
wire n_2251;
wire n_3096;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_3025;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_892;
wire n_3007;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1463;
wire n_1581;
wire n_1002;
wire n_2100;
wire n_3071;
wire n_2258;
wire n_1058;
wire n_1667;
wire n_2784;
wire n_2919;
wire n_3092;
wire n_1053;
wire n_1224;
wire n_2865;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_3146;
wire n_2241;
wire n_2757;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_1385;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_2942;
wire n_2987;
wire n_1527;
wire n_2042;
wire n_3106;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2862;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_1565;
wire n_2828;
wire n_1809;
wire n_1856;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_857;
wire n_2305;
wire n_2636;
wire n_2450;
wire n_1319;
wire n_2379;
wire n_2616;
wire n_2911;
wire n_2154;
wire n_1951;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_2293;
wire n_2837;
wire n_1393;
wire n_2319;
wire n_1775;
wire n_2979;
wire n_2028;
wire n_1368;
wire n_2762;
wire n_2808;
wire n_1276;
wire n_3009;
wire n_2548;
wire n_1412;
wire n_2679;
wire n_1709;
wire n_2676;
wire n_2108;
wire n_1538;
wire n_1162;
wire n_2930;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_3116;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_1038;
wire n_2967;
wire n_1369;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_2698;
wire n_1711;
wire n_870;
wire n_931;
wire n_1891;
wire n_1662;
wire n_1481;
wire n_2626;
wire n_3042;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_3047;
wire n_868;
wire n_2454;
wire n_2804;
wire n_914;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_3120;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_1888;
wire n_2009;
wire n_2222;
wire n_1892;
wire n_2990;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_1477;
wire n_3142;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_3119;
wire n_1189;
wire n_2690;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_1649;
wire n_3150;
wire n_2064;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_2621;
wire n_1759;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_913;
wire n_1537;
wire n_865;
wire n_2227;
wire n_2671;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_1829;
wire n_1464;
wire n_3133;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_2992;
wire n_1674;
wire n_1833;
wire n_3138;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_3128;
wire n_1734;
wire n_3038;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_3068;
wire n_1767;
wire n_3144;
wire n_2943;
wire n_2913;
wire n_2336;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_1233;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_2007;
wire n_949;
wire n_2539;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_2736;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_3158;
wire n_1624;
wire n_3000;
wire n_1510;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_1279;
wire n_1406;
wire n_3108;
wire n_3113;
wire n_3111;
wire n_2718;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_2577;
wire n_1760;
wire n_2875;
wire n_936;
wire n_1500;
wire n_2960;
wire n_1090;
wire n_2796;
wire n_2342;
wire n_2856;
wire n_1832;
wire n_1851;
wire n_999;
wire n_2046;
wire n_2848;
wire n_2741;
wire n_2937;
wire n_3003;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_3095;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_3030;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_2787;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_2846;
wire n_1781;
wire n_2084;
wire n_2925;
wire n_2035;
wire n_2061;
wire n_3075;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_2857;
wire n_1586;
wire n_959;
wire n_2459;
wire n_3031;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_2982;
wire n_1017;
wire n_2481;
wire n_2947;
wire n_2171;
wire n_978;
wire n_2768;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_1079;
wire n_2093;
wire n_2339;
wire n_1045;
wire n_1208;
wire n_2320;
wire n_2038;
wire n_2473;
wire n_2137;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_2029;
wire n_995;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_3021;
wire n_1989;
wire n_2359;
wire n_2941;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_3098;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_2312;
wire n_962;
wire n_1215;
wire n_3015;
wire n_1171;
wire n_1578;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_2882;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_2952;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_3058;
wire n_2812;
wire n_2048;
wire n_3109;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_3002;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_2565;
wire n_1159;
wire n_957;
wire n_2124;
wire n_3001;
wire n_2081;
wire n_3149;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_2418;
wire n_2519;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_2897;
wire n_2909;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_1237;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_2277;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_2090;
wire n_3153;
wire n_3045;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_2896;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_3065;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_3077;
wire n_2681;
wire n_1562;
wire n_3103;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_2878;
wire n_1823;
wire n_874;
wire n_2464;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_987;
wire n_1846;
wire n_3037;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_3154;
wire n_860;
wire n_2849;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_1849;
wire n_2410;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_2922;
wire n_1430;
wire n_2645;
wire n_2467;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_3029;
wire n_1552;
wire n_2508;
wire n_2593;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_2088;
wire n_2953;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_2658;
wire n_1717;
wire n_2895;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_3097;
wire n_1821;
wire n_2929;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_2740;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2890;
wire n_3059;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_3171;
wire n_1229;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2989;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_3026;
wire n_2216;
wire n_3020;
wire n_1757;
wire n_890;
wire n_1897;
wire n_1919;
wire n_1424;
wire n_1056;
wire n_960;
wire n_2933;
wire n_2308;
wire n_1893;
wire n_2910;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_2647;
wire n_3160;
wire n_1311;
wire n_2191;
wire n_2864;
wire n_2969;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_1346;
wire n_3053;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_3130;
wire n_2465;
wire n_2824;
wire n_3033;
wire n_2650;
wire n_912;
wire n_968;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_2923;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_2333;
wire n_885;
wire n_2916;
wire n_3166;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_1632;
wire n_3110;
wire n_2998;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_2402;
wire n_1157;
wire n_3073;
wire n_2403;
wire n_1050;
wire n_1954;
wire n_2265;
wire n_3162;
wire n_1608;
wire n_983;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_2870;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_3134;
wire n_2304;
wire n_2999;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_2637;
wire n_1974;
wire n_2463;
wire n_2086;
wire n_2289;
wire n_3080;
wire n_3051;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_2881;
wire n_1203;
wire n_1631;
wire n_2472;
wire n_1763;
wire n_2341;
wire n_3105;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_2993;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_2309;
wire n_2415;
wire n_2948;
wire n_3041;
wire n_2646;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_2123;
wire n_972;
wire n_2037;
wire n_2685;
wire n_3040;
wire n_1953;
wire n_1938;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_2903;
wire n_1967;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_1312;
wire n_1439;
wire n_2827;
wire n_1688;
wire n_3052;
wire n_945;
wire n_2997;
wire n_1504;
wire n_943;
wire n_992;
wire n_3067;
wire n_1932;
wire n_2755;
wire n_984;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_3167;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_3078;
wire n_2364;
wire n_2533;
wire n_3094;
wire n_896;
wire n_2310;
wire n_2780;
wire n_2287;
wire n_2860;
wire n_2291;
wire n_3099;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_2973;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_2318;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_2974;
wire n_988;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_2707;
wire n_2751;
wire n_2793;
wire n_2971;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_3147;
wire n_2758;
wire n_1458;
wire n_2471;
wire n_1472;
wire n_1176;
wire n_2298;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_2559;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2840;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_2893;
wire n_1188;
wire n_2588;
wire n_2962;
wire n_1722;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_2600;
wire n_2795;
wire n_1638;
wire n_1786;
wire n_2981;
wire n_2002;
wire n_2282;
wire n_2800;
wire n_2371;
wire n_2935;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_2352;
wire n_1413;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_3085;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_1895;
wire n_3123;
wire n_3137;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_939;
wire n_2361;
wire n_1088;
wire n_1173;
wire n_1232;
wire n_1603;
wire n_2638;
wire n_866;
wire n_969;
wire n_1401;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_2949;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_1653;
wire n_2270;
wire n_1506;
wire n_2653;
wire n_990;
wire n_2867;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_1465;
wire n_3145;
wire n_3124;
wire n_1122;
wire n_2608;
wire n_2657;
wire n_2995;
wire n_1375;
wire n_2494;
wire n_2649;
wire n_1102;
wire n_2852;
wire n_2392;
wire n_3093;
wire n_1843;
wire n_1499;
wire n_3061;
wire n_3155;
wire n_1187;
wire n_2633;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_1174;
wire n_2431;
wire n_2835;
wire n_2558;
wire n_1371;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_982;
wire n_2575;
wire n_2988;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_2766;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2722;
wire n_2117;
wire n_2745;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_1410;
wire n_1005;
wire n_1003;
wire n_3090;
wire n_2067;
wire n_1168;
wire n_2219;
wire n_2437;
wire n_2885;
wire n_2877;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_1584;
wire n_1726;
wire n_1835;
wire n_3035;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_2634;
wire n_910;
wire n_2232;
wire n_3034;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_2811;
wire n_1496;
wire n_1125;
wire n_2547;
wire n_3014;
wire n_1812;
wire n_2501;
wire n_3079;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_2121;
wire n_1803;
wire n_2665;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_1533;
wire n_2224;
wire n_2924;
wire n_2484;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_2994;
wire n_1067;
wire n_2946;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_3135;
wire n_2003;
wire n_1457;
wire n_2692;
wire n_3148;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_2264;
wire n_2754;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_872;
wire n_2012;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_2917;
wire n_869;
wire n_2965;
wire n_1703;
wire n_1352;
wire n_2926;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_3046;
wire n_1170;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_2103;
wire n_2160;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_855;
wire n_1178;
wire n_1461;
wire n_2697;
wire n_3074;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_2861;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2549;
wire n_2705;
wire n_3005;
wire n_2332;
wire n_1235;
wire n_980;
wire n_1115;
wire n_2433;
wire n_3129;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_2977;
wire n_2601;
wire n_3043;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_1334;
wire n_1907;
wire n_2686;
wire n_2528;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_2316;
wire n_3055;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_2906;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2817;
wire n_3139;
wire n_2773;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_2687;
wire n_3023;
wire n_1120;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_2850;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_2654;
wire n_997;
wire n_3104;
wire n_932;
wire n_3169;
wire n_3151;
wire n_3131;
wire n_2078;
wire n_1409;
wire n_1326;
wire n_3070;
wire n_2884;
wire n_1268;
wire n_2996;
wire n_2819;
wire n_3126;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_1718;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_1489;
wire n_1922;
wire n_2966;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_2950;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_3140;
wire n_3170;
wire n_2104;
wire n_2748;
wire n_2057;
wire n_3011;
wire n_1772;
wire n_905;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_2717;
wire n_2818;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_1901;
wire n_3069;
wire n_1900;
wire n_1620;
wire n_3032;
wire n_2889;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_3018;
wire n_1675;
wire n_3072;
wire n_1924;
wire n_2573;
wire n_3084;
wire n_3081;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_2939;
wire n_1745;
wire n_2735;
wire n_2497;
wire n_2006;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_3056;
wire n_1221;
wire n_2345;
wire n_2986;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_2726;
wire n_2774;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_3062;
wire n_3161;
wire n_2317;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_3017;
wire n_2476;
wire n_1770;
wire n_2781;
wire n_2456;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_2984;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_930;
wire n_1873;
wire n_1411;
wire n_3054;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_2854;
wire n_994;
wire n_1701;
wire n_2194;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_1567;
wire n_2567;
wire n_1247;
wire n_2709;
wire n_3102;
wire n_922;
wire n_3122;
wire n_1648;
wire n_1536;
wire n_3050;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_1246;
wire n_1478;
wire n_1339;
wire n_1797;
wire n_1769;
wire n_2957;
wire n_1210;
wire n_2964;
wire n_1364;
wire n_2956;
wire n_2357;
wire n_2183;
wire n_2742;
wire n_2673;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_1367;
wire n_928;
wire n_1943;
wire n_1460;
wire n_2018;
wire n_1555;
wire n_3117;
wire n_2834;
wire n_2531;
wire n_1589;
wire n_2961;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_2883;
wire n_3115;
wire n_2208;
wire n_3076;
wire n_1404;
wire n_3063;
wire n_2912;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_2931;
wire n_1652;
wire n_2209;
wire n_2809;
wire n_2050;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_3118;
wire n_2321;
wire n_1226;
wire n_1277;
wire n_2591;
wire n_2146;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_2940;
wire n_1546;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_979;
wire n_1515;
wire n_2841;
wire n_3165;
wire n_1627;
wire n_2918;
wire n_1245;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_2112;
wire n_1739;
wire n_2958;
wire n_2278;
wire n_2594;
wire n_3114;
wire n_3125;
wire n_2394;
wire n_1914;
wire n_2954;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_2381;
wire n_1654;
wire n_3004;
wire n_2569;
wire n_3112;
wire n_2349;
wire n_1103;
wire n_3132;
wire n_1379;
wire n_2734;
wire n_2196;
wire n_3024;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_2404;
wire n_2083;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_2655;
wire n_2027;
wire n_2642;
wire n_1130;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_1604;
wire n_1275;
wire n_2513;
wire n_2525;
wire n_3091;
wire n_2695;
wire n_1764;
wire n_2892;
wire n_3057;
wire n_3066;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1493;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2708;
wire n_2113;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_1996;
wire n_1505;
wire n_1181;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_1340;
wire n_2274;
wire n_2972;
wire n_1558;
wire n_2166;
wire n_2938;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_3152;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_2689;
wire n_2920;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_2991;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_3016;
wire n_1693;
wire n_2975;
wire n_2599;
wire n_2704;
wire n_904;
wire n_2839;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_2802;
wire n_1542;
wire n_1251;
wire n_3159;
wire n_2728;
wire n_2268;

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_426),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_200),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_820),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_727),
.Y(n_857)
);

INVx1_ASAP7_75t_SL g858 ( 
.A(n_822),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_750),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_311),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_747),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_590),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_778),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_29),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_719),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_708),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_798),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_677),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_810),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_836),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_785),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_217),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_723),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_611),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_755),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_63),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_800),
.Y(n_877)
);

CKINVDCx16_ASAP7_75t_R g878 ( 
.A(n_615),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_826),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_705),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_298),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_318),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_766),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_764),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_586),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_552),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_11),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_814),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_756),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_3),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_76),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_578),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_483),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_853),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_619),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_757),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_829),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_768),
.Y(n_898)
);

CKINVDCx16_ASAP7_75t_R g899 ( 
.A(n_452),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_470),
.Y(n_900)
);

INVxp67_ASAP7_75t_SL g901 ( 
.A(n_324),
.Y(n_901)
);

CKINVDCx20_ASAP7_75t_R g902 ( 
.A(n_239),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_155),
.Y(n_903)
);

BUFx10_ASAP7_75t_L g904 ( 
.A(n_667),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_254),
.Y(n_905)
);

CKINVDCx20_ASAP7_75t_R g906 ( 
.A(n_650),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_592),
.Y(n_907)
);

BUFx2_ASAP7_75t_R g908 ( 
.A(n_652),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_307),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_547),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_620),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_0),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_739),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_792),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_93),
.Y(n_915)
);

CKINVDCx16_ASAP7_75t_R g916 ( 
.A(n_195),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_824),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_791),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_74),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_716),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_233),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_453),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_771),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_563),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_348),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_541),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_91),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_752),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_758),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_532),
.Y(n_930)
);

BUFx10_ASAP7_75t_L g931 ( 
.A(n_706),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_219),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_264),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_603),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_720),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_816),
.Y(n_936)
);

CKINVDCx20_ASAP7_75t_R g937 ( 
.A(n_776),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_809),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_738),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_760),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_297),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_842),
.Y(n_942)
);

CKINVDCx20_ASAP7_75t_R g943 ( 
.A(n_0),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_643),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_724),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_321),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_833),
.Y(n_947)
);

CKINVDCx16_ASAP7_75t_R g948 ( 
.A(n_821),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_58),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_335),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_828),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_587),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_781),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_789),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_495),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_812),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_624),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_837),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_367),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_817),
.Y(n_960)
);

BUFx10_ASAP7_75t_L g961 ( 
.A(n_484),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_229),
.Y(n_962)
);

BUFx10_ASAP7_75t_L g963 ( 
.A(n_145),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_210),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_253),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_582),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_385),
.Y(n_967)
);

CKINVDCx20_ASAP7_75t_R g968 ( 
.A(n_285),
.Y(n_968)
);

INVx1_ASAP7_75t_SL g969 ( 
.A(n_273),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_711),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_519),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_725),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_425),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_585),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_288),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_594),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_384),
.Y(n_977)
);

CKINVDCx20_ASAP7_75t_R g978 ( 
.A(n_638),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_712),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_843),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_205),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_438),
.Y(n_982)
);

BUFx5_ASAP7_75t_L g983 ( 
.A(n_575),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_12),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_94),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_364),
.Y(n_986)
);

BUFx2_ASAP7_75t_L g987 ( 
.A(n_818),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_51),
.Y(n_988)
);

BUFx10_ASAP7_75t_L g989 ( 
.A(n_156),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_316),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_782),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_235),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_784),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_437),
.Y(n_994)
);

BUFx5_ASAP7_75t_L g995 ( 
.A(n_713),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_746),
.Y(n_996)
);

CKINVDCx20_ASAP7_75t_R g997 ( 
.A(n_515),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_690),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_763),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_257),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_405),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_408),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_570),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_681),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_762),
.Y(n_1005)
);

BUFx2_ASAP7_75t_L g1006 ( 
.A(n_205),
.Y(n_1006)
);

INVx1_ASAP7_75t_SL g1007 ( 
.A(n_767),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_823),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_275),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_498),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_413),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_749),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_561),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_167),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_802),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_217),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_834),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_308),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_31),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_709),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_170),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_533),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_589),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_194),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_722),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_559),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_795),
.Y(n_1027)
);

BUFx5_ASAP7_75t_L g1028 ( 
.A(n_703),
.Y(n_1028)
);

BUFx2_ASAP7_75t_L g1029 ( 
.A(n_794),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_93),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_148),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_721),
.Y(n_1032)
);

CKINVDCx20_ASAP7_75t_R g1033 ( 
.A(n_526),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_277),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_718),
.Y(n_1035)
);

CKINVDCx20_ASAP7_75t_R g1036 ( 
.A(n_172),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_572),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_71),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_396),
.Y(n_1039)
);

BUFx5_ASAP7_75t_L g1040 ( 
.A(n_54),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_774),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_737),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_120),
.Y(n_1043)
);

CKINVDCx16_ASAP7_75t_R g1044 ( 
.A(n_804),
.Y(n_1044)
);

CKINVDCx20_ASAP7_75t_R g1045 ( 
.A(n_779),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_803),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_717),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_504),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_707),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_398),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_813),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_186),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_819),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_372),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_714),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_206),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_350),
.Y(n_1057)
);

INVx1_ASAP7_75t_SL g1058 ( 
.A(n_844),
.Y(n_1058)
);

CKINVDCx16_ASAP7_75t_R g1059 ( 
.A(n_380),
.Y(n_1059)
);

BUFx2_ASAP7_75t_SL g1060 ( 
.A(n_524),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_132),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_753),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_849),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_754),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_177),
.Y(n_1065)
);

INVx2_ASAP7_75t_SL g1066 ( 
.A(n_790),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_759),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_496),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_769),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_676),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_9),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_773),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_352),
.Y(n_1073)
);

INVx1_ASAP7_75t_SL g1074 ( 
.A(n_831),
.Y(n_1074)
);

CKINVDCx20_ASAP7_75t_R g1075 ( 
.A(n_735),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_144),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_127),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_493),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_748),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_251),
.Y(n_1080)
);

INVx1_ASAP7_75t_SL g1081 ( 
.A(n_281),
.Y(n_1081)
);

BUFx10_ASAP7_75t_L g1082 ( 
.A(n_19),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_775),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_787),
.Y(n_1084)
);

CKINVDCx20_ASAP7_75t_R g1085 ( 
.A(n_772),
.Y(n_1085)
);

BUFx2_ASAP7_75t_L g1086 ( 
.A(n_741),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_740),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_319),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_266),
.Y(n_1089)
);

BUFx2_ASAP7_75t_L g1090 ( 
.A(n_729),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_734),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_190),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_554),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_292),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_22),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_598),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_19),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_731),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_840),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_9),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_505),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_490),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_825),
.Y(n_1103)
);

CKINVDCx14_ASAP7_75t_R g1104 ( 
.A(n_503),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_195),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_845),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_468),
.Y(n_1107)
);

CKINVDCx16_ASAP7_75t_R g1108 ( 
.A(n_374),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_409),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_783),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_797),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_807),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_745),
.Y(n_1113)
);

CKINVDCx20_ASAP7_75t_R g1114 ( 
.A(n_796),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_608),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_124),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_480),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_733),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_673),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_328),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_553),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_520),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_799),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_730),
.Y(n_1124)
);

BUFx10_ASAP7_75t_L g1125 ( 
.A(n_185),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_761),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_67),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_815),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_808),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_688),
.Y(n_1130)
);

CKINVDCx20_ASAP7_75t_R g1131 ( 
.A(n_167),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_732),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_715),
.Y(n_1133)
);

HB1xp67_ASAP7_75t_L g1134 ( 
.A(n_780),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_178),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_221),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_439),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_765),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_62),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_181),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_786),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_147),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_566),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_432),
.Y(n_1144)
);

CKINVDCx20_ASAP7_75t_R g1145 ( 
.A(n_152),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_282),
.Y(n_1146)
);

BUFx10_ASAP7_75t_L g1147 ( 
.A(n_145),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_744),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_743),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_418),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_455),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_306),
.Y(n_1152)
);

BUFx10_ASAP7_75t_L g1153 ( 
.A(n_263),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_164),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_334),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_806),
.Y(n_1156)
);

CKINVDCx20_ASAP7_75t_R g1157 ( 
.A(n_793),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_684),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_699),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_391),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_658),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_105),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_832),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_742),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_125),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_805),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_641),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_101),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_477),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_406),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_830),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_255),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_107),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_55),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_103),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_7),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_363),
.Y(n_1177)
);

INVxp67_ASAP7_75t_L g1178 ( 
.A(n_163),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_269),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_811),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_440),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_751),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_537),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_474),
.Y(n_1184)
);

CKINVDCx20_ASAP7_75t_R g1185 ( 
.A(n_576),
.Y(n_1185)
);

CKINVDCx20_ASAP7_75t_R g1186 ( 
.A(n_846),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_414),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_726),
.Y(n_1188)
);

CKINVDCx14_ASAP7_75t_R g1189 ( 
.A(n_168),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_777),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_354),
.Y(n_1191)
);

CKINVDCx14_ASAP7_75t_R g1192 ( 
.A(n_770),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_839),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_336),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_198),
.Y(n_1195)
);

CKINVDCx16_ASAP7_75t_R g1196 ( 
.A(n_788),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_407),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_693),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_635),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_728),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_331),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_63),
.Y(n_1202)
);

BUFx10_ASAP7_75t_L g1203 ( 
.A(n_534),
.Y(n_1203)
);

INVx2_ASAP7_75t_SL g1204 ( 
.A(n_827),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_127),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_472),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_736),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_654),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_24),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_801),
.Y(n_1210)
);

BUFx2_ASAP7_75t_L g1211 ( 
.A(n_616),
.Y(n_1211)
);

CKINVDCx16_ASAP7_75t_R g1212 ( 
.A(n_710),
.Y(n_1212)
);

INVx1_ASAP7_75t_SL g1213 ( 
.A(n_224),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1040),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1040),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1040),
.Y(n_1216)
);

INVx1_ASAP7_75t_SL g1217 ( 
.A(n_1006),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_854),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1040),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_1189),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_856),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1040),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_964),
.Y(n_1223)
);

INVxp67_ASAP7_75t_SL g1224 ( 
.A(n_870),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_964),
.Y(n_1225)
);

INVxp33_ASAP7_75t_SL g1226 ( 
.A(n_891),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_964),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1052),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_876),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_887),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_859),
.Y(n_1231)
);

BUFx3_ASAP7_75t_L g1232 ( 
.A(n_904),
.Y(n_1232)
);

INVx3_ASAP7_75t_L g1233 ( 
.A(n_963),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_903),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_981),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_984),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_860),
.Y(n_1237)
);

INVxp67_ASAP7_75t_SL g1238 ( 
.A(n_1041),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_988),
.Y(n_1239)
);

INVxp67_ASAP7_75t_SL g1240 ( 
.A(n_1134),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_904),
.Y(n_1241)
);

INVxp67_ASAP7_75t_SL g1242 ( 
.A(n_1149),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_916),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_992),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_861),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1019),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1024),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1061),
.Y(n_1248)
);

INVx1_ASAP7_75t_SL g1249 ( 
.A(n_902),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_906),
.Y(n_1250)
);

INVx3_ASAP7_75t_L g1251 ( 
.A(n_963),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1077),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1116),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1135),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1136),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1139),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1140),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1174),
.Y(n_1258)
);

CKINVDCx14_ASAP7_75t_R g1259 ( 
.A(n_1104),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1202),
.Y(n_1260)
);

CKINVDCx20_ASAP7_75t_R g1261 ( 
.A(n_937),
.Y(n_1261)
);

CKINVDCx16_ASAP7_75t_R g1262 ( 
.A(n_878),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1209),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_855),
.Y(n_1264)
);

INVxp67_ASAP7_75t_SL g1265 ( 
.A(n_1179),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_968),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_983),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_983),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_862),
.Y(n_1269)
);

CKINVDCx14_ASAP7_75t_R g1270 ( 
.A(n_1192),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_978),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_863),
.Y(n_1272)
);

INVxp67_ASAP7_75t_L g1273 ( 
.A(n_989),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_865),
.Y(n_1274)
);

INVxp67_ASAP7_75t_SL g1275 ( 
.A(n_974),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_989),
.Y(n_1276)
);

INVxp33_ASAP7_75t_SL g1277 ( 
.A(n_864),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1082),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_1218),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1223),
.Y(n_1280)
);

CKINVDCx16_ASAP7_75t_R g1281 ( 
.A(n_1250),
.Y(n_1281)
);

OA21x2_ASAP7_75t_L g1282 ( 
.A1(n_1215),
.A2(n_1222),
.B(n_1216),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1220),
.B(n_1211),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1225),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_1227),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1214),
.Y(n_1286)
);

OAI22x1_ASAP7_75t_L g1287 ( 
.A1(n_1217),
.A2(n_1213),
.B1(n_1095),
.B2(n_890),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1269),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1219),
.Y(n_1289)
);

NAND2xp33_ASAP7_75t_L g1290 ( 
.A(n_1264),
.B(n_1221),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1226),
.A2(n_899),
.B1(n_1044),
.B2(n_948),
.Y(n_1291)
);

OA21x2_ASAP7_75t_L g1292 ( 
.A1(n_1274),
.A2(n_873),
.B(n_869),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1231),
.B(n_1066),
.Y(n_1293)
);

OA21x2_ASAP7_75t_L g1294 ( 
.A1(n_1267),
.A2(n_884),
.B(n_880),
.Y(n_1294)
);

OA21x2_ASAP7_75t_L g1295 ( 
.A1(n_1268),
.A2(n_889),
.B(n_886),
.Y(n_1295)
);

BUFx8_ASAP7_75t_L g1296 ( 
.A(n_1276),
.Y(n_1296)
);

OA21x2_ASAP7_75t_L g1297 ( 
.A1(n_1229),
.A2(n_920),
.B(n_900),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1230),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1237),
.B(n_1204),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1277),
.B(n_987),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1245),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1224),
.A2(n_883),
.B(n_857),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_1232),
.Y(n_1303)
);

INVx2_ASAP7_75t_SL g1304 ( 
.A(n_1241),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1259),
.B(n_1029),
.Y(n_1305)
);

INVx2_ASAP7_75t_SL g1306 ( 
.A(n_1233),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1234),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1235),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1272),
.B(n_1086),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1228),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1238),
.A2(n_918),
.B(n_894),
.Y(n_1311)
);

BUFx6f_ASAP7_75t_L g1312 ( 
.A(n_1236),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_1239),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1244),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1246),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1275),
.B(n_1090),
.Y(n_1316)
);

INVx5_ASAP7_75t_L g1317 ( 
.A(n_1233),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1270),
.B(n_1067),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_1247),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1248),
.Y(n_1320)
);

BUFx8_ASAP7_75t_L g1321 ( 
.A(n_1252),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1253),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1240),
.B(n_1121),
.Y(n_1323)
);

AOI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1262),
.A2(n_1108),
.B1(n_1196),
.B2(n_1059),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1254),
.Y(n_1325)
);

BUFx8_ASAP7_75t_L g1326 ( 
.A(n_1255),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1298),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1307),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1286),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1289),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_1313),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1306),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1303),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1308),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_1305),
.Y(n_1335)
);

AOI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1300),
.A2(n_1265),
.B1(n_1242),
.B2(n_1033),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1280),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1315),
.Y(n_1338)
);

NAND2xp33_ASAP7_75t_SL g1339 ( 
.A(n_1291),
.B(n_1243),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1283),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1320),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1325),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1317),
.B(n_1251),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1284),
.Y(n_1344)
);

XNOR2xp5_ASAP7_75t_L g1345 ( 
.A(n_1324),
.B(n_1261),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1288),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1285),
.Y(n_1347)
);

INVx3_ASAP7_75t_L g1348 ( 
.A(n_1312),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1310),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1312),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_L g1351 ( 
.A(n_1319),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1319),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1317),
.B(n_1251),
.Y(n_1353)
);

AND2x6_ASAP7_75t_L g1354 ( 
.A(n_1323),
.B(n_1057),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1287),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1304),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1294),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1314),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1322),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1295),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1282),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1293),
.B(n_1113),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1316),
.B(n_1278),
.Y(n_1363)
);

INVx3_ASAP7_75t_L g1364 ( 
.A(n_1297),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_L g1365 ( 
.A(n_1299),
.B(n_1278),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1309),
.B(n_1273),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1318),
.B(n_1292),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1302),
.B(n_1212),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1311),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1321),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1290),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1326),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1279),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1301),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1296),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1281),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1279),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1298),
.Y(n_1378)
);

INVx3_ASAP7_75t_L g1379 ( 
.A(n_1313),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_SL g1380 ( 
.A(n_1300),
.B(n_931),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1298),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1306),
.B(n_1263),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1298),
.Y(n_1383)
);

AND2x6_ASAP7_75t_L g1384 ( 
.A(n_1305),
.B(n_1057),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1298),
.Y(n_1385)
);

BUFx6f_ASAP7_75t_L g1386 ( 
.A(n_1312),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1298),
.Y(n_1387)
);

OA21x2_ASAP7_75t_L g1388 ( 
.A1(n_1302),
.A2(n_901),
.B(n_924),
.Y(n_1388)
);

XOR2xp5_ASAP7_75t_L g1389 ( 
.A(n_1281),
.B(n_1266),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1286),
.Y(n_1390)
);

CKINVDCx8_ASAP7_75t_R g1391 ( 
.A(n_1281),
.Y(n_1391)
);

BUFx6f_ASAP7_75t_L g1392 ( 
.A(n_1312),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1306),
.B(n_1249),
.Y(n_1393)
);

BUFx2_ASAP7_75t_L g1394 ( 
.A(n_1303),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_SL g1395 ( 
.A(n_1371),
.B(n_1365),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1366),
.B(n_1271),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1329),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1363),
.B(n_926),
.Y(n_1398)
);

INVx3_ASAP7_75t_L g1399 ( 
.A(n_1351),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1336),
.B(n_1393),
.Y(n_1400)
);

INVx1_ASAP7_75t_SL g1401 ( 
.A(n_1394),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1330),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1335),
.B(n_908),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1327),
.Y(n_1404)
);

INVxp67_ASAP7_75t_L g1405 ( 
.A(n_1333),
.Y(n_1405)
);

OR2x6_ASAP7_75t_L g1406 ( 
.A(n_1370),
.B(n_1372),
.Y(n_1406)
);

AND2x6_ASAP7_75t_L g1407 ( 
.A(n_1369),
.B(n_929),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1328),
.Y(n_1408)
);

INVx3_ASAP7_75t_L g1409 ( 
.A(n_1351),
.Y(n_1409)
);

OR2x6_ASAP7_75t_L g1410 ( 
.A(n_1376),
.B(n_1060),
.Y(n_1410)
);

BUFx6f_ASAP7_75t_L g1411 ( 
.A(n_1386),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1361),
.A2(n_1020),
.B1(n_1039),
.B2(n_982),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1334),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1338),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1341),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_SL g1416 ( 
.A(n_1377),
.B(n_997),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1342),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1367),
.A2(n_1101),
.B1(n_1167),
.B2(n_1098),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1390),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1359),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1337),
.Y(n_1421)
);

AND2x4_ASAP7_75t_L g1422 ( 
.A(n_1331),
.B(n_1256),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1346),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1378),
.Y(n_1424)
);

INVx4_ASAP7_75t_L g1425 ( 
.A(n_1392),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_1391),
.Y(n_1426)
);

BUFx2_ASAP7_75t_L g1427 ( 
.A(n_1340),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1380),
.B(n_1260),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1344),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1355),
.Y(n_1430)
);

AOI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1339),
.A2(n_1075),
.B1(n_1085),
.B2(n_1045),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1373),
.Y(n_1432)
);

NAND3xp33_ASAP7_75t_L g1433 ( 
.A(n_1381),
.B(n_905),
.C(n_872),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1383),
.Y(n_1434)
);

BUFx6f_ASAP7_75t_L g1435 ( 
.A(n_1386),
.Y(n_1435)
);

OR2x6_ASAP7_75t_L g1436 ( 
.A(n_1375),
.B(n_1178),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1358),
.Y(n_1437)
);

NAND2xp33_ASAP7_75t_L g1438 ( 
.A(n_1357),
.B(n_1354),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1362),
.B(n_934),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1385),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1387),
.Y(n_1441)
);

INVx2_ASAP7_75t_SL g1442 ( 
.A(n_1382),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1392),
.Y(n_1443)
);

NAND3xp33_ASAP7_75t_L g1444 ( 
.A(n_1332),
.B(n_915),
.C(n_912),
.Y(n_1444)
);

BUFx3_ASAP7_75t_L g1445 ( 
.A(n_1379),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1360),
.A2(n_1193),
.B1(n_939),
.B2(n_951),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1374),
.B(n_1356),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1350),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1352),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1354),
.B(n_950),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1347),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1354),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1357),
.B(n_1364),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1349),
.Y(n_1454)
);

INVx4_ASAP7_75t_L g1455 ( 
.A(n_1348),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1343),
.Y(n_1456)
);

INVx3_ASAP7_75t_L g1457 ( 
.A(n_1353),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1384),
.B(n_953),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1384),
.B(n_954),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1388),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1368),
.Y(n_1461)
);

OR2x6_ASAP7_75t_L g1462 ( 
.A(n_1389),
.B(n_1258),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1384),
.Y(n_1463)
);

INVx5_ASAP7_75t_L g1464 ( 
.A(n_1345),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1329),
.Y(n_1465)
);

INVx2_ASAP7_75t_SL g1466 ( 
.A(n_1393),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1361),
.A2(n_959),
.B1(n_970),
.B2(n_966),
.Y(n_1467)
);

CKINVDCx20_ASAP7_75t_R g1468 ( 
.A(n_1391),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_SL g1469 ( 
.A(n_1371),
.B(n_1093),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1394),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1327),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_SL g1472 ( 
.A(n_1371),
.B(n_1111),
.Y(n_1472)
);

AND2x4_ASAP7_75t_L g1473 ( 
.A(n_1331),
.B(n_1257),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1371),
.A2(n_1157),
.B1(n_1185),
.B2(n_1114),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1365),
.B(n_975),
.Y(n_1475)
);

INVx3_ASAP7_75t_L g1476 ( 
.A(n_1351),
.Y(n_1476)
);

INVx3_ASAP7_75t_L g1477 ( 
.A(n_1351),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1329),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_1371),
.B(n_1186),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1329),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1336),
.B(n_919),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_1371),
.B(n_858),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1365),
.B(n_976),
.Y(n_1483)
);

INVxp33_ASAP7_75t_L g1484 ( 
.A(n_1393),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1371),
.B(n_969),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1327),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1336),
.B(n_921),
.Y(n_1487)
);

INVx5_ASAP7_75t_L g1488 ( 
.A(n_1351),
.Y(n_1488)
);

NAND2xp33_ASAP7_75t_SL g1489 ( 
.A(n_1380),
.B(n_943),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1366),
.B(n_971),
.Y(n_1490)
);

INVx1_ASAP7_75t_SL g1491 ( 
.A(n_1393),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1329),
.Y(n_1492)
);

NOR2x1p5_ASAP7_75t_L g1493 ( 
.A(n_1375),
.B(n_1195),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1393),
.B(n_1082),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1365),
.B(n_977),
.Y(n_1495)
);

NAND3xp33_ASAP7_75t_L g1496 ( 
.A(n_1336),
.B(n_932),
.C(n_927),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1327),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1327),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1361),
.A2(n_990),
.B1(n_1004),
.B2(n_994),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1327),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1365),
.B(n_1009),
.Y(n_1501)
);

AND2x6_ASAP7_75t_L g1502 ( 
.A(n_1369),
.B(n_1010),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_SL g1503 ( 
.A(n_1371),
.B(n_1058),
.Y(n_1503)
);

INVx3_ASAP7_75t_L g1504 ( 
.A(n_1351),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1329),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1327),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1366),
.B(n_1007),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1361),
.A2(n_1015),
.B1(n_1023),
.B2(n_1013),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1351),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1404),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1397),
.Y(n_1511)
);

AOI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1461),
.A2(n_1081),
.B1(n_1074),
.B2(n_1035),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1402),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1484),
.B(n_1014),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1490),
.B(n_1025),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1507),
.B(n_1047),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1395),
.B(n_1054),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1470),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1475),
.B(n_1055),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1419),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1483),
.B(n_1063),
.Y(n_1521)
);

INVxp67_ASAP7_75t_L g1522 ( 
.A(n_1494),
.Y(n_1522)
);

NOR2xp67_ASAP7_75t_L g1523 ( 
.A(n_1405),
.B(n_866),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1465),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1478),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_SL g1526 ( 
.A(n_1466),
.B(n_867),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1495),
.B(n_1072),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1480),
.Y(n_1528)
);

A2O1A1Ixp33_ASAP7_75t_L g1529 ( 
.A1(n_1400),
.A2(n_1079),
.B(n_1088),
.C(n_1073),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1501),
.B(n_1096),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1398),
.B(n_1106),
.Y(n_1531)
);

AND2x6_ASAP7_75t_SL g1532 ( 
.A(n_1462),
.B(n_1107),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1453),
.B(n_1117),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1408),
.B(n_1119),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_SL g1535 ( 
.A(n_1491),
.B(n_1432),
.Y(n_1535)
);

AND2x2_ASAP7_75t_SL g1536 ( 
.A(n_1416),
.B(n_1120),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1413),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1414),
.B(n_1128),
.Y(n_1538)
);

INVx2_ASAP7_75t_SL g1539 ( 
.A(n_1411),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1474),
.B(n_1036),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_SL g1541 ( 
.A(n_1447),
.B(n_868),
.Y(n_1541)
);

NOR3xp33_ASAP7_75t_L g1542 ( 
.A(n_1396),
.B(n_949),
.C(n_933),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1492),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_SL g1544 ( 
.A(n_1457),
.B(n_871),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1415),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1417),
.B(n_1129),
.Y(n_1546)
);

AND2x6_ASAP7_75t_L g1547 ( 
.A(n_1463),
.B(n_1130),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1423),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1401),
.B(n_1125),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_L g1550 ( 
.A(n_1469),
.B(n_1080),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1505),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_SL g1552 ( 
.A(n_1442),
.B(n_874),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1424),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_L g1554 ( 
.A(n_1472),
.B(n_1131),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1434),
.B(n_1132),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1440),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1471),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1486),
.B(n_1137),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1497),
.B(n_1141),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_1479),
.B(n_875),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1498),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_1431),
.B(n_1145),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_SL g1563 ( 
.A(n_1426),
.B(n_931),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1500),
.B(n_1143),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_SL g1565 ( 
.A(n_1441),
.B(n_877),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_SL g1566 ( 
.A(n_1506),
.B(n_879),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1467),
.A2(n_1155),
.B1(n_1159),
.B2(n_1148),
.Y(n_1567)
);

INVx2_ASAP7_75t_SL g1568 ( 
.A(n_1411),
.Y(n_1568)
);

NOR2xp67_ASAP7_75t_L g1569 ( 
.A(n_1444),
.B(n_881),
.Y(n_1569)
);

BUFx12f_ASAP7_75t_L g1570 ( 
.A(n_1406),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1403),
.B(n_1125),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1481),
.B(n_962),
.Y(n_1572)
);

INVxp67_ASAP7_75t_SL g1573 ( 
.A(n_1438),
.Y(n_1573)
);

INVx2_ASAP7_75t_SL g1574 ( 
.A(n_1435),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1420),
.Y(n_1575)
);

INVx6_ASAP7_75t_L g1576 ( 
.A(n_1488),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1439),
.B(n_1163),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1421),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1427),
.B(n_1147),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_SL g1580 ( 
.A(n_1456),
.B(n_882),
.Y(n_1580)
);

INVxp67_ASAP7_75t_L g1581 ( 
.A(n_1428),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_SL g1582 ( 
.A(n_1454),
.B(n_885),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1487),
.B(n_965),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1429),
.Y(n_1584)
);

NAND2xp33_ASAP7_75t_SL g1585 ( 
.A(n_1452),
.B(n_888),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1499),
.B(n_1170),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1437),
.Y(n_1587)
);

INVx4_ASAP7_75t_L g1588 ( 
.A(n_1488),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1448),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1449),
.Y(n_1590)
);

AOI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1482),
.A2(n_1182),
.B1(n_1183),
.B2(n_1171),
.Y(n_1591)
);

A2O1A1Ixp33_ASAP7_75t_L g1592 ( 
.A1(n_1496),
.A2(n_1188),
.B(n_1191),
.C(n_1187),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1485),
.B(n_985),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1422),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1473),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1430),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1508),
.A2(n_1502),
.B1(n_1407),
.B2(n_1446),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1412),
.B(n_1199),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1435),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1418),
.B(n_1201),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1503),
.B(n_1206),
.Y(n_1601)
);

O2A1O1Ixp33_ASAP7_75t_L g1602 ( 
.A1(n_1450),
.A2(n_1210),
.B(n_893),
.C(n_895),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1407),
.B(n_892),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_R g1604 ( 
.A(n_1468),
.B(n_896),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1407),
.B(n_897),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1502),
.B(n_898),
.Y(n_1606)
);

INVx2_ASAP7_75t_SL g1607 ( 
.A(n_1509),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1455),
.B(n_907),
.Y(n_1608)
);

NAND3xp33_ASAP7_75t_L g1609 ( 
.A(n_1433),
.B(n_1489),
.C(n_1464),
.Y(n_1609)
);

NAND2xp33_ASAP7_75t_SL g1610 ( 
.A(n_1493),
.B(n_909),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1410),
.B(n_1147),
.Y(n_1611)
);

O2A1O1Ixp33_ASAP7_75t_L g1612 ( 
.A1(n_1458),
.A2(n_1459),
.B(n_1460),
.C(n_1410),
.Y(n_1612)
);

INVx1_ASAP7_75t_SL g1613 ( 
.A(n_1399),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1502),
.B(n_910),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1409),
.B(n_911),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1451),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_SL g1617 ( 
.A(n_1425),
.B(n_913),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_SL g1618 ( 
.A(n_1451),
.B(n_914),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1443),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_SL g1620 ( 
.A(n_1476),
.B(n_917),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_SL g1621 ( 
.A(n_1477),
.B(n_922),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1504),
.B(n_923),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1445),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1464),
.B(n_1000),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1436),
.B(n_925),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_SL g1626 ( 
.A(n_1462),
.B(n_928),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1436),
.B(n_930),
.Y(n_1627)
);

BUFx5_ASAP7_75t_L g1628 ( 
.A(n_1406),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1397),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1490),
.B(n_935),
.Y(n_1630)
);

O2A1O1Ixp33_ASAP7_75t_L g1631 ( 
.A1(n_1398),
.A2(n_938),
.B(n_940),
.C(n_936),
.Y(n_1631)
);

NAND2xp33_ASAP7_75t_R g1632 ( 
.A(n_1470),
.B(n_941),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1404),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1490),
.B(n_942),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1397),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1490),
.B(n_944),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1397),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1404),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1397),
.Y(n_1639)
);

BUFx6f_ASAP7_75t_SL g1640 ( 
.A(n_1406),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1490),
.B(n_945),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1484),
.B(n_1016),
.Y(n_1642)
);

INVx2_ASAP7_75t_SL g1643 ( 
.A(n_1466),
.Y(n_1643)
);

INVxp67_ASAP7_75t_SL g1644 ( 
.A(n_1453),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1490),
.B(n_946),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1466),
.B(n_947),
.Y(n_1646)
);

INVx3_ASAP7_75t_L g1647 ( 
.A(n_1411),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1490),
.B(n_952),
.Y(n_1648)
);

INVx4_ASAP7_75t_L g1649 ( 
.A(n_1488),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1404),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1397),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1404),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1490),
.B(n_955),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1445),
.B(n_1021),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1490),
.B(n_956),
.Y(n_1655)
);

INVx4_ASAP7_75t_L g1656 ( 
.A(n_1488),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1404),
.Y(n_1657)
);

AOI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1461),
.A2(n_958),
.B1(n_960),
.B2(n_957),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1490),
.B(n_967),
.Y(n_1659)
);

INVxp67_ASAP7_75t_L g1660 ( 
.A(n_1494),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_SL g1661 ( 
.A(n_1466),
.B(n_972),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1491),
.B(n_1205),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1404),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1397),
.Y(n_1664)
);

INVx2_ASAP7_75t_SL g1665 ( 
.A(n_1466),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1490),
.B(n_973),
.Y(n_1666)
);

INVx2_ASAP7_75t_SL g1667 ( 
.A(n_1466),
.Y(n_1667)
);

INVxp67_ASAP7_75t_L g1668 ( 
.A(n_1494),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1510),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1511),
.Y(n_1670)
);

AOI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1644),
.A2(n_1091),
.B(n_1057),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1515),
.B(n_979),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1623),
.B(n_1643),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1516),
.B(n_980),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1518),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_SL g1676 ( 
.A(n_1536),
.B(n_961),
.Y(n_1676)
);

AOI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1562),
.A2(n_1208),
.B1(n_986),
.B2(n_993),
.Y(n_1677)
);

OR2x6_ASAP7_75t_L g1678 ( 
.A(n_1570),
.B(n_1091),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1581),
.B(n_1550),
.Y(n_1679)
);

AND2x2_ASAP7_75t_SL g1680 ( 
.A(n_1540),
.B(n_1091),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1537),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1545),
.Y(n_1682)
);

BUFx6f_ASAP7_75t_L g1683 ( 
.A(n_1576),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1630),
.B(n_991),
.Y(n_1684)
);

NOR3xp33_ASAP7_75t_SL g1685 ( 
.A(n_1632),
.B(n_1031),
.C(n_1030),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1548),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1553),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1634),
.B(n_996),
.Y(n_1688)
);

NOR2x2_ASAP7_75t_L g1689 ( 
.A(n_1556),
.B(n_1619),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1557),
.Y(n_1690)
);

BUFx8_ASAP7_75t_L g1691 ( 
.A(n_1640),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_L g1692 ( 
.A(n_1554),
.B(n_1038),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1572),
.A2(n_983),
.B1(n_1028),
.B2(n_995),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1561),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1633),
.Y(n_1695)
);

OR2x4_ASAP7_75t_L g1696 ( 
.A(n_1583),
.B(n_1126),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1665),
.B(n_267),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_SL g1698 ( 
.A(n_1522),
.B(n_961),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1638),
.Y(n_1699)
);

CKINVDCx20_ASAP7_75t_R g1700 ( 
.A(n_1604),
.Y(n_1700)
);

INVx1_ASAP7_75t_SL g1701 ( 
.A(n_1596),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1636),
.B(n_998),
.Y(n_1702)
);

AND2x4_ASAP7_75t_L g1703 ( 
.A(n_1667),
.B(n_268),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1513),
.Y(n_1704)
);

INVx5_ASAP7_75t_L g1705 ( 
.A(n_1576),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1650),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1652),
.Y(n_1707)
);

INVx2_ASAP7_75t_SL g1708 ( 
.A(n_1599),
.Y(n_1708)
);

NAND2x1p5_ASAP7_75t_L g1709 ( 
.A(n_1588),
.B(n_1126),
.Y(n_1709)
);

BUFx12f_ASAP7_75t_SL g1710 ( 
.A(n_1649),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1641),
.B(n_999),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_1532),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_L g1713 ( 
.A(n_1514),
.B(n_1043),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1657),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1520),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1645),
.B(n_1001),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1648),
.B(n_1002),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1524),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1525),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1653),
.B(n_1003),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_1624),
.Y(n_1721)
);

BUFx6f_ASAP7_75t_L g1722 ( 
.A(n_1656),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1660),
.B(n_1668),
.Y(n_1723)
);

BUFx4f_ASAP7_75t_L g1724 ( 
.A(n_1547),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1663),
.Y(n_1725)
);

BUFx6f_ASAP7_75t_L g1726 ( 
.A(n_1539),
.Y(n_1726)
);

AND2x4_ASAP7_75t_L g1727 ( 
.A(n_1594),
.B(n_270),
.Y(n_1727)
);

A2O1A1Ixp33_ASAP7_75t_L g1728 ( 
.A1(n_1593),
.A2(n_1180),
.B(n_1181),
.C(n_1177),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1528),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1589),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1549),
.B(n_1153),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1542),
.A2(n_995),
.B1(n_1028),
.B2(n_983),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1595),
.B(n_271),
.Y(n_1733)
);

BUFx3_ASAP7_75t_L g1734 ( 
.A(n_1647),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1568),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1543),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1575),
.Y(n_1737)
);

INVx2_ASAP7_75t_SL g1738 ( 
.A(n_1574),
.Y(n_1738)
);

OR2x2_ASAP7_75t_SL g1739 ( 
.A(n_1609),
.B(n_1153),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1584),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1551),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1662),
.B(n_1056),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1535),
.B(n_1065),
.Y(n_1743)
);

BUFx3_ASAP7_75t_L g1744 ( 
.A(n_1628),
.Y(n_1744)
);

AND2x4_ASAP7_75t_L g1745 ( 
.A(n_1607),
.B(n_272),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1655),
.B(n_1005),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_1628),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_SL g1748 ( 
.A(n_1659),
.B(n_1203),
.Y(n_1748)
);

INVx3_ASAP7_75t_L g1749 ( 
.A(n_1616),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1666),
.B(n_1008),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_SL g1751 ( 
.A(n_1628),
.B(n_1203),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1573),
.B(n_1011),
.Y(n_1752)
);

AND2x6_ASAP7_75t_SL g1753 ( 
.A(n_1654),
.B(n_1071),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1571),
.B(n_1642),
.Y(n_1754)
);

INVxp67_ASAP7_75t_L g1755 ( 
.A(n_1579),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1519),
.B(n_1012),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1578),
.Y(n_1757)
);

INVx3_ASAP7_75t_L g1758 ( 
.A(n_1613),
.Y(n_1758)
);

BUFx6f_ASAP7_75t_L g1759 ( 
.A(n_1587),
.Y(n_1759)
);

NAND2xp33_ASAP7_75t_SL g1760 ( 
.A(n_1560),
.B(n_1017),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_SL g1761 ( 
.A(n_1628),
.B(n_1018),
.Y(n_1761)
);

AOI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1541),
.A2(n_1169),
.B1(n_1184),
.B2(n_1166),
.Y(n_1762)
);

NOR2x2_ASAP7_75t_L g1763 ( 
.A(n_1629),
.B(n_1076),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1521),
.B(n_1527),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1635),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1637),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_SL g1767 ( 
.A(n_1658),
.B(n_1022),
.Y(n_1767)
);

AOI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1580),
.A2(n_1194),
.B1(n_1197),
.B2(n_1190),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_SL g1769 ( 
.A(n_1512),
.B(n_1026),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_1610),
.Y(n_1770)
);

HB1xp67_ASAP7_75t_L g1771 ( 
.A(n_1590),
.Y(n_1771)
);

A2O1A1Ixp33_ASAP7_75t_L g1772 ( 
.A1(n_1529),
.A2(n_1200),
.B(n_1198),
.C(n_1032),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_SL g1773 ( 
.A(n_1597),
.B(n_1027),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_L g1774 ( 
.A(n_1664),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1530),
.B(n_1034),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1639),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1651),
.Y(n_1777)
);

INVx1_ASAP7_75t_SL g1778 ( 
.A(n_1611),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_SL g1779 ( 
.A(n_1569),
.B(n_1037),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1531),
.B(n_1042),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1523),
.B(n_1089),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1517),
.B(n_1046),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_SL g1783 ( 
.A(n_1612),
.B(n_1048),
.Y(n_1783)
);

BUFx6f_ASAP7_75t_L g1784 ( 
.A(n_1547),
.Y(n_1784)
);

AND2x4_ASAP7_75t_L g1785 ( 
.A(n_1552),
.B(n_274),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1534),
.B(n_1049),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1669),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1681),
.Y(n_1788)
);

INVxp67_ASAP7_75t_L g1789 ( 
.A(n_1675),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1682),
.Y(n_1790)
);

INVx4_ASAP7_75t_L g1791 ( 
.A(n_1705),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_SL g1792 ( 
.A1(n_1680),
.A2(n_1563),
.B1(n_1625),
.B2(n_1601),
.Y(n_1792)
);

AND3x1_ASAP7_75t_SL g1793 ( 
.A(n_1686),
.B(n_1097),
.C(n_1092),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1687),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_SL g1795 ( 
.A(n_1721),
.B(n_1615),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1690),
.Y(n_1796)
);

INVx4_ASAP7_75t_L g1797 ( 
.A(n_1705),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_SL g1798 ( 
.A(n_1754),
.B(n_1622),
.Y(n_1798)
);

AOI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1692),
.A2(n_1585),
.B1(n_1626),
.B2(n_1526),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1694),
.Y(n_1800)
);

NOR2xp33_ASAP7_75t_L g1801 ( 
.A(n_1679),
.B(n_1646),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1695),
.Y(n_1802)
);

OR2x6_ASAP7_75t_L g1803 ( 
.A(n_1683),
.B(n_1627),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1764),
.B(n_1538),
.Y(n_1804)
);

BUFx6f_ASAP7_75t_L g1805 ( 
.A(n_1683),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1699),
.Y(n_1806)
);

HB1xp67_ASAP7_75t_L g1807 ( 
.A(n_1701),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1713),
.B(n_1546),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1706),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1707),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1714),
.B(n_1725),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1730),
.B(n_1555),
.Y(n_1812)
);

BUFx3_ASAP7_75t_L g1813 ( 
.A(n_1722),
.Y(n_1813)
);

NOR2xp33_ASAP7_75t_L g1814 ( 
.A(n_1755),
.B(n_1661),
.Y(n_1814)
);

BUFx6f_ASAP7_75t_L g1815 ( 
.A(n_1722),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1731),
.B(n_1558),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1737),
.Y(n_1817)
);

NAND3xp33_ASAP7_75t_L g1818 ( 
.A(n_1677),
.B(n_1591),
.C(n_1592),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1672),
.B(n_1559),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_SL g1820 ( 
.A(n_1758),
.B(n_1759),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1740),
.Y(n_1821)
);

INVx4_ASAP7_75t_L g1822 ( 
.A(n_1726),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1670),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1774),
.Y(n_1824)
);

INVx3_ASAP7_75t_L g1825 ( 
.A(n_1734),
.Y(n_1825)
);

CKINVDCx5p33_ASAP7_75t_R g1826 ( 
.A(n_1700),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_L g1827 ( 
.A(n_1743),
.B(n_1676),
.Y(n_1827)
);

AOI22x1_ASAP7_75t_L g1828 ( 
.A1(n_1671),
.A2(n_1631),
.B1(n_1547),
.B2(n_1602),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1674),
.B(n_1564),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1741),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1778),
.B(n_1566),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1704),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1781),
.B(n_1577),
.Y(n_1833)
);

BUFx2_ASAP7_75t_L g1834 ( 
.A(n_1689),
.Y(n_1834)
);

INVxp67_ASAP7_75t_SL g1835 ( 
.A(n_1771),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1715),
.Y(n_1836)
);

INVx5_ASAP7_75t_L g1837 ( 
.A(n_1726),
.Y(n_1837)
);

INVxp67_ASAP7_75t_SL g1838 ( 
.A(n_1735),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_L g1839 ( 
.A(n_1742),
.B(n_1582),
.Y(n_1839)
);

BUFx6f_ASAP7_75t_L g1840 ( 
.A(n_1708),
.Y(n_1840)
);

BUFx2_ASAP7_75t_L g1841 ( 
.A(n_1673),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1718),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1684),
.B(n_1533),
.Y(n_1843)
);

BUFx2_ASAP7_75t_L g1844 ( 
.A(n_1710),
.Y(n_1844)
);

AOI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1785),
.A2(n_1544),
.B1(n_1618),
.B2(n_1617),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1757),
.Y(n_1846)
);

INVx4_ASAP7_75t_L g1847 ( 
.A(n_1747),
.Y(n_1847)
);

INVxp67_ASAP7_75t_L g1848 ( 
.A(n_1723),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1766),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_L g1850 ( 
.A(n_1696),
.B(n_1565),
.Y(n_1850)
);

NAND3xp33_ASAP7_75t_L g1851 ( 
.A(n_1693),
.B(n_1685),
.C(n_1732),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_SL g1852 ( 
.A(n_1759),
.B(n_1770),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1776),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1688),
.B(n_1702),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1719),
.Y(n_1855)
);

BUFx4f_ASAP7_75t_L g1856 ( 
.A(n_1784),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1711),
.B(n_1586),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1729),
.B(n_1603),
.Y(n_1858)
);

BUFx4f_ASAP7_75t_L g1859 ( 
.A(n_1784),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1736),
.Y(n_1860)
);

INVx1_ASAP7_75t_SL g1861 ( 
.A(n_1763),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1716),
.B(n_1608),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1717),
.B(n_1620),
.Y(n_1863)
);

BUFx6f_ASAP7_75t_L g1864 ( 
.A(n_1738),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1777),
.Y(n_1865)
);

AOI22xp5_ASAP7_75t_L g1866 ( 
.A1(n_1748),
.A2(n_1621),
.B1(n_1606),
.B2(n_1614),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1765),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1749),
.Y(n_1868)
);

OR2x6_ASAP7_75t_L g1869 ( 
.A(n_1744),
.B(n_1605),
.Y(n_1869)
);

INVx3_ASAP7_75t_L g1870 ( 
.A(n_1691),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1727),
.B(n_1600),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1733),
.Y(n_1872)
);

BUFx3_ASAP7_75t_L g1873 ( 
.A(n_1697),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1720),
.B(n_1567),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1703),
.Y(n_1875)
);

BUFx2_ASAP7_75t_L g1876 ( 
.A(n_1745),
.Y(n_1876)
);

INVxp67_ASAP7_75t_L g1877 ( 
.A(n_1678),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1698),
.B(n_1598),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1782),
.B(n_1100),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1746),
.B(n_1050),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_1753),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1752),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1750),
.B(n_1051),
.Y(n_1883)
);

OAI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1756),
.A2(n_1062),
.B1(n_1064),
.B2(n_1053),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1775),
.B(n_1068),
.Y(n_1885)
);

HB1xp67_ASAP7_75t_L g1886 ( 
.A(n_1739),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1786),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_L g1888 ( 
.A1(n_1773),
.A2(n_995),
.B1(n_1028),
.B2(n_983),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1780),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_SL g1890 ( 
.A(n_1724),
.B(n_1069),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1751),
.B(n_1105),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1769),
.B(n_1127),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1783),
.Y(n_1893)
);

AND2x4_ASAP7_75t_L g1894 ( 
.A(n_1678),
.B(n_276),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1761),
.Y(n_1895)
);

INVx1_ASAP7_75t_SL g1896 ( 
.A(n_1712),
.Y(n_1896)
);

BUFx2_ASAP7_75t_L g1897 ( 
.A(n_1760),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1709),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1779),
.Y(n_1899)
);

AOI22xp33_ASAP7_75t_L g1900 ( 
.A1(n_1767),
.A2(n_1028),
.B1(n_995),
.B2(n_1070),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1762),
.Y(n_1901)
);

INVx3_ASAP7_75t_L g1902 ( 
.A(n_1728),
.Y(n_1902)
);

BUFx6f_ASAP7_75t_L g1903 ( 
.A(n_1772),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1768),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1754),
.B(n_1078),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1669),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1669),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1669),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1669),
.Y(n_1909)
);

INVxp33_ASAP7_75t_L g1910 ( 
.A(n_1675),
.Y(n_1910)
);

AOI22xp5_ASAP7_75t_L g1911 ( 
.A1(n_1692),
.A2(n_1164),
.B1(n_1161),
.B2(n_1084),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1669),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1754),
.B(n_1083),
.Y(n_1913)
);

BUFx6f_ASAP7_75t_L g1914 ( 
.A(n_1705),
.Y(n_1914)
);

AOI211x1_ASAP7_75t_L g1915 ( 
.A1(n_1811),
.A2(n_1154),
.B(n_1162),
.C(n_1142),
.Y(n_1915)
);

OAI21x1_ASAP7_75t_L g1916 ( 
.A1(n_1828),
.A2(n_1028),
.B(n_995),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1807),
.B(n_1165),
.Y(n_1917)
);

NOR2xp33_ASAP7_75t_L g1918 ( 
.A(n_1827),
.B(n_1087),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1787),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1796),
.Y(n_1920)
);

AOI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1804),
.A2(n_1133),
.B(n_1126),
.Y(n_1921)
);

AOI22xp33_ASAP7_75t_L g1922 ( 
.A1(n_1892),
.A2(n_1168),
.B1(n_1173),
.B2(n_1172),
.Y(n_1922)
);

NOR2xp67_ASAP7_75t_L g1923 ( 
.A(n_1848),
.B(n_278),
.Y(n_1923)
);

AOI21xp5_ASAP7_75t_L g1924 ( 
.A1(n_1854),
.A2(n_1207),
.B(n_1133),
.Y(n_1924)
);

BUFx2_ASAP7_75t_L g1925 ( 
.A(n_1834),
.Y(n_1925)
);

AO21x2_ASAP7_75t_L g1926 ( 
.A1(n_1893),
.A2(n_1099),
.B(n_1094),
.Y(n_1926)
);

AOI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1843),
.A2(n_1829),
.B(n_1819),
.Y(n_1927)
);

AO31x2_ASAP7_75t_L g1928 ( 
.A1(n_1850),
.A2(n_1207),
.A3(n_1133),
.B(n_280),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1808),
.B(n_1175),
.Y(n_1929)
);

INVx3_ASAP7_75t_L g1930 ( 
.A(n_1791),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1889),
.B(n_1176),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1816),
.B(n_1102),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1879),
.B(n_1103),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1887),
.B(n_1109),
.Y(n_1934)
);

AO31x2_ASAP7_75t_L g1935 ( 
.A1(n_1862),
.A2(n_1207),
.A3(n_283),
.B(n_284),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1800),
.Y(n_1936)
);

BUFx2_ASAP7_75t_L g1937 ( 
.A(n_1841),
.Y(n_1937)
);

OAI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1833),
.A2(n_1818),
.B(n_1857),
.Y(n_1938)
);

OA21x2_ASAP7_75t_L g1939 ( 
.A1(n_1888),
.A2(n_1112),
.B(n_1110),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1882),
.B(n_1115),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1802),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1801),
.B(n_1118),
.Y(n_1942)
);

OAI21xp5_ASAP7_75t_SL g1943 ( 
.A1(n_1792),
.A2(n_1799),
.B(n_1839),
.Y(n_1943)
);

BUFx3_ASAP7_75t_L g1944 ( 
.A(n_1914),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1871),
.B(n_1122),
.Y(n_1945)
);

O2A1O1Ixp5_ASAP7_75t_L g1946 ( 
.A1(n_1902),
.A2(n_1124),
.B(n_1138),
.C(n_1123),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1812),
.B(n_1144),
.Y(n_1947)
);

OAI21xp5_ASAP7_75t_L g1948 ( 
.A1(n_1874),
.A2(n_1150),
.B(n_1146),
.Y(n_1948)
);

OAI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1851),
.A2(n_1152),
.B(n_1151),
.Y(n_1949)
);

OAI21xp33_ASAP7_75t_L g1950 ( 
.A1(n_1911),
.A2(n_1158),
.B(n_1156),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1824),
.B(n_1160),
.Y(n_1951)
);

OAI21x1_ASAP7_75t_L g1952 ( 
.A1(n_1895),
.A2(n_286),
.B(n_279),
.Y(n_1952)
);

OAI21x1_ASAP7_75t_L g1953 ( 
.A1(n_1866),
.A2(n_289),
.B(n_287),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1835),
.B(n_1),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1878),
.B(n_1),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1872),
.B(n_2),
.Y(n_1956)
);

BUFx6f_ASAP7_75t_L g1957 ( 
.A(n_1914),
.Y(n_1957)
);

INVx5_ASAP7_75t_L g1958 ( 
.A(n_1815),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1863),
.B(n_2),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1831),
.B(n_3),
.Y(n_1960)
);

INVx2_ASAP7_75t_SL g1961 ( 
.A(n_1837),
.Y(n_1961)
);

OAI21x1_ASAP7_75t_L g1962 ( 
.A1(n_1830),
.A2(n_291),
.B(n_290),
.Y(n_1962)
);

O2A1O1Ixp5_ASAP7_75t_L g1963 ( 
.A1(n_1798),
.A2(n_6),
.B(n_4),
.C(n_5),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1806),
.Y(n_1964)
);

A2O1A1Ixp33_ASAP7_75t_L g1965 ( 
.A1(n_1845),
.A2(n_6),
.B(n_4),
.C(n_5),
.Y(n_1965)
);

OA21x2_ASAP7_75t_L g1966 ( 
.A1(n_1900),
.A2(n_294),
.B(n_293),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1905),
.B(n_7),
.Y(n_1967)
);

OAI21x1_ASAP7_75t_L g1968 ( 
.A1(n_1846),
.A2(n_296),
.B(n_295),
.Y(n_1968)
);

INVx3_ASAP7_75t_L g1969 ( 
.A(n_1797),
.Y(n_1969)
);

OAI22xp5_ASAP7_75t_L g1970 ( 
.A1(n_1838),
.A2(n_1814),
.B1(n_1875),
.B2(n_1876),
.Y(n_1970)
);

OAI21x1_ASAP7_75t_L g1971 ( 
.A1(n_1849),
.A2(n_300),
.B(n_299),
.Y(n_1971)
);

BUFx6f_ASAP7_75t_L g1972 ( 
.A(n_1815),
.Y(n_1972)
);

AOI221x1_ASAP7_75t_L g1973 ( 
.A1(n_1904),
.A2(n_11),
.B1(n_8),
.B2(n_10),
.C(n_12),
.Y(n_1973)
);

AO31x2_ASAP7_75t_L g1974 ( 
.A1(n_1901),
.A2(n_302),
.A3(n_303),
.B(n_301),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1913),
.B(n_8),
.Y(n_1975)
);

INVx1_ASAP7_75t_SL g1976 ( 
.A(n_1837),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1880),
.B(n_10),
.Y(n_1977)
);

AOI21x1_ASAP7_75t_L g1978 ( 
.A1(n_1897),
.A2(n_305),
.B(n_304),
.Y(n_1978)
);

AOI221xp5_ASAP7_75t_L g1979 ( 
.A1(n_1886),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.C(n_16),
.Y(n_1979)
);

A2O1A1Ixp33_ASAP7_75t_L g1980 ( 
.A1(n_1899),
.A2(n_1883),
.B(n_1885),
.C(n_1858),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1909),
.Y(n_1981)
);

AO21x2_ASAP7_75t_L g1982 ( 
.A1(n_1817),
.A2(n_310),
.B(n_309),
.Y(n_1982)
);

AO31x2_ASAP7_75t_L g1983 ( 
.A1(n_1788),
.A2(n_313),
.A3(n_314),
.B(n_312),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1912),
.B(n_1795),
.Y(n_1984)
);

NOR3xp33_ASAP7_75t_L g1985 ( 
.A(n_1890),
.B(n_13),
.C(n_14),
.Y(n_1985)
);

A2O1A1Ixp33_ASAP7_75t_L g1986 ( 
.A1(n_1903),
.A2(n_17),
.B(n_15),
.C(n_16),
.Y(n_1986)
);

A2O1A1Ixp33_ASAP7_75t_L g1987 ( 
.A1(n_1903),
.A2(n_20),
.B(n_17),
.C(n_18),
.Y(n_1987)
);

OAI21x1_ASAP7_75t_L g1988 ( 
.A1(n_1853),
.A2(n_317),
.B(n_315),
.Y(n_1988)
);

INVx3_ASAP7_75t_L g1989 ( 
.A(n_1840),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1823),
.B(n_18),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1832),
.B(n_1836),
.Y(n_1991)
);

OAI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1789),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_1992)
);

NAND2x1p5_ASAP7_75t_L g1993 ( 
.A(n_1822),
.B(n_320),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1790),
.Y(n_1994)
);

OAI21xp5_ASAP7_75t_L g1995 ( 
.A1(n_1884),
.A2(n_1891),
.B(n_1820),
.Y(n_1995)
);

HB1xp67_ASAP7_75t_L g1996 ( 
.A(n_1984),
.Y(n_1996)
);

CKINVDCx5p33_ASAP7_75t_R g1997 ( 
.A(n_1944),
.Y(n_1997)
);

BUFx3_ASAP7_75t_L g1998 ( 
.A(n_1958),
.Y(n_1998)
);

HB1xp67_ASAP7_75t_L g1999 ( 
.A(n_1970),
.Y(n_1999)
);

AND2x6_ASAP7_75t_L g2000 ( 
.A(n_1994),
.B(n_1894),
.Y(n_2000)
);

HB1xp67_ASAP7_75t_L g2001 ( 
.A(n_1920),
.Y(n_2001)
);

INVx4_ASAP7_75t_L g2002 ( 
.A(n_1958),
.Y(n_2002)
);

AND2x4_ASAP7_75t_L g2003 ( 
.A(n_1937),
.B(n_1989),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1941),
.Y(n_2004)
);

BUFx6f_ASAP7_75t_L g2005 ( 
.A(n_1972),
.Y(n_2005)
);

AND2x4_ASAP7_75t_L g2006 ( 
.A(n_1961),
.B(n_1847),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1990),
.B(n_1821),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1981),
.Y(n_2008)
);

OR2x2_ASAP7_75t_L g2009 ( 
.A(n_1955),
.B(n_1794),
.Y(n_2009)
);

HB1xp67_ASAP7_75t_L g2010 ( 
.A(n_1919),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1991),
.B(n_1809),
.Y(n_2011)
);

OR2x2_ASAP7_75t_L g2012 ( 
.A(n_1959),
.B(n_1810),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1936),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1964),
.Y(n_2014)
);

INVx3_ASAP7_75t_L g2015 ( 
.A(n_1972),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1916),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1928),
.Y(n_2017)
);

CKINVDCx6p67_ASAP7_75t_R g2018 ( 
.A(n_1957),
.Y(n_2018)
);

AOI22xp33_ASAP7_75t_SL g2019 ( 
.A1(n_1918),
.A2(n_1861),
.B1(n_1881),
.B2(n_1873),
.Y(n_2019)
);

BUFx2_ASAP7_75t_L g2020 ( 
.A(n_1925),
.Y(n_2020)
);

O2A1O1Ixp5_ASAP7_75t_L g2021 ( 
.A1(n_1965),
.A2(n_1852),
.B(n_1865),
.C(n_1906),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1932),
.B(n_1945),
.Y(n_2022)
);

INVx5_ASAP7_75t_L g2023 ( 
.A(n_1957),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1956),
.B(n_1907),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1938),
.B(n_1908),
.Y(n_2025)
);

INVxp67_ASAP7_75t_SL g2026 ( 
.A(n_1927),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1928),
.Y(n_2027)
);

BUFx2_ASAP7_75t_L g2028 ( 
.A(n_1976),
.Y(n_2028)
);

OR2x2_ASAP7_75t_L g2029 ( 
.A(n_1954),
.B(n_1910),
.Y(n_2029)
);

AND2x4_ASAP7_75t_L g2030 ( 
.A(n_1930),
.B(n_1813),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1980),
.B(n_1842),
.Y(n_2031)
);

INVx2_ASAP7_75t_SL g2032 ( 
.A(n_1969),
.Y(n_2032)
);

BUFx6f_ASAP7_75t_L g2033 ( 
.A(n_1917),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1943),
.B(n_1855),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1935),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1929),
.B(n_1860),
.Y(n_2036)
);

AND2x4_ASAP7_75t_L g2037 ( 
.A(n_1923),
.B(n_1844),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1942),
.B(n_1867),
.Y(n_2038)
);

A2O1A1Ixp33_ASAP7_75t_SL g2039 ( 
.A1(n_1985),
.A2(n_1877),
.B(n_1898),
.C(n_1870),
.Y(n_2039)
);

AOI21xp5_ASAP7_75t_L g2040 ( 
.A1(n_1946),
.A2(n_1869),
.B(n_1859),
.Y(n_2040)
);

BUFx4_ASAP7_75t_SL g2041 ( 
.A(n_1986),
.Y(n_2041)
);

AOI21xp5_ASAP7_75t_L g2042 ( 
.A1(n_1924),
.A2(n_1869),
.B(n_1856),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1977),
.B(n_1826),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1996),
.B(n_1951),
.Y(n_2044)
);

BUFx2_ASAP7_75t_L g2045 ( 
.A(n_2020),
.Y(n_2045)
);

OAI22xp5_ASAP7_75t_L g2046 ( 
.A1(n_2034),
.A2(n_1960),
.B1(n_1987),
.B2(n_1979),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_2001),
.Y(n_2047)
);

OR2x2_ASAP7_75t_L g2048 ( 
.A(n_2009),
.B(n_1967),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_2007),
.B(n_1995),
.Y(n_2049)
);

BUFx3_ASAP7_75t_L g2050 ( 
.A(n_2005),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_2025),
.B(n_1975),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_2010),
.B(n_1915),
.Y(n_2052)
);

BUFx3_ASAP7_75t_L g2053 ( 
.A(n_2005),
.Y(n_2053)
);

A2O1A1Ixp33_ASAP7_75t_L g2054 ( 
.A1(n_2021),
.A2(n_1963),
.B(n_1953),
.C(n_1949),
.Y(n_2054)
);

AND2x4_ASAP7_75t_L g2055 ( 
.A(n_2003),
.B(n_1935),
.Y(n_2055)
);

NOR2xp33_ASAP7_75t_L g2056 ( 
.A(n_2043),
.B(n_1896),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_2024),
.B(n_1983),
.Y(n_2057)
);

A2O1A1Ixp33_ASAP7_75t_L g2058 ( 
.A1(n_2026),
.A2(n_1948),
.B(n_1950),
.C(n_1921),
.Y(n_2058)
);

O2A1O1Ixp33_ASAP7_75t_L g2059 ( 
.A1(n_2039),
.A2(n_1992),
.B(n_1931),
.C(n_1940),
.Y(n_2059)
);

BUFx3_ASAP7_75t_L g2060 ( 
.A(n_2030),
.Y(n_2060)
);

AOI21xp5_ASAP7_75t_SL g2061 ( 
.A1(n_2040),
.A2(n_1973),
.B(n_1993),
.Y(n_2061)
);

AOI21xp5_ASAP7_75t_L g2062 ( 
.A1(n_2031),
.A2(n_1966),
.B(n_1926),
.Y(n_2062)
);

NOR2xp33_ASAP7_75t_L g2063 ( 
.A(n_2033),
.B(n_1933),
.Y(n_2063)
);

AND2x4_ASAP7_75t_L g2064 ( 
.A(n_2011),
.B(n_1983),
.Y(n_2064)
);

AND2x4_ASAP7_75t_L g2065 ( 
.A(n_2028),
.B(n_1974),
.Y(n_2065)
);

AOI21x1_ASAP7_75t_SL g2066 ( 
.A1(n_2037),
.A2(n_1934),
.B(n_1947),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_2022),
.B(n_1999),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_2004),
.Y(n_2068)
);

A2O1A1Ixp33_ASAP7_75t_L g2069 ( 
.A1(n_2042),
.A2(n_1922),
.B(n_1988),
.C(n_1968),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_2008),
.B(n_1982),
.Y(n_2070)
);

INVxp67_ASAP7_75t_L g2071 ( 
.A(n_2029),
.Y(n_2071)
);

AND2x2_ASAP7_75t_SL g2072 ( 
.A(n_2002),
.B(n_1939),
.Y(n_2072)
);

OA21x2_ASAP7_75t_L g2073 ( 
.A1(n_2017),
.A2(n_1971),
.B(n_1962),
.Y(n_2073)
);

A2O1A1Ixp33_ASAP7_75t_L g2074 ( 
.A1(n_2041),
.A2(n_1952),
.B(n_1793),
.C(n_1868),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_SL g2075 ( 
.A(n_2012),
.B(n_1978),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_2013),
.B(n_1974),
.Y(n_2076)
);

AND2x4_ASAP7_75t_L g2077 ( 
.A(n_2014),
.B(n_1840),
.Y(n_2077)
);

O2A1O1Ixp33_ASAP7_75t_L g2078 ( 
.A1(n_2038),
.A2(n_1803),
.B(n_1825),
.C(n_24),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_2033),
.B(n_1803),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_2036),
.B(n_1864),
.Y(n_2080)
);

O2A1O1Ixp33_ASAP7_75t_L g2081 ( 
.A1(n_2027),
.A2(n_2035),
.B(n_2032),
.C(n_1998),
.Y(n_2081)
);

CKINVDCx5p33_ASAP7_75t_R g2082 ( 
.A(n_1997),
.Y(n_2082)
);

AOI21xp5_ASAP7_75t_L g2083 ( 
.A1(n_2016),
.A2(n_1864),
.B(n_1805),
.Y(n_2083)
);

AND2x4_ASAP7_75t_L g2084 ( 
.A(n_2023),
.B(n_1805),
.Y(n_2084)
);

INVx3_ASAP7_75t_L g2085 ( 
.A(n_2015),
.Y(n_2085)
);

AOI21xp5_ASAP7_75t_L g2086 ( 
.A1(n_2000),
.A2(n_323),
.B(n_322),
.Y(n_2086)
);

OAI22xp5_ASAP7_75t_SL g2087 ( 
.A1(n_2019),
.A2(n_25),
.B1(n_21),
.B2(n_23),
.Y(n_2087)
);

INVx8_ASAP7_75t_L g2088 ( 
.A(n_2023),
.Y(n_2088)
);

AND2x2_ASAP7_75t_L g2089 ( 
.A(n_2006),
.B(n_23),
.Y(n_2089)
);

NAND2x1p5_ASAP7_75t_L g2090 ( 
.A(n_2000),
.B(n_2018),
.Y(n_2090)
);

BUFx6f_ASAP7_75t_L g2091 ( 
.A(n_2000),
.Y(n_2091)
);

A2O1A1Ixp33_ASAP7_75t_L g2092 ( 
.A1(n_2021),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_2092)
);

NOR2x1_ASAP7_75t_L g2093 ( 
.A(n_2031),
.B(n_26),
.Y(n_2093)
);

HB1xp67_ASAP7_75t_L g2094 ( 
.A(n_1996),
.Y(n_2094)
);

AOI22xp33_ASAP7_75t_SL g2095 ( 
.A1(n_2046),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_2068),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_2047),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2094),
.Y(n_2098)
);

INVx3_ASAP7_75t_L g2099 ( 
.A(n_2060),
.Y(n_2099)
);

BUFx2_ASAP7_75t_L g2100 ( 
.A(n_2045),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2070),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2076),
.Y(n_2102)
);

INVx2_ASAP7_75t_SL g2103 ( 
.A(n_2088),
.Y(n_2103)
);

AOI22xp33_ASAP7_75t_SL g2104 ( 
.A1(n_2087),
.A2(n_31),
.B1(n_28),
.B2(n_30),
.Y(n_2104)
);

NOR2xp33_ASAP7_75t_L g2105 ( 
.A(n_2051),
.B(n_30),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_2064),
.Y(n_2106)
);

AND2x4_ASAP7_75t_L g2107 ( 
.A(n_2055),
.B(n_325),
.Y(n_2107)
);

OAI21x1_ASAP7_75t_L g2108 ( 
.A1(n_2062),
.A2(n_327),
.B(n_326),
.Y(n_2108)
);

NOR2xp33_ASAP7_75t_L g2109 ( 
.A(n_2071),
.B(n_32),
.Y(n_2109)
);

BUFx3_ASAP7_75t_L g2110 ( 
.A(n_2050),
.Y(n_2110)
);

INVx3_ASAP7_75t_L g2111 ( 
.A(n_2088),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2057),
.Y(n_2112)
);

OR2x2_ASAP7_75t_L g2113 ( 
.A(n_2049),
.B(n_32),
.Y(n_2113)
);

OR2x2_ASAP7_75t_L g2114 ( 
.A(n_2067),
.B(n_2048),
.Y(n_2114)
);

OAI21x1_ASAP7_75t_L g2115 ( 
.A1(n_2083),
.A2(n_330),
.B(n_329),
.Y(n_2115)
);

HB1xp67_ASAP7_75t_L g2116 ( 
.A(n_2065),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2081),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2052),
.Y(n_2118)
);

INVxp67_ASAP7_75t_L g2119 ( 
.A(n_2044),
.Y(n_2119)
);

OA21x2_ASAP7_75t_L g2120 ( 
.A1(n_2075),
.A2(n_41),
.B(n_33),
.Y(n_2120)
);

BUFx3_ASAP7_75t_L g2121 ( 
.A(n_2053),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_2079),
.B(n_33),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_2073),
.Y(n_2123)
);

BUFx3_ASAP7_75t_L g2124 ( 
.A(n_2082),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2080),
.Y(n_2125)
);

INVx1_ASAP7_75t_SL g2126 ( 
.A(n_2077),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2093),
.Y(n_2127)
);

OAI21x1_ASAP7_75t_L g2128 ( 
.A1(n_2066),
.A2(n_333),
.B(n_332),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_2085),
.Y(n_2129)
);

AO21x1_ASAP7_75t_SL g2130 ( 
.A1(n_2061),
.A2(n_34),
.B(n_35),
.Y(n_2130)
);

HB1xp67_ASAP7_75t_L g2131 ( 
.A(n_2091),
.Y(n_2131)
);

CKINVDCx5p33_ASAP7_75t_R g2132 ( 
.A(n_2084),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2072),
.Y(n_2133)
);

AND2x4_ASAP7_75t_L g2134 ( 
.A(n_2091),
.B(n_337),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2078),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2090),
.Y(n_2136)
);

OR2x6_ASAP7_75t_L g2137 ( 
.A(n_2086),
.B(n_338),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_2089),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2092),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2069),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2054),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2074),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_2063),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_2056),
.B(n_34),
.Y(n_2144)
);

INVx5_ASAP7_75t_L g2145 ( 
.A(n_2059),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2058),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2068),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2068),
.Y(n_2148)
);

OAI22xp33_ASAP7_75t_L g2149 ( 
.A1(n_2046),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2068),
.Y(n_2150)
);

OAI21x1_ASAP7_75t_L g2151 ( 
.A1(n_2062),
.A2(n_340),
.B(n_339),
.Y(n_2151)
);

INVx3_ASAP7_75t_L g2152 ( 
.A(n_2060),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2068),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2068),
.Y(n_2154)
);

OAI21x1_ASAP7_75t_L g2155 ( 
.A1(n_2062),
.A2(n_342),
.B(n_341),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_2045),
.B(n_36),
.Y(n_2156)
);

OAI21xp5_ASAP7_75t_L g2157 ( 
.A1(n_2059),
.A2(n_37),
.B(n_38),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2068),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2068),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2068),
.Y(n_2160)
);

OAI22xp5_ASAP7_75t_L g2161 ( 
.A1(n_2092),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2068),
.Y(n_2162)
);

AO21x2_ASAP7_75t_L g2163 ( 
.A1(n_2062),
.A2(n_39),
.B(n_40),
.Y(n_2163)
);

AO21x2_ASAP7_75t_L g2164 ( 
.A1(n_2062),
.A2(n_41),
.B(n_42),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2045),
.B(n_42),
.Y(n_2165)
);

CKINVDCx20_ASAP7_75t_R g2166 ( 
.A(n_2082),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2068),
.Y(n_2167)
);

BUFx2_ASAP7_75t_L g2168 ( 
.A(n_2045),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2068),
.Y(n_2169)
);

HB1xp67_ASAP7_75t_L g2170 ( 
.A(n_2094),
.Y(n_2170)
);

BUFx2_ASAP7_75t_L g2171 ( 
.A(n_2117),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2100),
.B(n_2168),
.Y(n_2172)
);

BUFx2_ASAP7_75t_L g2173 ( 
.A(n_2116),
.Y(n_2173)
);

BUFx2_ASAP7_75t_L g2174 ( 
.A(n_2136),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2147),
.Y(n_2175)
);

NOR2x1_ASAP7_75t_L g2176 ( 
.A(n_2118),
.B(n_43),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2148),
.Y(n_2177)
);

BUFx2_ASAP7_75t_L g2178 ( 
.A(n_2170),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_2097),
.Y(n_2179)
);

BUFx2_ASAP7_75t_L g2180 ( 
.A(n_2106),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2150),
.Y(n_2181)
);

INVx3_ASAP7_75t_L g2182 ( 
.A(n_2111),
.Y(n_2182)
);

CKINVDCx6p67_ASAP7_75t_R g2183 ( 
.A(n_2166),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2153),
.Y(n_2184)
);

NOR2xp33_ASAP7_75t_L g2185 ( 
.A(n_2125),
.B(n_43),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2154),
.Y(n_2186)
);

BUFx2_ASAP7_75t_L g2187 ( 
.A(n_2102),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_2096),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_2114),
.B(n_44),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_2119),
.B(n_44),
.Y(n_2190)
);

HB1xp67_ASAP7_75t_L g2191 ( 
.A(n_2101),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2158),
.Y(n_2192)
);

BUFx3_ASAP7_75t_L g2193 ( 
.A(n_2124),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_2169),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_2159),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2160),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_2112),
.B(n_45),
.Y(n_2197)
);

AO31x2_ASAP7_75t_L g2198 ( 
.A1(n_2140),
.A2(n_2123),
.A3(n_2141),
.B(n_2146),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_2162),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2167),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_2098),
.Y(n_2201)
);

INVx1_ASAP7_75t_SL g2202 ( 
.A(n_2110),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2133),
.Y(n_2203)
);

NOR2x1_ASAP7_75t_L g2204 ( 
.A(n_2127),
.B(n_45),
.Y(n_2204)
);

AOI22xp33_ASAP7_75t_L g2205 ( 
.A1(n_2145),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_2129),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2105),
.B(n_46),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2113),
.B(n_47),
.Y(n_2208)
);

OR2x2_ASAP7_75t_L g2209 ( 
.A(n_2126),
.B(n_2143),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_2099),
.B(n_48),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2138),
.Y(n_2211)
);

AND2x4_ASAP7_75t_L g2212 ( 
.A(n_2131),
.B(n_49),
.Y(n_2212)
);

HB1xp67_ASAP7_75t_L g2213 ( 
.A(n_2120),
.Y(n_2213)
);

INVxp67_ASAP7_75t_SL g2214 ( 
.A(n_2152),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2121),
.B(n_49),
.Y(n_2215)
);

OR2x2_ASAP7_75t_L g2216 ( 
.A(n_2135),
.B(n_50),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_2163),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_2164),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2109),
.Y(n_2219)
);

AND2x2_ASAP7_75t_L g2220 ( 
.A(n_2103),
.B(n_50),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_2156),
.B(n_51),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2165),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2132),
.B(n_52),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_2122),
.B(n_52),
.Y(n_2224)
);

HB1xp67_ASAP7_75t_L g2225 ( 
.A(n_2142),
.Y(n_2225)
);

OR2x2_ASAP7_75t_L g2226 ( 
.A(n_2144),
.B(n_53),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2145),
.B(n_53),
.Y(n_2227)
);

OR2x2_ASAP7_75t_L g2228 ( 
.A(n_2139),
.B(n_54),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_2130),
.B(n_55),
.Y(n_2229)
);

CKINVDCx5p33_ASAP7_75t_R g2230 ( 
.A(n_2134),
.Y(n_2230)
);

INVx1_ASAP7_75t_SL g2231 ( 
.A(n_2107),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_2108),
.B(n_56),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2151),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2157),
.B(n_56),
.Y(n_2234)
);

OR2x2_ASAP7_75t_L g2235 ( 
.A(n_2155),
.B(n_2128),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_2149),
.B(n_57),
.Y(n_2236)
);

INVx1_ASAP7_75t_SL g2237 ( 
.A(n_2137),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2115),
.Y(n_2238)
);

INVx3_ASAP7_75t_L g2239 ( 
.A(n_2137),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_2161),
.Y(n_2240)
);

AND2x2_ASAP7_75t_L g2241 ( 
.A(n_2095),
.B(n_57),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2104),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2147),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2147),
.Y(n_2244)
);

AO21x2_ASAP7_75t_L g2245 ( 
.A1(n_2123),
.A2(n_58),
.B(n_59),
.Y(n_2245)
);

AND2x2_ASAP7_75t_L g2246 ( 
.A(n_2100),
.B(n_59),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2147),
.Y(n_2247)
);

BUFx3_ASAP7_75t_L g2248 ( 
.A(n_2166),
.Y(n_2248)
);

INVx2_ASAP7_75t_SL g2249 ( 
.A(n_2100),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_2118),
.B(n_60),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2100),
.B(n_60),
.Y(n_2251)
);

AND2x2_ASAP7_75t_L g2252 ( 
.A(n_2100),
.B(n_61),
.Y(n_2252)
);

INVx3_ASAP7_75t_L g2253 ( 
.A(n_2111),
.Y(n_2253)
);

OR2x2_ASAP7_75t_L g2254 ( 
.A(n_2112),
.B(n_61),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2147),
.Y(n_2255)
);

INVx2_ASAP7_75t_L g2256 ( 
.A(n_2100),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_2100),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2147),
.Y(n_2258)
);

HB1xp67_ASAP7_75t_L g2259 ( 
.A(n_2170),
.Y(n_2259)
);

AOI22xp33_ASAP7_75t_L g2260 ( 
.A1(n_2146),
.A2(n_65),
.B1(n_62),
.B2(n_64),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2100),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_2100),
.B(n_64),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_2100),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_2100),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2147),
.Y(n_2265)
);

BUFx3_ASAP7_75t_L g2266 ( 
.A(n_2166),
.Y(n_2266)
);

OAI22xp33_ASAP7_75t_L g2267 ( 
.A1(n_2145),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_2100),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_2174),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_2172),
.B(n_66),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_2195),
.Y(n_2271)
);

AND2x4_ASAP7_75t_L g2272 ( 
.A(n_2249),
.B(n_2239),
.Y(n_2272)
);

INVx4_ASAP7_75t_R g2273 ( 
.A(n_2248),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_2173),
.B(n_68),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_2199),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2198),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2175),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_2198),
.Y(n_2278)
);

AOI22xp5_ASAP7_75t_L g2279 ( 
.A1(n_2234),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_2203),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2177),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2181),
.Y(n_2282)
);

HB1xp67_ASAP7_75t_L g2283 ( 
.A(n_2171),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2184),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2186),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2178),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_2256),
.B(n_69),
.Y(n_2287)
);

AND2x2_ASAP7_75t_L g2288 ( 
.A(n_2257),
.B(n_70),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_2261),
.B(n_71),
.Y(n_2289)
);

INVxp67_ASAP7_75t_L g2290 ( 
.A(n_2225),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_2192),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_2263),
.B(n_72),
.Y(n_2292)
);

OR2x2_ASAP7_75t_L g2293 ( 
.A(n_2259),
.B(n_72),
.Y(n_2293)
);

NOR4xp25_ASAP7_75t_SL g2294 ( 
.A(n_2171),
.B(n_2214),
.C(n_2233),
.D(n_2238),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_2264),
.B(n_73),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_2196),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2268),
.B(n_73),
.Y(n_2297)
);

BUFx12f_ASAP7_75t_L g2298 ( 
.A(n_2226),
.Y(n_2298)
);

OR2x2_ASAP7_75t_L g2299 ( 
.A(n_2209),
.B(n_74),
.Y(n_2299)
);

OR2x2_ASAP7_75t_L g2300 ( 
.A(n_2211),
.B(n_75),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2180),
.B(n_75),
.Y(n_2301)
);

AND2x4_ASAP7_75t_L g2302 ( 
.A(n_2182),
.B(n_2253),
.Y(n_2302)
);

AO31x2_ASAP7_75t_L g2303 ( 
.A1(n_2217),
.A2(n_78),
.A3(n_76),
.B(n_77),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_2200),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2243),
.Y(n_2305)
);

AND2x2_ASAP7_75t_L g2306 ( 
.A(n_2222),
.B(n_2187),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2213),
.B(n_77),
.Y(n_2307)
);

HB1xp67_ASAP7_75t_L g2308 ( 
.A(n_2191),
.Y(n_2308)
);

AND2x2_ASAP7_75t_L g2309 ( 
.A(n_2206),
.B(n_78),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_2201),
.B(n_79),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2244),
.Y(n_2311)
);

AND2x2_ASAP7_75t_L g2312 ( 
.A(n_2188),
.B(n_79),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2194),
.B(n_80),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_2247),
.Y(n_2314)
);

OR2x2_ASAP7_75t_L g2315 ( 
.A(n_2179),
.B(n_80),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_2255),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2258),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2265),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2254),
.Y(n_2319)
);

BUFx6f_ASAP7_75t_L g2320 ( 
.A(n_2212),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2218),
.Y(n_2321)
);

AND2x2_ASAP7_75t_L g2322 ( 
.A(n_2202),
.B(n_81),
.Y(n_2322)
);

AND2x2_ASAP7_75t_L g2323 ( 
.A(n_2189),
.B(n_2237),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_2216),
.Y(n_2324)
);

INVx3_ASAP7_75t_L g2325 ( 
.A(n_2193),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2197),
.Y(n_2326)
);

HB1xp67_ASAP7_75t_L g2327 ( 
.A(n_2176),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2219),
.B(n_81),
.Y(n_2328)
);

INVx2_ASAP7_75t_SL g2329 ( 
.A(n_2266),
.Y(n_2329)
);

AOI22xp33_ASAP7_75t_L g2330 ( 
.A1(n_2240),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_2330)
);

AO21x2_ASAP7_75t_L g2331 ( 
.A1(n_2250),
.A2(n_82),
.B(n_83),
.Y(n_2331)
);

AND2x2_ASAP7_75t_L g2332 ( 
.A(n_2231),
.B(n_84),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_2185),
.B(n_85),
.Y(n_2333)
);

INVx2_ASAP7_75t_SL g2334 ( 
.A(n_2183),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_2228),
.Y(n_2335)
);

AND2x2_ASAP7_75t_L g2336 ( 
.A(n_2246),
.B(n_2251),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2190),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2252),
.B(n_85),
.Y(n_2338)
);

INVx3_ASAP7_75t_L g2339 ( 
.A(n_2210),
.Y(n_2339)
);

INVxp67_ASAP7_75t_L g2340 ( 
.A(n_2204),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2245),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2262),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2208),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2235),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2227),
.Y(n_2345)
);

BUFx6f_ASAP7_75t_L g2346 ( 
.A(n_2220),
.Y(n_2346)
);

INVx3_ASAP7_75t_L g2347 ( 
.A(n_2215),
.Y(n_2347)
);

AND2x2_ASAP7_75t_L g2348 ( 
.A(n_2223),
.B(n_86),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_2221),
.B(n_86),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2232),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_2229),
.Y(n_2351)
);

INVx3_ASAP7_75t_L g2352 ( 
.A(n_2230),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2207),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2242),
.B(n_87),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2224),
.B(n_87),
.Y(n_2355)
);

AND2x2_ASAP7_75t_L g2356 ( 
.A(n_2241),
.B(n_88),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2267),
.B(n_88),
.Y(n_2357)
);

AOI22xp33_ASAP7_75t_L g2358 ( 
.A1(n_2236),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2205),
.Y(n_2359)
);

OR2x2_ASAP7_75t_SL g2360 ( 
.A(n_2260),
.B(n_89),
.Y(n_2360)
);

BUFx4f_ASAP7_75t_SL g2361 ( 
.A(n_2183),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_2174),
.Y(n_2362)
);

NOR2x1_ASAP7_75t_L g2363 ( 
.A(n_2171),
.B(n_90),
.Y(n_2363)
);

AND2x2_ASAP7_75t_L g2364 ( 
.A(n_2172),
.B(n_92),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2175),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_2174),
.Y(n_2366)
);

INVxp67_ASAP7_75t_SL g2367 ( 
.A(n_2225),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2172),
.B(n_92),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2259),
.B(n_94),
.Y(n_2369)
);

AND2x2_ASAP7_75t_L g2370 ( 
.A(n_2172),
.B(n_95),
.Y(n_2370)
);

AND2x2_ASAP7_75t_L g2371 ( 
.A(n_2172),
.B(n_95),
.Y(n_2371)
);

BUFx3_ASAP7_75t_L g2372 ( 
.A(n_2183),
.Y(n_2372)
);

INVxp67_ASAP7_75t_SL g2373 ( 
.A(n_2225),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_2174),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_2259),
.B(n_96),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_2172),
.B(n_96),
.Y(n_2376)
);

AND2x2_ASAP7_75t_L g2377 ( 
.A(n_2172),
.B(n_97),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2175),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2175),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2175),
.Y(n_2380)
);

AND2x2_ASAP7_75t_L g2381 ( 
.A(n_2172),
.B(n_97),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2175),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2259),
.B(n_98),
.Y(n_2383)
);

OR2x2_ASAP7_75t_L g2384 ( 
.A(n_2259),
.B(n_98),
.Y(n_2384)
);

NOR2x1_ASAP7_75t_L g2385 ( 
.A(n_2171),
.B(n_99),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2175),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2175),
.Y(n_2387)
);

BUFx6f_ASAP7_75t_L g2388 ( 
.A(n_2212),
.Y(n_2388)
);

OAI22xp5_ASAP7_75t_L g2389 ( 
.A1(n_2234),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2175),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2175),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2277),
.Y(n_2392)
);

HB1xp67_ASAP7_75t_L g2393 ( 
.A(n_2283),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2281),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2345),
.B(n_100),
.Y(n_2395)
);

INVx1_ASAP7_75t_SL g2396 ( 
.A(n_2361),
.Y(n_2396)
);

AND2x4_ASAP7_75t_L g2397 ( 
.A(n_2334),
.B(n_102),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2282),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2327),
.B(n_102),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_2276),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_L g2401 ( 
.A(n_2290),
.B(n_103),
.Y(n_2401)
);

AND2x2_ASAP7_75t_L g2402 ( 
.A(n_2351),
.B(n_104),
.Y(n_2402)
);

INVxp67_ASAP7_75t_SL g2403 ( 
.A(n_2340),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_2353),
.B(n_104),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_2278),
.Y(n_2405)
);

OR2x2_ASAP7_75t_L g2406 ( 
.A(n_2324),
.B(n_105),
.Y(n_2406)
);

INVxp67_ASAP7_75t_L g2407 ( 
.A(n_2363),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2284),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_2269),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2285),
.Y(n_2410)
);

INVx2_ASAP7_75t_SL g2411 ( 
.A(n_2273),
.Y(n_2411)
);

INVx3_ASAP7_75t_L g2412 ( 
.A(n_2302),
.Y(n_2412)
);

AND2x2_ASAP7_75t_L g2413 ( 
.A(n_2286),
.B(n_106),
.Y(n_2413)
);

AND2x2_ASAP7_75t_L g2414 ( 
.A(n_2350),
.B(n_106),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_2307),
.B(n_107),
.Y(n_2415)
);

HB1xp67_ASAP7_75t_L g2416 ( 
.A(n_2308),
.Y(n_2416)
);

AND2x2_ASAP7_75t_L g2417 ( 
.A(n_2335),
.B(n_108),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2343),
.B(n_108),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_2362),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2366),
.Y(n_2420)
);

AND2x2_ASAP7_75t_L g2421 ( 
.A(n_2374),
.B(n_109),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2272),
.B(n_109),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_2367),
.B(n_110),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_2271),
.Y(n_2424)
);

INVx1_ASAP7_75t_SL g2425 ( 
.A(n_2372),
.Y(n_2425)
);

INVxp67_ASAP7_75t_SL g2426 ( 
.A(n_2385),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2373),
.B(n_2341),
.Y(n_2427)
);

AND2x2_ASAP7_75t_L g2428 ( 
.A(n_2306),
.B(n_2323),
.Y(n_2428)
);

AND2x2_ASAP7_75t_L g2429 ( 
.A(n_2339),
.B(n_110),
.Y(n_2429)
);

INVxp67_ASAP7_75t_SL g2430 ( 
.A(n_2347),
.Y(n_2430)
);

INVx2_ASAP7_75t_SL g2431 ( 
.A(n_2320),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2305),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2319),
.B(n_111),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2317),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2318),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2312),
.B(n_111),
.Y(n_2436)
);

INVxp67_ASAP7_75t_SL g2437 ( 
.A(n_2346),
.Y(n_2437)
);

BUFx2_ASAP7_75t_L g2438 ( 
.A(n_2298),
.Y(n_2438)
);

INVx4_ASAP7_75t_L g2439 ( 
.A(n_2320),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_2275),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2365),
.Y(n_2441)
);

AND2x2_ASAP7_75t_L g2442 ( 
.A(n_2336),
.B(n_112),
.Y(n_2442)
);

HB1xp67_ASAP7_75t_L g2443 ( 
.A(n_2291),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2378),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2379),
.Y(n_2445)
);

INVx3_ASAP7_75t_L g2446 ( 
.A(n_2388),
.Y(n_2446)
);

INVx3_ASAP7_75t_L g2447 ( 
.A(n_2388),
.Y(n_2447)
);

NOR2xp67_ASAP7_75t_L g2448 ( 
.A(n_2321),
.B(n_112),
.Y(n_2448)
);

AND2x2_ASAP7_75t_L g2449 ( 
.A(n_2342),
.B(n_113),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_2280),
.Y(n_2450)
);

AND2x4_ASAP7_75t_L g2451 ( 
.A(n_2325),
.B(n_113),
.Y(n_2451)
);

INVx1_ASAP7_75t_SL g2452 ( 
.A(n_2274),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2380),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2337),
.B(n_114),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2313),
.B(n_114),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2309),
.B(n_115),
.Y(n_2456)
);

HB1xp67_ASAP7_75t_L g2457 ( 
.A(n_2296),
.Y(n_2457)
);

AND2x2_ASAP7_75t_L g2458 ( 
.A(n_2326),
.B(n_115),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2382),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2344),
.Y(n_2460)
);

INVxp67_ASAP7_75t_SL g2461 ( 
.A(n_2346),
.Y(n_2461)
);

HB1xp67_ASAP7_75t_L g2462 ( 
.A(n_2304),
.Y(n_2462)
);

INVxp67_ASAP7_75t_L g2463 ( 
.A(n_2331),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2311),
.Y(n_2464)
);

OR2x2_ASAP7_75t_L g2465 ( 
.A(n_2299),
.B(n_116),
.Y(n_2465)
);

AND2x4_ASAP7_75t_L g2466 ( 
.A(n_2329),
.B(n_2352),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_2310),
.B(n_116),
.Y(n_2467)
);

OR2x2_ASAP7_75t_L g2468 ( 
.A(n_2314),
.B(n_117),
.Y(n_2468)
);

AND2x4_ASAP7_75t_L g2469 ( 
.A(n_2301),
.B(n_117),
.Y(n_2469)
);

AND2x2_ASAP7_75t_L g2470 ( 
.A(n_2270),
.B(n_118),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2386),
.Y(n_2471)
);

INVxp67_ASAP7_75t_L g2472 ( 
.A(n_2315),
.Y(n_2472)
);

AND2x2_ASAP7_75t_L g2473 ( 
.A(n_2364),
.B(n_118),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2387),
.Y(n_2474)
);

NAND2xp33_ASAP7_75t_L g2475 ( 
.A(n_2357),
.B(n_119),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2316),
.Y(n_2476)
);

AND2x2_ASAP7_75t_L g2477 ( 
.A(n_2368),
.B(n_119),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_2390),
.Y(n_2478)
);

AND2x2_ASAP7_75t_L g2479 ( 
.A(n_2370),
.B(n_120),
.Y(n_2479)
);

AND2x2_ASAP7_75t_L g2480 ( 
.A(n_2371),
.B(n_121),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_2369),
.B(n_121),
.Y(n_2481)
);

HB1xp67_ASAP7_75t_L g2482 ( 
.A(n_2391),
.Y(n_2482)
);

AND2x2_ASAP7_75t_L g2483 ( 
.A(n_2376),
.B(n_122),
.Y(n_2483)
);

NOR2xp33_ASAP7_75t_L g2484 ( 
.A(n_2354),
.B(n_122),
.Y(n_2484)
);

AND2x2_ASAP7_75t_L g2485 ( 
.A(n_2377),
.B(n_123),
.Y(n_2485)
);

AND2x2_ASAP7_75t_L g2486 ( 
.A(n_2381),
.B(n_123),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2300),
.Y(n_2487)
);

NOR2xp33_ASAP7_75t_L g2488 ( 
.A(n_2333),
.B(n_124),
.Y(n_2488)
);

AND2x2_ASAP7_75t_L g2489 ( 
.A(n_2287),
.B(n_125),
.Y(n_2489)
);

O2A1O1Ixp33_ASAP7_75t_L g2490 ( 
.A1(n_2389),
.A2(n_129),
.B(n_130),
.C(n_128),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2303),
.Y(n_2491)
);

AND2x2_ASAP7_75t_L g2492 ( 
.A(n_2288),
.B(n_126),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2289),
.B(n_126),
.Y(n_2493)
);

AND2x4_ASAP7_75t_L g2494 ( 
.A(n_2292),
.B(n_128),
.Y(n_2494)
);

INVx1_ASAP7_75t_SL g2495 ( 
.A(n_2293),
.Y(n_2495)
);

OR2x2_ASAP7_75t_L g2496 ( 
.A(n_2384),
.B(n_129),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2303),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2295),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_2297),
.Y(n_2499)
);

AND2x2_ASAP7_75t_L g2500 ( 
.A(n_2328),
.B(n_130),
.Y(n_2500)
);

BUFx2_ASAP7_75t_L g2501 ( 
.A(n_2332),
.Y(n_2501)
);

OR2x2_ASAP7_75t_L g2502 ( 
.A(n_2375),
.B(n_131),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2322),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_2383),
.Y(n_2504)
);

AND2x4_ASAP7_75t_L g2505 ( 
.A(n_2359),
.B(n_131),
.Y(n_2505)
);

AND2x2_ASAP7_75t_L g2506 ( 
.A(n_2294),
.B(n_2349),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2338),
.Y(n_2507)
);

AND2x2_ASAP7_75t_L g2508 ( 
.A(n_2348),
.B(n_132),
.Y(n_2508)
);

OR2x2_ASAP7_75t_L g2509 ( 
.A(n_2355),
.B(n_133),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2356),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2360),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2279),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2358),
.Y(n_2513)
);

OR2x2_ASAP7_75t_L g2514 ( 
.A(n_2330),
.B(n_133),
.Y(n_2514)
);

AND2x4_ASAP7_75t_L g2515 ( 
.A(n_2334),
.B(n_134),
.Y(n_2515)
);

NOR2xp33_ASAP7_75t_L g2516 ( 
.A(n_2361),
.B(n_134),
.Y(n_2516)
);

AND2x2_ASAP7_75t_L g2517 ( 
.A(n_2351),
.B(n_135),
.Y(n_2517)
);

AND2x2_ASAP7_75t_L g2518 ( 
.A(n_2351),
.B(n_135),
.Y(n_2518)
);

OR2x2_ASAP7_75t_L g2519 ( 
.A(n_2324),
.B(n_136),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2345),
.B(n_136),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2276),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2277),
.Y(n_2522)
);

AND2x2_ASAP7_75t_L g2523 ( 
.A(n_2351),
.B(n_137),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2345),
.B(n_137),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2277),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2277),
.Y(n_2526)
);

AND2x2_ASAP7_75t_L g2527 ( 
.A(n_2351),
.B(n_138),
.Y(n_2527)
);

AND2x2_ASAP7_75t_L g2528 ( 
.A(n_2351),
.B(n_138),
.Y(n_2528)
);

BUFx2_ASAP7_75t_L g2529 ( 
.A(n_2340),
.Y(n_2529)
);

INVx2_ASAP7_75t_SL g2530 ( 
.A(n_2273),
.Y(n_2530)
);

AND2x2_ASAP7_75t_L g2531 ( 
.A(n_2351),
.B(n_139),
.Y(n_2531)
);

CKINVDCx11_ASAP7_75t_R g2532 ( 
.A(n_2298),
.Y(n_2532)
);

HB1xp67_ASAP7_75t_L g2533 ( 
.A(n_2283),
.Y(n_2533)
);

INVx2_ASAP7_75t_SL g2534 ( 
.A(n_2273),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2277),
.Y(n_2535)
);

INVx2_ASAP7_75t_L g2536 ( 
.A(n_2276),
.Y(n_2536)
);

HB1xp67_ASAP7_75t_L g2537 ( 
.A(n_2283),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2276),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2277),
.Y(n_2539)
);

INVx2_ASAP7_75t_L g2540 ( 
.A(n_2276),
.Y(n_2540)
);

BUFx3_ASAP7_75t_L g2541 ( 
.A(n_2372),
.Y(n_2541)
);

NOR2x1p5_ASAP7_75t_L g2542 ( 
.A(n_2372),
.B(n_139),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_2345),
.B(n_140),
.Y(n_2543)
);

HB1xp67_ASAP7_75t_L g2544 ( 
.A(n_2283),
.Y(n_2544)
);

AND2x2_ASAP7_75t_L g2545 ( 
.A(n_2351),
.B(n_140),
.Y(n_2545)
);

AND2x4_ASAP7_75t_SL g2546 ( 
.A(n_2325),
.B(n_141),
.Y(n_2546)
);

OR2x2_ASAP7_75t_L g2547 ( 
.A(n_2324),
.B(n_141),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2276),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2345),
.B(n_142),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2277),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2345),
.B(n_142),
.Y(n_2551)
);

INVx4_ASAP7_75t_L g2552 ( 
.A(n_2361),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2276),
.Y(n_2553)
);

INVx2_ASAP7_75t_SL g2554 ( 
.A(n_2273),
.Y(n_2554)
);

OR2x2_ASAP7_75t_L g2555 ( 
.A(n_2324),
.B(n_143),
.Y(n_2555)
);

INVx3_ASAP7_75t_L g2556 ( 
.A(n_2302),
.Y(n_2556)
);

AND2x2_ASAP7_75t_L g2557 ( 
.A(n_2351),
.B(n_143),
.Y(n_2557)
);

INVx2_ASAP7_75t_SL g2558 ( 
.A(n_2273),
.Y(n_2558)
);

BUFx6f_ASAP7_75t_L g2559 ( 
.A(n_2372),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2277),
.Y(n_2560)
);

INVx3_ASAP7_75t_L g2561 ( 
.A(n_2302),
.Y(n_2561)
);

OR2x2_ASAP7_75t_L g2562 ( 
.A(n_2324),
.B(n_144),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2482),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2392),
.Y(n_2564)
);

HB1xp67_ASAP7_75t_L g2565 ( 
.A(n_2529),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2394),
.Y(n_2566)
);

NOR3xp33_ASAP7_75t_L g2567 ( 
.A(n_2475),
.B(n_146),
.C(n_147),
.Y(n_2567)
);

AOI21xp5_ASAP7_75t_L g2568 ( 
.A1(n_2426),
.A2(n_146),
.B(n_148),
.Y(n_2568)
);

INVx3_ASAP7_75t_L g2569 ( 
.A(n_2552),
.Y(n_2569)
);

OAI31xp33_ASAP7_75t_L g2570 ( 
.A1(n_2506),
.A2(n_2407),
.A3(n_2463),
.B(n_2511),
.Y(n_2570)
);

INVx3_ASAP7_75t_L g2571 ( 
.A(n_2559),
.Y(n_2571)
);

INVxp67_ASAP7_75t_SL g2572 ( 
.A(n_2448),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_L g2573 ( 
.A(n_2403),
.B(n_149),
.Y(n_2573)
);

INVxp67_ASAP7_75t_SL g2574 ( 
.A(n_2393),
.Y(n_2574)
);

NAND3xp33_ASAP7_75t_L g2575 ( 
.A(n_2490),
.B(n_149),
.C(n_150),
.Y(n_2575)
);

AND2x4_ASAP7_75t_L g2576 ( 
.A(n_2411),
.B(n_150),
.Y(n_2576)
);

AOI22xp33_ASAP7_75t_L g2577 ( 
.A1(n_2512),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_2577)
);

OR2x6_ASAP7_75t_L g2578 ( 
.A(n_2530),
.B(n_151),
.Y(n_2578)
);

INVx1_ASAP7_75t_SL g2579 ( 
.A(n_2532),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2398),
.Y(n_2580)
);

INVxp67_ASAP7_75t_SL g2581 ( 
.A(n_2533),
.Y(n_2581)
);

AO21x2_ASAP7_75t_L g2582 ( 
.A1(n_2423),
.A2(n_153),
.B(n_154),
.Y(n_2582)
);

INVx5_ASAP7_75t_L g2583 ( 
.A(n_2559),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2408),
.Y(n_2584)
);

HB1xp67_ASAP7_75t_L g2585 ( 
.A(n_2537),
.Y(n_2585)
);

AOI22xp5_ASAP7_75t_L g2586 ( 
.A1(n_2430),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_2586)
);

AND2x2_ASAP7_75t_L g2587 ( 
.A(n_2428),
.B(n_157),
.Y(n_2587)
);

HB1xp67_ASAP7_75t_L g2588 ( 
.A(n_2544),
.Y(n_2588)
);

INVx2_ASAP7_75t_L g2589 ( 
.A(n_2438),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2410),
.Y(n_2590)
);

AO21x2_ASAP7_75t_L g2591 ( 
.A1(n_2399),
.A2(n_157),
.B(n_158),
.Y(n_2591)
);

NOR2xp67_ASAP7_75t_L g2592 ( 
.A(n_2534),
.B(n_158),
.Y(n_2592)
);

AOI222xp33_ASAP7_75t_L g2593 ( 
.A1(n_2513),
.A2(n_161),
.B1(n_163),
.B2(n_159),
.C1(n_160),
.C2(n_162),
.Y(n_2593)
);

INVx2_ASAP7_75t_L g2594 ( 
.A(n_2439),
.Y(n_2594)
);

AND2x2_ASAP7_75t_L g2595 ( 
.A(n_2412),
.B(n_159),
.Y(n_2595)
);

INVx2_ASAP7_75t_L g2596 ( 
.A(n_2446),
.Y(n_2596)
);

INVx2_ASAP7_75t_L g2597 ( 
.A(n_2447),
.Y(n_2597)
);

OR2x2_ASAP7_75t_L g2598 ( 
.A(n_2409),
.B(n_2419),
.Y(n_2598)
);

BUFx2_ASAP7_75t_L g2599 ( 
.A(n_2554),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2432),
.Y(n_2600)
);

OAI33xp33_ASAP7_75t_L g2601 ( 
.A1(n_2491),
.A2(n_162),
.A3(n_165),
.B1(n_160),
.B2(n_161),
.B3(n_164),
.Y(n_2601)
);

HB1xp67_ASAP7_75t_L g2602 ( 
.A(n_2416),
.Y(n_2602)
);

INVxp67_ASAP7_75t_SL g2603 ( 
.A(n_2558),
.Y(n_2603)
);

INVx3_ASAP7_75t_L g2604 ( 
.A(n_2541),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2434),
.Y(n_2605)
);

INVx2_ASAP7_75t_SL g2606 ( 
.A(n_2466),
.Y(n_2606)
);

OAI221xp5_ASAP7_75t_L g2607 ( 
.A1(n_2437),
.A2(n_168),
.B1(n_165),
.B2(n_166),
.C(n_169),
.Y(n_2607)
);

INVx2_ASAP7_75t_SL g2608 ( 
.A(n_2396),
.Y(n_2608)
);

AOI22xp33_ASAP7_75t_L g2609 ( 
.A1(n_2507),
.A2(n_170),
.B1(n_166),
.B2(n_169),
.Y(n_2609)
);

AOI22xp5_ASAP7_75t_L g2610 ( 
.A1(n_2461),
.A2(n_173),
.B1(n_171),
.B2(n_172),
.Y(n_2610)
);

AND2x2_ASAP7_75t_L g2611 ( 
.A(n_2556),
.B(n_171),
.Y(n_2611)
);

INVx2_ASAP7_75t_L g2612 ( 
.A(n_2431),
.Y(n_2612)
);

HB1xp67_ASAP7_75t_L g2613 ( 
.A(n_2501),
.Y(n_2613)
);

OAI222xp33_ASAP7_75t_L g2614 ( 
.A1(n_2452),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.C1(n_174),
.C2(n_176),
.Y(n_2614)
);

INVx4_ASAP7_75t_L g2615 ( 
.A(n_2451),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_2561),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2435),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2400),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2441),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2444),
.Y(n_2620)
);

AND2x4_ASAP7_75t_L g2621 ( 
.A(n_2425),
.B(n_173),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2405),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_2487),
.B(n_174),
.Y(n_2623)
);

OAI211xp5_ASAP7_75t_L g2624 ( 
.A1(n_2427),
.A2(n_179),
.B(n_175),
.C(n_176),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2521),
.Y(n_2625)
);

AOI222xp33_ASAP7_75t_L g2626 ( 
.A1(n_2488),
.A2(n_2484),
.B1(n_2472),
.B2(n_2415),
.C1(n_2481),
.C2(n_2495),
.Y(n_2626)
);

AOI22xp33_ASAP7_75t_L g2627 ( 
.A1(n_2504),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_2627)
);

INVxp67_ASAP7_75t_SL g2628 ( 
.A(n_2542),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2536),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2445),
.Y(n_2630)
);

BUFx3_ASAP7_75t_L g2631 ( 
.A(n_2546),
.Y(n_2631)
);

INVx2_ASAP7_75t_L g2632 ( 
.A(n_2538),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2453),
.Y(n_2633)
);

INVx2_ASAP7_75t_L g2634 ( 
.A(n_2540),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2459),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2471),
.Y(n_2636)
);

AO21x2_ASAP7_75t_L g2637 ( 
.A1(n_2401),
.A2(n_180),
.B(n_182),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2474),
.Y(n_2638)
);

AND2x2_ASAP7_75t_L g2639 ( 
.A(n_2420),
.B(n_182),
.Y(n_2639)
);

AND2x2_ASAP7_75t_L g2640 ( 
.A(n_2503),
.B(n_183),
.Y(n_2640)
);

AND2x2_ASAP7_75t_L g2641 ( 
.A(n_2510),
.B(n_183),
.Y(n_2641)
);

OR2x2_ASAP7_75t_L g2642 ( 
.A(n_2424),
.B(n_184),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2522),
.Y(n_2643)
);

AND2x2_ASAP7_75t_L g2644 ( 
.A(n_2498),
.B(n_184),
.Y(n_2644)
);

INVxp67_ASAP7_75t_SL g2645 ( 
.A(n_2443),
.Y(n_2645)
);

INVx1_ASAP7_75t_SL g2646 ( 
.A(n_2397),
.Y(n_2646)
);

AOI21x1_ASAP7_75t_L g2647 ( 
.A1(n_2395),
.A2(n_2524),
.B(n_2520),
.Y(n_2647)
);

BUFx2_ASAP7_75t_L g2648 ( 
.A(n_2515),
.Y(n_2648)
);

OAI21x1_ASAP7_75t_SL g2649 ( 
.A1(n_2433),
.A2(n_185),
.B(n_186),
.Y(n_2649)
);

AND2x4_ASAP7_75t_L g2650 ( 
.A(n_2499),
.B(n_187),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2525),
.Y(n_2651)
);

BUFx3_ASAP7_75t_L g2652 ( 
.A(n_2494),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2526),
.Y(n_2653)
);

HB1xp67_ASAP7_75t_L g2654 ( 
.A(n_2457),
.Y(n_2654)
);

INVx2_ASAP7_75t_L g2655 ( 
.A(n_2548),
.Y(n_2655)
);

OR2x2_ASAP7_75t_L g2656 ( 
.A(n_2440),
.B(n_187),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_L g2657 ( 
.A(n_2414),
.B(n_188),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2535),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2539),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2553),
.Y(n_2660)
);

INVx3_ASAP7_75t_L g2661 ( 
.A(n_2505),
.Y(n_2661)
);

BUFx2_ASAP7_75t_L g2662 ( 
.A(n_2462),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2550),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2560),
.Y(n_2664)
);

AOI221xp5_ASAP7_75t_SL g2665 ( 
.A1(n_2497),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.C(n_191),
.Y(n_2665)
);

INVx2_ASAP7_75t_SL g2666 ( 
.A(n_2422),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2478),
.Y(n_2667)
);

INVxp67_ASAP7_75t_SL g2668 ( 
.A(n_2468),
.Y(n_2668)
);

INVx2_ASAP7_75t_SL g2669 ( 
.A(n_2429),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2449),
.B(n_189),
.Y(n_2670)
);

NAND4xp25_ASAP7_75t_L g2671 ( 
.A(n_2516),
.B(n_193),
.C(n_194),
.D(n_192),
.Y(n_2671)
);

AND2x2_ASAP7_75t_L g2672 ( 
.A(n_2460),
.B(n_191),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_2454),
.B(n_192),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2450),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2464),
.Y(n_2675)
);

AO21x2_ASAP7_75t_L g2676 ( 
.A1(n_2418),
.A2(n_193),
.B(n_196),
.Y(n_2676)
);

AOI31xp33_ASAP7_75t_L g2677 ( 
.A1(n_2514),
.A2(n_198),
.A3(n_196),
.B(n_197),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2476),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2406),
.Y(n_2679)
);

AND2x2_ASAP7_75t_L g2680 ( 
.A(n_2458),
.B(n_197),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_L g2681 ( 
.A(n_2404),
.B(n_199),
.Y(n_2681)
);

AND4x1_ASAP7_75t_L g2682 ( 
.A(n_2442),
.B(n_2500),
.C(n_2517),
.D(n_2402),
.Y(n_2682)
);

INVx1_ASAP7_75t_SL g2683 ( 
.A(n_2465),
.Y(n_2683)
);

INVx2_ASAP7_75t_L g2684 ( 
.A(n_2519),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2547),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2613),
.Y(n_2686)
);

OR2x2_ASAP7_75t_L g2687 ( 
.A(n_2683),
.B(n_2555),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2602),
.Y(n_2688)
);

NOR2xp33_ASAP7_75t_L g2689 ( 
.A(n_2579),
.B(n_2543),
.Y(n_2689)
);

BUFx3_ASAP7_75t_L g2690 ( 
.A(n_2583),
.Y(n_2690)
);

AND2x2_ASAP7_75t_L g2691 ( 
.A(n_2599),
.B(n_2413),
.Y(n_2691)
);

OR2x2_ASAP7_75t_L g2692 ( 
.A(n_2565),
.B(n_2684),
.Y(n_2692)
);

AND2x2_ASAP7_75t_L g2693 ( 
.A(n_2603),
.B(n_2421),
.Y(n_2693)
);

INVx2_ASAP7_75t_L g2694 ( 
.A(n_2583),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2585),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2588),
.Y(n_2696)
);

AND2x2_ASAP7_75t_L g2697 ( 
.A(n_2589),
.B(n_2417),
.Y(n_2697)
);

AND2x2_ASAP7_75t_L g2698 ( 
.A(n_2604),
.B(n_2531),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2654),
.Y(n_2699)
);

AND2x2_ASAP7_75t_L g2700 ( 
.A(n_2594),
.B(n_2545),
.Y(n_2700)
);

AND2x2_ASAP7_75t_L g2701 ( 
.A(n_2606),
.B(n_2608),
.Y(n_2701)
);

INVx3_ASAP7_75t_L g2702 ( 
.A(n_2615),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2662),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2572),
.B(n_2549),
.Y(n_2704)
);

NAND2x1p5_ASAP7_75t_L g2705 ( 
.A(n_2571),
.B(n_2562),
.Y(n_2705)
);

OR2x2_ASAP7_75t_L g2706 ( 
.A(n_2668),
.B(n_2551),
.Y(n_2706)
);

INVx3_ASAP7_75t_L g2707 ( 
.A(n_2569),
.Y(n_2707)
);

INVx1_ASAP7_75t_SL g2708 ( 
.A(n_2648),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2628),
.B(n_2518),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2645),
.Y(n_2710)
);

AND2x2_ASAP7_75t_L g2711 ( 
.A(n_2661),
.B(n_2523),
.Y(n_2711)
);

AND2x2_ASAP7_75t_L g2712 ( 
.A(n_2612),
.B(n_2527),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2574),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2669),
.B(n_2626),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2581),
.B(n_2528),
.Y(n_2715)
);

NOR2x1_ASAP7_75t_L g2716 ( 
.A(n_2592),
.B(n_2496),
.Y(n_2716)
);

AND2x2_ASAP7_75t_L g2717 ( 
.A(n_2596),
.B(n_2557),
.Y(n_2717)
);

AND2x4_ASAP7_75t_L g2718 ( 
.A(n_2652),
.B(n_2469),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2591),
.B(n_2489),
.Y(n_2719)
);

AND2x2_ASAP7_75t_L g2720 ( 
.A(n_2597),
.B(n_2492),
.Y(n_2720)
);

AND2x2_ASAP7_75t_L g2721 ( 
.A(n_2616),
.B(n_2493),
.Y(n_2721)
);

AND2x2_ASAP7_75t_L g2722 ( 
.A(n_2666),
.B(n_2508),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2564),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2566),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2580),
.Y(n_2725)
);

INVxp67_ASAP7_75t_L g2726 ( 
.A(n_2578),
.Y(n_2726)
);

NOR2xp33_ASAP7_75t_L g2727 ( 
.A(n_2682),
.B(n_2502),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2679),
.B(n_2470),
.Y(n_2728)
);

OR2x2_ASAP7_75t_L g2729 ( 
.A(n_2685),
.B(n_2509),
.Y(n_2729)
);

HB1xp67_ASAP7_75t_L g2730 ( 
.A(n_2563),
.Y(n_2730)
);

OR2x6_ASAP7_75t_L g2731 ( 
.A(n_2578),
.B(n_2473),
.Y(n_2731)
);

AND2x2_ASAP7_75t_L g2732 ( 
.A(n_2646),
.B(n_2477),
.Y(n_2732)
);

AND2x2_ASAP7_75t_L g2733 ( 
.A(n_2631),
.B(n_2479),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2582),
.B(n_2637),
.Y(n_2734)
);

HB1xp67_ASAP7_75t_L g2735 ( 
.A(n_2598),
.Y(n_2735)
);

AND2x2_ASAP7_75t_L g2736 ( 
.A(n_2587),
.B(n_2480),
.Y(n_2736)
);

NOR2x1p5_ASAP7_75t_L g2737 ( 
.A(n_2671),
.B(n_2467),
.Y(n_2737)
);

INVx2_ASAP7_75t_L g2738 ( 
.A(n_2642),
.Y(n_2738)
);

AND2x2_ASAP7_75t_L g2739 ( 
.A(n_2641),
.B(n_2483),
.Y(n_2739)
);

AND2x2_ASAP7_75t_L g2740 ( 
.A(n_2595),
.B(n_2485),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2584),
.Y(n_2741)
);

AND2x2_ASAP7_75t_L g2742 ( 
.A(n_2611),
.B(n_2486),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2676),
.B(n_2436),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2570),
.B(n_2455),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2590),
.Y(n_2745)
);

AND2x2_ASAP7_75t_L g2746 ( 
.A(n_2690),
.B(n_2647),
.Y(n_2746)
);

INVx1_ASAP7_75t_SL g2747 ( 
.A(n_2716),
.Y(n_2747)
);

NOR2xp33_ASAP7_75t_L g2748 ( 
.A(n_2707),
.B(n_2573),
.Y(n_2748)
);

AOI22xp5_ASAP7_75t_L g2749 ( 
.A1(n_2727),
.A2(n_2567),
.B1(n_2665),
.B2(n_2575),
.Y(n_2749)
);

OR2x2_ASAP7_75t_L g2750 ( 
.A(n_2708),
.B(n_2678),
.Y(n_2750)
);

INVx2_ASAP7_75t_L g2751 ( 
.A(n_2694),
.Y(n_2751)
);

INVx2_ASAP7_75t_L g2752 ( 
.A(n_2702),
.Y(n_2752)
);

AND2x2_ASAP7_75t_L g2753 ( 
.A(n_2701),
.B(n_2576),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2735),
.Y(n_2754)
);

AND2x2_ASAP7_75t_L g2755 ( 
.A(n_2691),
.B(n_2726),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2730),
.Y(n_2756)
);

AND2x2_ASAP7_75t_L g2757 ( 
.A(n_2693),
.B(n_2674),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2732),
.B(n_2568),
.Y(n_2758)
);

AND2x2_ASAP7_75t_L g2759 ( 
.A(n_2733),
.B(n_2675),
.Y(n_2759)
);

NOR2xp33_ASAP7_75t_SL g2760 ( 
.A(n_2718),
.B(n_2614),
.Y(n_2760)
);

AND2x2_ASAP7_75t_L g2761 ( 
.A(n_2698),
.B(n_2621),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2739),
.B(n_2677),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2713),
.Y(n_2763)
);

INVxp67_ASAP7_75t_L g2764 ( 
.A(n_2731),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2710),
.Y(n_2765)
);

OR2x2_ASAP7_75t_L g2766 ( 
.A(n_2692),
.B(n_2667),
.Y(n_2766)
);

OR2x2_ASAP7_75t_L g2767 ( 
.A(n_2715),
.B(n_2623),
.Y(n_2767)
);

AOI22x1_ASAP7_75t_SL g2768 ( 
.A1(n_2703),
.A2(n_2593),
.B1(n_2605),
.B2(n_2600),
.Y(n_2768)
);

OR2x2_ASAP7_75t_L g2769 ( 
.A(n_2686),
.B(n_2656),
.Y(n_2769)
);

INVx2_ASAP7_75t_L g2770 ( 
.A(n_2731),
.Y(n_2770)
);

AND2x2_ASAP7_75t_SL g2771 ( 
.A(n_2734),
.B(n_2577),
.Y(n_2771)
);

AND2x2_ASAP7_75t_L g2772 ( 
.A(n_2711),
.B(n_2680),
.Y(n_2772)
);

HB1xp67_ASAP7_75t_L g2773 ( 
.A(n_2705),
.Y(n_2773)
);

AND2x2_ASAP7_75t_L g2774 ( 
.A(n_2720),
.B(n_2644),
.Y(n_2774)
);

INVx1_ASAP7_75t_SL g2775 ( 
.A(n_2687),
.Y(n_2775)
);

BUFx6f_ASAP7_75t_L g2776 ( 
.A(n_2699),
.Y(n_2776)
);

INVx2_ASAP7_75t_SL g2777 ( 
.A(n_2722),
.Y(n_2777)
);

AND2x2_ASAP7_75t_L g2778 ( 
.A(n_2753),
.B(n_2721),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2755),
.Y(n_2779)
);

OAI32xp33_ASAP7_75t_L g2780 ( 
.A1(n_2747),
.A2(n_2744),
.A3(n_2714),
.B1(n_2719),
.B2(n_2743),
.Y(n_2780)
);

AND2x2_ASAP7_75t_L g2781 ( 
.A(n_2761),
.B(n_2697),
.Y(n_2781)
);

NOR2xp33_ASAP7_75t_L g2782 ( 
.A(n_2764),
.B(n_2709),
.Y(n_2782)
);

AOI21xp33_ASAP7_75t_L g2783 ( 
.A1(n_2771),
.A2(n_2695),
.B(n_2688),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_L g2784 ( 
.A(n_2760),
.B(n_2712),
.Y(n_2784)
);

INVx2_ASAP7_75t_L g2785 ( 
.A(n_2770),
.Y(n_2785)
);

INVx2_ASAP7_75t_L g2786 ( 
.A(n_2751),
.Y(n_2786)
);

AND2x2_ASAP7_75t_L g2787 ( 
.A(n_2772),
.B(n_2700),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2754),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2752),
.Y(n_2789)
);

AND2x2_ASAP7_75t_L g2790 ( 
.A(n_2773),
.B(n_2774),
.Y(n_2790)
);

NAND2xp33_ASAP7_75t_R g2791 ( 
.A(n_2768),
.B(n_2689),
.Y(n_2791)
);

BUFx2_ASAP7_75t_L g2792 ( 
.A(n_2746),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2777),
.B(n_2775),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2756),
.Y(n_2794)
);

AO21x1_ASAP7_75t_L g2795 ( 
.A1(n_2749),
.A2(n_2704),
.B(n_2696),
.Y(n_2795)
);

INVx2_ASAP7_75t_L g2796 ( 
.A(n_2776),
.Y(n_2796)
);

INVx1_ASAP7_75t_SL g2797 ( 
.A(n_2750),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2779),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2793),
.Y(n_2799)
);

OR2x2_ASAP7_75t_L g2800 ( 
.A(n_2797),
.B(n_2762),
.Y(n_2800)
);

AND2x2_ASAP7_75t_L g2801 ( 
.A(n_2790),
.B(n_2759),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2785),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2792),
.B(n_2776),
.Y(n_2803)
);

OR2x2_ASAP7_75t_L g2804 ( 
.A(n_2784),
.B(n_2769),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2788),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2786),
.Y(n_2806)
);

OR2x2_ASAP7_75t_L g2807 ( 
.A(n_2789),
.B(n_2766),
.Y(n_2807)
);

AOI222xp33_ASAP7_75t_L g2808 ( 
.A1(n_2799),
.A2(n_2780),
.B1(n_2782),
.B2(n_2763),
.C1(n_2765),
.C2(n_2794),
.Y(n_2808)
);

OAI21xp33_ASAP7_75t_L g2809 ( 
.A1(n_2801),
.A2(n_2783),
.B(n_2787),
.Y(n_2809)
);

NOR2xp33_ASAP7_75t_L g2810 ( 
.A(n_2803),
.B(n_2778),
.Y(n_2810)
);

AND2x2_ASAP7_75t_L g2811 ( 
.A(n_2802),
.B(n_2781),
.Y(n_2811)
);

AOI21xp33_ASAP7_75t_L g2812 ( 
.A1(n_2800),
.A2(n_2791),
.B(n_2795),
.Y(n_2812)
);

OAI22xp5_ASAP7_75t_L g2813 ( 
.A1(n_2804),
.A2(n_2758),
.B1(n_2796),
.B2(n_2748),
.Y(n_2813)
);

AOI22xp5_ASAP7_75t_L g2814 ( 
.A1(n_2798),
.A2(n_2757),
.B1(n_2738),
.B2(n_2601),
.Y(n_2814)
);

OAI221xp5_ASAP7_75t_L g2815 ( 
.A1(n_2807),
.A2(n_2767),
.B1(n_2586),
.B2(n_2610),
.C(n_2706),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_L g2816 ( 
.A(n_2806),
.B(n_2717),
.Y(n_2816)
);

HB1xp67_ASAP7_75t_L g2817 ( 
.A(n_2811),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2816),
.Y(n_2818)
);

AND2x2_ASAP7_75t_L g2819 ( 
.A(n_2810),
.B(n_2736),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_2809),
.B(n_2740),
.Y(n_2820)
);

NOR2xp33_ASAP7_75t_L g2821 ( 
.A(n_2812),
.B(n_2728),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2808),
.B(n_2742),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2813),
.Y(n_2823)
);

O2A1O1Ixp5_ASAP7_75t_L g2824 ( 
.A1(n_2814),
.A2(n_2805),
.B(n_2624),
.C(n_2724),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_2815),
.B(n_2729),
.Y(n_2825)
);

NOR2xp33_ASAP7_75t_L g2826 ( 
.A(n_2812),
.B(n_2723),
.Y(n_2826)
);

CKINVDCx20_ASAP7_75t_R g2827 ( 
.A(n_2810),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_2809),
.B(n_2737),
.Y(n_2828)
);

INVx2_ASAP7_75t_L g2829 ( 
.A(n_2811),
.Y(n_2829)
);

INVxp67_ASAP7_75t_L g2830 ( 
.A(n_2810),
.Y(n_2830)
);

INVx1_ASAP7_75t_SL g2831 ( 
.A(n_2811),
.Y(n_2831)
);

OAI21xp33_ASAP7_75t_L g2832 ( 
.A1(n_2809),
.A2(n_2741),
.B(n_2725),
.Y(n_2832)
);

AND2x2_ASAP7_75t_L g2833 ( 
.A(n_2811),
.B(n_2745),
.Y(n_2833)
);

AND2x2_ASAP7_75t_L g2834 ( 
.A(n_2811),
.B(n_2640),
.Y(n_2834)
);

NOR2xp33_ASAP7_75t_L g2835 ( 
.A(n_2827),
.B(n_2681),
.Y(n_2835)
);

HB1xp67_ASAP7_75t_L g2836 ( 
.A(n_2817),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_SL g2837 ( 
.A(n_2831),
.B(n_2819),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2834),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2829),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_L g2840 ( 
.A(n_2833),
.B(n_2822),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_2830),
.B(n_2617),
.Y(n_2841)
);

NAND3xp33_ASAP7_75t_L g2842 ( 
.A(n_2824),
.B(n_2607),
.C(n_2609),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2820),
.Y(n_2843)
);

INVx3_ASAP7_75t_SL g2844 ( 
.A(n_2823),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_2821),
.B(n_2619),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2828),
.Y(n_2846)
);

INVxp67_ASAP7_75t_SL g2847 ( 
.A(n_2825),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2832),
.Y(n_2848)
);

NAND2x1p5_ASAP7_75t_L g2849 ( 
.A(n_2818),
.B(n_2639),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2826),
.Y(n_2850)
);

OR2x2_ASAP7_75t_L g2851 ( 
.A(n_2831),
.B(n_2620),
.Y(n_2851)
);

O2A1O1Ixp5_ASAP7_75t_L g2852 ( 
.A1(n_2824),
.A2(n_2618),
.B(n_2625),
.C(n_2622),
.Y(n_2852)
);

AND2x2_ASAP7_75t_L g2853 ( 
.A(n_2819),
.B(n_2630),
.Y(n_2853)
);

AOI221xp5_ASAP7_75t_L g2854 ( 
.A1(n_2824),
.A2(n_2649),
.B1(n_2627),
.B2(n_2670),
.C(n_2657),
.Y(n_2854)
);

INVx2_ASAP7_75t_L g2855 ( 
.A(n_2849),
.Y(n_2855)
);

AND2x2_ASAP7_75t_L g2856 ( 
.A(n_2838),
.B(n_2643),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2836),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_L g2858 ( 
.A(n_2835),
.B(n_2651),
.Y(n_2858)
);

AOI211xp5_ASAP7_75t_L g2859 ( 
.A1(n_2837),
.A2(n_2673),
.B(n_2672),
.C(n_2456),
.Y(n_2859)
);

NAND4xp25_ASAP7_75t_L g2860 ( 
.A(n_2840),
.B(n_2650),
.C(n_2653),
.D(n_2633),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_L g2861 ( 
.A(n_2854),
.B(n_2659),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_L g2862 ( 
.A(n_2844),
.B(n_2663),
.Y(n_2862)
);

AND2x2_ASAP7_75t_L g2863 ( 
.A(n_2853),
.B(n_2839),
.Y(n_2863)
);

OR2x2_ASAP7_75t_L g2864 ( 
.A(n_2842),
.B(n_2635),
.Y(n_2864)
);

AOI211x1_ASAP7_75t_L g2865 ( 
.A1(n_2848),
.A2(n_2638),
.B(n_2658),
.C(n_2636),
.Y(n_2865)
);

NOR3xp33_ASAP7_75t_SL g2866 ( 
.A(n_2847),
.B(n_2664),
.C(n_199),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_L g2867 ( 
.A(n_2843),
.B(n_2632),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2850),
.B(n_2634),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_SL g2869 ( 
.A(n_2852),
.B(n_2629),
.Y(n_2869)
);

NOR3xp33_ASAP7_75t_L g2870 ( 
.A(n_2846),
.B(n_2655),
.C(n_2660),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2851),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2845),
.Y(n_2872)
);

NOR2xp33_ASAP7_75t_L g2873 ( 
.A(n_2841),
.B(n_200),
.Y(n_2873)
);

OR2x2_ASAP7_75t_L g2874 ( 
.A(n_2836),
.B(n_201),
.Y(n_2874)
);

AOI22xp5_ASAP7_75t_L g2875 ( 
.A1(n_2842),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.Y(n_2875)
);

NAND3xp33_ASAP7_75t_L g2876 ( 
.A(n_2866),
.B(n_202),
.C(n_203),
.Y(n_2876)
);

NOR2xp33_ASAP7_75t_L g2877 ( 
.A(n_2857),
.B(n_204),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_SL g2878 ( 
.A(n_2855),
.B(n_204),
.Y(n_2878)
);

NAND3xp33_ASAP7_75t_L g2879 ( 
.A(n_2875),
.B(n_2874),
.C(n_2873),
.Y(n_2879)
);

NOR4xp75_ASAP7_75t_L g2880 ( 
.A(n_2862),
.B(n_208),
.C(n_206),
.D(n_207),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_SL g2881 ( 
.A(n_2859),
.B(n_207),
.Y(n_2881)
);

NAND4xp25_ASAP7_75t_L g2882 ( 
.A(n_2870),
.B(n_2864),
.C(n_2861),
.D(n_2865),
.Y(n_2882)
);

NOR4xp25_ASAP7_75t_L g2883 ( 
.A(n_2871),
.B(n_210),
.C(n_208),
.D(n_209),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2863),
.Y(n_2884)
);

NAND4xp25_ASAP7_75t_SL g2885 ( 
.A(n_2867),
.B(n_212),
.C(n_209),
.D(n_211),
.Y(n_2885)
);

NOR3xp33_ASAP7_75t_L g2886 ( 
.A(n_2872),
.B(n_213),
.C(n_212),
.Y(n_2886)
);

NOR3xp33_ASAP7_75t_L g2887 ( 
.A(n_2868),
.B(n_2858),
.C(n_2869),
.Y(n_2887)
);

OAI211xp5_ASAP7_75t_SL g2888 ( 
.A1(n_2856),
.A2(n_214),
.B(n_211),
.C(n_213),
.Y(n_2888)
);

NAND3xp33_ASAP7_75t_SL g2889 ( 
.A(n_2860),
.B(n_214),
.C(n_215),
.Y(n_2889)
);

NOR3x1_ASAP7_75t_L g2890 ( 
.A(n_2862),
.B(n_215),
.C(n_216),
.Y(n_2890)
);

OAI21xp5_ASAP7_75t_L g2891 ( 
.A1(n_2857),
.A2(n_219),
.B(n_218),
.Y(n_2891)
);

NAND3xp33_ASAP7_75t_SL g2892 ( 
.A(n_2857),
.B(n_216),
.C(n_218),
.Y(n_2892)
);

AOI21xp5_ASAP7_75t_L g2893 ( 
.A1(n_2869),
.A2(n_220),
.B(n_221),
.Y(n_2893)
);

OAI221xp5_ASAP7_75t_L g2894 ( 
.A1(n_2857),
.A2(n_223),
.B1(n_220),
.B2(n_222),
.C(n_224),
.Y(n_2894)
);

INVx2_ASAP7_75t_L g2895 ( 
.A(n_2874),
.Y(n_2895)
);

NAND3xp33_ASAP7_75t_SL g2896 ( 
.A(n_2857),
.B(n_222),
.C(n_223),
.Y(n_2896)
);

AND2x2_ASAP7_75t_L g2897 ( 
.A(n_2863),
.B(n_225),
.Y(n_2897)
);

NAND4xp25_ASAP7_75t_L g2898 ( 
.A(n_2870),
.B(n_227),
.C(n_225),
.D(n_226),
.Y(n_2898)
);

OAI21xp5_ASAP7_75t_SL g2899 ( 
.A1(n_2857),
.A2(n_226),
.B(n_227),
.Y(n_2899)
);

NOR2xp67_ASAP7_75t_L g2900 ( 
.A(n_2857),
.B(n_229),
.Y(n_2900)
);

OAI211xp5_ASAP7_75t_L g2901 ( 
.A1(n_2857),
.A2(n_231),
.B(n_228),
.C(n_230),
.Y(n_2901)
);

NOR2xp33_ASAP7_75t_SL g2902 ( 
.A(n_2855),
.B(n_228),
.Y(n_2902)
);

NOR2xp33_ASAP7_75t_L g2903 ( 
.A(n_2857),
.B(n_230),
.Y(n_2903)
);

NOR2xp67_ASAP7_75t_SL g2904 ( 
.A(n_2857),
.B(n_231),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_SL g2905 ( 
.A(n_2857),
.B(n_232),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2874),
.Y(n_2906)
);

AOI221xp5_ASAP7_75t_SL g2907 ( 
.A1(n_2857),
.A2(n_234),
.B1(n_232),
.B2(n_233),
.C(n_235),
.Y(n_2907)
);

NAND4xp25_ASAP7_75t_L g2908 ( 
.A(n_2870),
.B(n_237),
.C(n_234),
.D(n_236),
.Y(n_2908)
);

NAND3x1_ASAP7_75t_L g2909 ( 
.A(n_2863),
.B(n_236),
.C(n_237),
.Y(n_2909)
);

NAND3xp33_ASAP7_75t_L g2910 ( 
.A(n_2866),
.B(n_238),
.C(n_239),
.Y(n_2910)
);

NOR2x1_ASAP7_75t_L g2911 ( 
.A(n_2874),
.B(n_238),
.Y(n_2911)
);

O2A1O1Ixp33_ASAP7_75t_L g2912 ( 
.A1(n_2857),
.A2(n_242),
.B(n_240),
.C(n_241),
.Y(n_2912)
);

NAND5xp2_ASAP7_75t_L g2913 ( 
.A(n_2857),
.B(n_242),
.C(n_240),
.D(n_241),
.E(n_243),
.Y(n_2913)
);

NAND4xp25_ASAP7_75t_L g2914 ( 
.A(n_2870),
.B(n_245),
.C(n_243),
.D(n_244),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2900),
.B(n_2897),
.Y(n_2915)
);

A2O1A1Ixp33_ASAP7_75t_L g2916 ( 
.A1(n_2912),
.A2(n_246),
.B(n_244),
.C(n_245),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2909),
.Y(n_2917)
);

NOR2x1_ASAP7_75t_L g2918 ( 
.A(n_2911),
.B(n_246),
.Y(n_2918)
);

NOR2x1_ASAP7_75t_L g2919 ( 
.A(n_2892),
.B(n_247),
.Y(n_2919)
);

NOR3x1_ASAP7_75t_L g2920 ( 
.A(n_2876),
.B(n_247),
.C(n_248),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_SL g2921 ( 
.A(n_2883),
.B(n_248),
.Y(n_2921)
);

INVxp67_ASAP7_75t_L g2922 ( 
.A(n_2913),
.Y(n_2922)
);

AND2x4_ASAP7_75t_L g2923 ( 
.A(n_2880),
.B(n_249),
.Y(n_2923)
);

NOR3xp33_ASAP7_75t_L g2924 ( 
.A(n_2882),
.B(n_249),
.C(n_250),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2904),
.Y(n_2925)
);

AOI22xp5_ASAP7_75t_L g2926 ( 
.A1(n_2884),
.A2(n_252),
.B1(n_250),
.B2(n_251),
.Y(n_2926)
);

NOR2x1_ASAP7_75t_L g2927 ( 
.A(n_2896),
.B(n_252),
.Y(n_2927)
);

AOI221x1_ASAP7_75t_L g2928 ( 
.A1(n_2887),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.C(n_256),
.Y(n_2928)
);

OAI21xp5_ASAP7_75t_SL g2929 ( 
.A1(n_2910),
.A2(n_2889),
.B(n_2879),
.Y(n_2929)
);

AND2x2_ASAP7_75t_L g2930 ( 
.A(n_2895),
.B(n_256),
.Y(n_2930)
);

NOR2xp67_ASAP7_75t_L g2931 ( 
.A(n_2885),
.B(n_257),
.Y(n_2931)
);

NAND2xp33_ASAP7_75t_L g2932 ( 
.A(n_2886),
.B(n_258),
.Y(n_2932)
);

OAI322xp33_ASAP7_75t_L g2933 ( 
.A1(n_2881),
.A2(n_263),
.A3(n_262),
.B1(n_260),
.B2(n_258),
.C1(n_259),
.C2(n_261),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2877),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2903),
.Y(n_2935)
);

NOR2x1p5_ASAP7_75t_L g2936 ( 
.A(n_2914),
.B(n_259),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2890),
.Y(n_2937)
);

OAI322xp33_ASAP7_75t_L g2938 ( 
.A1(n_2893),
.A2(n_266),
.A3(n_265),
.B1(n_262),
.B2(n_260),
.C1(n_261),
.C2(n_264),
.Y(n_2938)
);

AOI22xp33_ASAP7_75t_L g2939 ( 
.A1(n_2906),
.A2(n_265),
.B1(n_848),
.B2(n_847),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_SL g2940 ( 
.A(n_2907),
.B(n_2902),
.Y(n_2940)
);

XNOR2x1_ASAP7_75t_L g2941 ( 
.A(n_2891),
.B(n_343),
.Y(n_2941)
);

OAI322xp33_ASAP7_75t_L g2942 ( 
.A1(n_2878),
.A2(n_351),
.A3(n_349),
.B1(n_346),
.B2(n_344),
.C1(n_345),
.C2(n_347),
.Y(n_2942)
);

AOI22x1_ASAP7_75t_L g2943 ( 
.A1(n_2888),
.A2(n_356),
.B1(n_353),
.B2(n_355),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_L g2944 ( 
.A(n_2899),
.B(n_357),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2901),
.Y(n_2945)
);

INVx2_ASAP7_75t_L g2946 ( 
.A(n_2905),
.Y(n_2946)
);

AND2x2_ASAP7_75t_L g2947 ( 
.A(n_2898),
.B(n_358),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2908),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_L g2949 ( 
.A(n_2894),
.B(n_359),
.Y(n_2949)
);

OAI211xp5_ASAP7_75t_L g2950 ( 
.A1(n_2882),
.A2(n_362),
.B(n_360),
.C(n_361),
.Y(n_2950)
);

HB1xp67_ASAP7_75t_L g2951 ( 
.A(n_2900),
.Y(n_2951)
);

NAND4xp25_ASAP7_75t_SL g2952 ( 
.A(n_2876),
.B(n_368),
.C(n_365),
.D(n_366),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2909),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_L g2954 ( 
.A(n_2900),
.B(n_369),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2909),
.Y(n_2955)
);

NOR2x1_ASAP7_75t_L g2956 ( 
.A(n_2900),
.B(n_370),
.Y(n_2956)
);

OR2x2_ASAP7_75t_L g2957 ( 
.A(n_2917),
.B(n_2953),
.Y(n_2957)
);

NOR2xp67_ASAP7_75t_L g2958 ( 
.A(n_2955),
.B(n_371),
.Y(n_2958)
);

INVxp67_ASAP7_75t_SL g2959 ( 
.A(n_2918),
.Y(n_2959)
);

NAND3xp33_ASAP7_75t_SL g2960 ( 
.A(n_2924),
.B(n_373),
.C(n_375),
.Y(n_2960)
);

NAND3x1_ASAP7_75t_SL g2961 ( 
.A(n_2956),
.B(n_376),
.C(n_377),
.Y(n_2961)
);

NOR2xp33_ASAP7_75t_L g2962 ( 
.A(n_2922),
.B(n_378),
.Y(n_2962)
);

NOR2xp67_ASAP7_75t_L g2963 ( 
.A(n_2951),
.B(n_379),
.Y(n_2963)
);

XNOR2xp5_ASAP7_75t_L g2964 ( 
.A(n_2936),
.B(n_381),
.Y(n_2964)
);

NOR2x1_ASAP7_75t_L g2965 ( 
.A(n_2915),
.B(n_382),
.Y(n_2965)
);

NOR2x1_ASAP7_75t_SL g2966 ( 
.A(n_2921),
.B(n_383),
.Y(n_2966)
);

AND4x2_ASAP7_75t_L g2967 ( 
.A(n_2919),
.B(n_2927),
.C(n_2920),
.D(n_2929),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2923),
.Y(n_2968)
);

NAND2xp5_ASAP7_75t_L g2969 ( 
.A(n_2923),
.B(n_386),
.Y(n_2969)
);

OAI21xp5_ASAP7_75t_L g2970 ( 
.A1(n_2931),
.A2(n_387),
.B(n_388),
.Y(n_2970)
);

NOR4xp75_ASAP7_75t_L g2971 ( 
.A(n_2940),
.B(n_392),
.C(n_389),
.D(n_390),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_2930),
.Y(n_2972)
);

AND3x2_ASAP7_75t_L g2973 ( 
.A(n_2925),
.B(n_393),
.C(n_394),
.Y(n_2973)
);

NOR3x1_ASAP7_75t_L g2974 ( 
.A(n_2950),
.B(n_395),
.C(n_397),
.Y(n_2974)
);

NAND4xp75_ASAP7_75t_L g2975 ( 
.A(n_2928),
.B(n_2945),
.C(n_2937),
.D(n_2948),
.Y(n_2975)
);

NAND3xp33_ASAP7_75t_SL g2976 ( 
.A(n_2916),
.B(n_399),
.C(n_400),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2954),
.Y(n_2977)
);

NOR3xp33_ASAP7_75t_L g2978 ( 
.A(n_2949),
.B(n_401),
.C(n_402),
.Y(n_2978)
);

OR2x2_ASAP7_75t_L g2979 ( 
.A(n_2944),
.B(n_841),
.Y(n_2979)
);

INVx2_ASAP7_75t_L g2980 ( 
.A(n_2943),
.Y(n_2980)
);

INVx2_ASAP7_75t_SL g2981 ( 
.A(n_2946),
.Y(n_2981)
);

NAND3xp33_ASAP7_75t_L g2982 ( 
.A(n_2932),
.B(n_403),
.C(n_404),
.Y(n_2982)
);

NAND3xp33_ASAP7_75t_SL g2983 ( 
.A(n_2934),
.B(n_410),
.C(n_411),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2933),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2947),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2938),
.Y(n_2986)
);

NOR2x1p5_ASAP7_75t_L g2987 ( 
.A(n_2935),
.B(n_412),
.Y(n_2987)
);

INVx1_ASAP7_75t_SL g2988 ( 
.A(n_2941),
.Y(n_2988)
);

NOR2x1_ASAP7_75t_L g2989 ( 
.A(n_2952),
.B(n_415),
.Y(n_2989)
);

NOR2xp67_ASAP7_75t_L g2990 ( 
.A(n_2926),
.B(n_416),
.Y(n_2990)
);

AND2x2_ASAP7_75t_L g2991 ( 
.A(n_2939),
.B(n_417),
.Y(n_2991)
);

NOR2xp67_ASAP7_75t_L g2992 ( 
.A(n_2942),
.B(n_419),
.Y(n_2992)
);

NAND4xp25_ASAP7_75t_L g2993 ( 
.A(n_2924),
.B(n_422),
.C(n_420),
.D(n_421),
.Y(n_2993)
);

NOR3xp33_ASAP7_75t_L g2994 ( 
.A(n_2929),
.B(n_423),
.C(n_424),
.Y(n_2994)
);

NOR2x1_ASAP7_75t_L g2995 ( 
.A(n_2918),
.B(n_427),
.Y(n_2995)
);

NOR2x1p5_ASAP7_75t_L g2996 ( 
.A(n_2915),
.B(n_428),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2923),
.B(n_429),
.Y(n_2997)
);

NOR2x1_ASAP7_75t_L g2998 ( 
.A(n_2918),
.B(n_430),
.Y(n_2998)
);

NAND3xp33_ASAP7_75t_L g2999 ( 
.A(n_2928),
.B(n_431),
.C(n_433),
.Y(n_2999)
);

AND2x4_ASAP7_75t_L g3000 ( 
.A(n_2956),
.B(n_434),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2918),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2918),
.Y(n_3002)
);

NOR2x1_ASAP7_75t_L g3003 ( 
.A(n_2918),
.B(n_435),
.Y(n_3003)
);

NAND4xp75_ASAP7_75t_L g3004 ( 
.A(n_2918),
.B(n_442),
.C(n_436),
.D(n_441),
.Y(n_3004)
);

AOI21xp5_ASAP7_75t_SL g3005 ( 
.A1(n_2928),
.A2(n_838),
.B(n_835),
.Y(n_3005)
);

NAND3xp33_ASAP7_75t_SL g3006 ( 
.A(n_2953),
.B(n_443),
.C(n_444),
.Y(n_3006)
);

NAND3x1_ASAP7_75t_L g3007 ( 
.A(n_2918),
.B(n_445),
.C(n_446),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2968),
.Y(n_3008)
);

CKINVDCx5p33_ASAP7_75t_R g3009 ( 
.A(n_2981),
.Y(n_3009)
);

OAI21xp5_ASAP7_75t_L g3010 ( 
.A1(n_3007),
.A2(n_447),
.B(n_448),
.Y(n_3010)
);

INVx2_ASAP7_75t_L g3011 ( 
.A(n_2973),
.Y(n_3011)
);

NOR3xp33_ASAP7_75t_SL g3012 ( 
.A(n_2975),
.B(n_449),
.C(n_450),
.Y(n_3012)
);

OR2x2_ASAP7_75t_L g3013 ( 
.A(n_3001),
.B(n_451),
.Y(n_3013)
);

OR2x6_ASAP7_75t_L g3014 ( 
.A(n_3002),
.B(n_851),
.Y(n_3014)
);

OAI22xp5_ASAP7_75t_L g3015 ( 
.A1(n_2957),
.A2(n_457),
.B1(n_454),
.B2(n_456),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2959),
.Y(n_3016)
);

NOR2xp67_ASAP7_75t_L g3017 ( 
.A(n_2999),
.B(n_459),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2995),
.Y(n_3018)
);

INVx2_ASAP7_75t_SL g3019 ( 
.A(n_2998),
.Y(n_3019)
);

AOI22xp5_ASAP7_75t_L g3020 ( 
.A1(n_2962),
.A2(n_461),
.B1(n_458),
.B2(n_460),
.Y(n_3020)
);

NAND2x1p5_ASAP7_75t_L g3021 ( 
.A(n_3003),
.B(n_462),
.Y(n_3021)
);

OAI22xp5_ASAP7_75t_L g3022 ( 
.A1(n_2986),
.A2(n_465),
.B1(n_463),
.B2(n_464),
.Y(n_3022)
);

CKINVDCx5p33_ASAP7_75t_R g3023 ( 
.A(n_2972),
.Y(n_3023)
);

OAI21xp5_ASAP7_75t_L g3024 ( 
.A1(n_3005),
.A2(n_466),
.B(n_467),
.Y(n_3024)
);

AOI211xp5_ASAP7_75t_L g3025 ( 
.A1(n_3006),
.A2(n_473),
.B(n_469),
.C(n_471),
.Y(n_3025)
);

OR2x2_ASAP7_75t_L g3026 ( 
.A(n_2969),
.B(n_475),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_SL g3027 ( 
.A(n_3000),
.B(n_476),
.Y(n_3027)
);

NOR2xp67_ASAP7_75t_SL g3028 ( 
.A(n_3004),
.B(n_478),
.Y(n_3028)
);

NAND4xp75_ASAP7_75t_L g3029 ( 
.A(n_2965),
.B(n_482),
.C(n_479),
.D(n_481),
.Y(n_3029)
);

OAI21xp5_ASAP7_75t_L g3030 ( 
.A1(n_2958),
.A2(n_485),
.B(n_486),
.Y(n_3030)
);

INVx2_ASAP7_75t_L g3031 ( 
.A(n_2987),
.Y(n_3031)
);

NOR2xp33_ASAP7_75t_L g3032 ( 
.A(n_2997),
.B(n_2984),
.Y(n_3032)
);

INVx2_ASAP7_75t_L g3033 ( 
.A(n_3000),
.Y(n_3033)
);

NAND2xp33_ASAP7_75t_SL g3034 ( 
.A(n_2996),
.B(n_487),
.Y(n_3034)
);

INVx2_ASAP7_75t_SL g3035 ( 
.A(n_2989),
.Y(n_3035)
);

NOR2x1_ASAP7_75t_L g3036 ( 
.A(n_2963),
.B(n_488),
.Y(n_3036)
);

NAND3x1_ASAP7_75t_SL g3037 ( 
.A(n_2970),
.B(n_489),
.C(n_491),
.Y(n_3037)
);

INVx2_ASAP7_75t_L g3038 ( 
.A(n_2979),
.Y(n_3038)
);

AOI22xp5_ASAP7_75t_L g3039 ( 
.A1(n_2994),
.A2(n_497),
.B1(n_492),
.B2(n_494),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_SL g3040 ( 
.A(n_2980),
.B(n_499),
.Y(n_3040)
);

AND2x2_ASAP7_75t_L g3041 ( 
.A(n_2966),
.B(n_500),
.Y(n_3041)
);

AOI211xp5_ASAP7_75t_L g3042 ( 
.A1(n_2960),
.A2(n_506),
.B(n_501),
.C(n_502),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2967),
.Y(n_3043)
);

NAND4xp75_ASAP7_75t_L g3044 ( 
.A(n_2990),
.B(n_509),
.C(n_507),
.D(n_508),
.Y(n_3044)
);

NOR3xp33_ASAP7_75t_L g3045 ( 
.A(n_2961),
.B(n_510),
.C(n_511),
.Y(n_3045)
);

AOI22xp5_ASAP7_75t_L g3046 ( 
.A1(n_2978),
.A2(n_514),
.B1(n_512),
.B2(n_513),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2964),
.Y(n_3047)
);

AND3x2_ASAP7_75t_L g3048 ( 
.A(n_2985),
.B(n_528),
.C(n_516),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2991),
.B(n_517),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_L g3050 ( 
.A(n_2992),
.B(n_518),
.Y(n_3050)
);

AND2x4_ASAP7_75t_L g3051 ( 
.A(n_3008),
.B(n_2971),
.Y(n_3051)
);

NAND2xp5_ASAP7_75t_L g3052 ( 
.A(n_3009),
.B(n_2977),
.Y(n_3052)
);

INVxp33_ASAP7_75t_L g3053 ( 
.A(n_3036),
.Y(n_3053)
);

INVx2_ASAP7_75t_L g3054 ( 
.A(n_3048),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_3021),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_3013),
.Y(n_3056)
);

INVx2_ASAP7_75t_L g3057 ( 
.A(n_3014),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_3026),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_3016),
.Y(n_3059)
);

AND3x4_ASAP7_75t_L g3060 ( 
.A(n_3045),
.B(n_2974),
.C(n_2988),
.Y(n_3060)
);

XNOR2x1_ASAP7_75t_L g3061 ( 
.A(n_3023),
.B(n_3043),
.Y(n_3061)
);

NOR2x1_ASAP7_75t_L g3062 ( 
.A(n_3018),
.B(n_2982),
.Y(n_3062)
);

OA22x2_ASAP7_75t_L g3063 ( 
.A1(n_3024),
.A2(n_2976),
.B1(n_2993),
.B2(n_2983),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_3011),
.Y(n_3064)
);

NAND4xp75_ASAP7_75t_L g3065 ( 
.A(n_3012),
.B(n_852),
.C(n_523),
.D(n_521),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_3049),
.Y(n_3066)
);

INVx2_ASAP7_75t_SL g3067 ( 
.A(n_3041),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_SL g3068 ( 
.A(n_3019),
.B(n_3035),
.Y(n_3068)
);

AND2x2_ASAP7_75t_L g3069 ( 
.A(n_3033),
.B(n_522),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_3014),
.Y(n_3070)
);

NOR2x1_ASAP7_75t_L g3071 ( 
.A(n_3029),
.B(n_525),
.Y(n_3071)
);

NOR2x1p5_ASAP7_75t_L g3072 ( 
.A(n_3044),
.B(n_527),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_3027),
.Y(n_3073)
);

AOI22xp5_ASAP7_75t_L g3074 ( 
.A1(n_3032),
.A2(n_531),
.B1(n_529),
.B2(n_530),
.Y(n_3074)
);

XNOR2x1_ASAP7_75t_L g3075 ( 
.A(n_3017),
.B(n_535),
.Y(n_3075)
);

AOI211xp5_ASAP7_75t_L g3076 ( 
.A1(n_3022),
.A2(n_539),
.B(n_536),
.C(n_538),
.Y(n_3076)
);

BUFx12f_ASAP7_75t_L g3077 ( 
.A(n_3034),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_SL g3078 ( 
.A(n_3010),
.B(n_540),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_3050),
.Y(n_3079)
);

OAI22xp33_ASAP7_75t_SL g3080 ( 
.A1(n_3040),
.A2(n_544),
.B1(n_542),
.B2(n_543),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_3031),
.Y(n_3081)
);

AND2x2_ASAP7_75t_L g3082 ( 
.A(n_3038),
.B(n_545),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_3028),
.B(n_3030),
.Y(n_3083)
);

NOR3xp33_ASAP7_75t_L g3084 ( 
.A(n_3047),
.B(n_546),
.C(n_548),
.Y(n_3084)
);

AND2x4_ASAP7_75t_L g3085 ( 
.A(n_3046),
.B(n_850),
.Y(n_3085)
);

AND2x4_ASAP7_75t_L g3086 ( 
.A(n_3039),
.B(n_549),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_L g3087 ( 
.A(n_3069),
.B(n_3082),
.Y(n_3087)
);

AOI311xp33_ASAP7_75t_L g3088 ( 
.A1(n_3064),
.A2(n_3059),
.A3(n_3081),
.B(n_3073),
.C(n_3056),
.Y(n_3088)
);

AND2x4_ASAP7_75t_L g3089 ( 
.A(n_3054),
.B(n_3072),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_SL g3090 ( 
.A(n_3080),
.B(n_3025),
.Y(n_3090)
);

BUFx3_ASAP7_75t_L g3091 ( 
.A(n_3077),
.Y(n_3091)
);

XNOR2xp5_ASAP7_75t_L g3092 ( 
.A(n_3061),
.B(n_3037),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_3067),
.B(n_3042),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_3068),
.Y(n_3094)
);

OAI22x1_ASAP7_75t_L g3095 ( 
.A1(n_3060),
.A2(n_3020),
.B1(n_3015),
.B2(n_555),
.Y(n_3095)
);

AOI211xp5_ASAP7_75t_SL g3096 ( 
.A1(n_3052),
.A2(n_556),
.B(n_550),
.C(n_551),
.Y(n_3096)
);

NOR3xp33_ASAP7_75t_L g3097 ( 
.A(n_3062),
.B(n_557),
.C(n_558),
.Y(n_3097)
);

INVxp33_ASAP7_75t_SL g3098 ( 
.A(n_3055),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_3051),
.Y(n_3099)
);

XOR2x1_ASAP7_75t_L g3100 ( 
.A(n_3075),
.B(n_560),
.Y(n_3100)
);

AOI22xp33_ASAP7_75t_L g3101 ( 
.A1(n_3086),
.A2(n_565),
.B1(n_562),
.B2(n_564),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_3063),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_3071),
.Y(n_3103)
);

AOI211xp5_ASAP7_75t_L g3104 ( 
.A1(n_3053),
.A2(n_569),
.B(n_567),
.C(n_568),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_3057),
.Y(n_3105)
);

BUFx2_ASAP7_75t_L g3106 ( 
.A(n_3070),
.Y(n_3106)
);

AOI21xp5_ASAP7_75t_L g3107 ( 
.A1(n_3078),
.A2(n_571),
.B(n_573),
.Y(n_3107)
);

AND2x2_ASAP7_75t_L g3108 ( 
.A(n_3058),
.B(n_574),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_3083),
.Y(n_3109)
);

NOR2x1p5_ASAP7_75t_L g3110 ( 
.A(n_3065),
.B(n_577),
.Y(n_3110)
);

OAI211xp5_ASAP7_75t_L g3111 ( 
.A1(n_3076),
.A2(n_581),
.B(n_579),
.C(n_580),
.Y(n_3111)
);

INVx3_ASAP7_75t_L g3112 ( 
.A(n_3085),
.Y(n_3112)
);

OAI22xp33_ASAP7_75t_L g3113 ( 
.A1(n_3079),
.A2(n_588),
.B1(n_583),
.B2(n_584),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_3066),
.Y(n_3114)
);

OR2x2_ASAP7_75t_L g3115 ( 
.A(n_3094),
.B(n_3084),
.Y(n_3115)
);

AOI211xp5_ASAP7_75t_L g3116 ( 
.A1(n_3111),
.A2(n_3074),
.B(n_595),
.C(n_591),
.Y(n_3116)
);

AOI22xp33_ASAP7_75t_L g3117 ( 
.A1(n_3098),
.A2(n_597),
.B1(n_593),
.B2(n_596),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_3106),
.Y(n_3118)
);

BUFx12f_ASAP7_75t_L g3119 ( 
.A(n_3091),
.Y(n_3119)
);

NAND4xp75_ASAP7_75t_L g3120 ( 
.A(n_3102),
.B(n_601),
.C(n_599),
.D(n_600),
.Y(n_3120)
);

NAND4xp75_ASAP7_75t_L g3121 ( 
.A(n_3105),
.B(n_605),
.C(n_602),
.D(n_604),
.Y(n_3121)
);

NAND4xp75_ASAP7_75t_L g3122 ( 
.A(n_3099),
.B(n_609),
.C(n_606),
.D(n_607),
.Y(n_3122)
);

OAI31xp33_ASAP7_75t_SL g3123 ( 
.A1(n_3100),
.A2(n_613),
.A3(n_610),
.B(n_612),
.Y(n_3123)
);

AOI211xp5_ASAP7_75t_L g3124 ( 
.A1(n_3103),
.A2(n_618),
.B(n_614),
.C(n_617),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_3087),
.Y(n_3125)
);

NAND3xp33_ASAP7_75t_L g3126 ( 
.A(n_3088),
.B(n_621),
.C(n_622),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_3108),
.B(n_623),
.Y(n_3127)
);

XNOR2x1_ASAP7_75t_L g3128 ( 
.A(n_3118),
.B(n_3092),
.Y(n_3128)
);

AOI211xp5_ASAP7_75t_L g3129 ( 
.A1(n_3126),
.A2(n_3107),
.B(n_3109),
.C(n_3114),
.Y(n_3129)
);

OR4x1_ASAP7_75t_L g3130 ( 
.A(n_3125),
.B(n_3119),
.C(n_3123),
.D(n_3089),
.Y(n_3130)
);

NAND4xp25_ASAP7_75t_L g3131 ( 
.A(n_3116),
.B(n_3093),
.C(n_3089),
.D(n_3090),
.Y(n_3131)
);

OAI321xp33_ASAP7_75t_L g3132 ( 
.A1(n_3115),
.A2(n_3101),
.A3(n_3113),
.B1(n_3104),
.B2(n_3095),
.C(n_3110),
.Y(n_3132)
);

OAI221xp5_ASAP7_75t_L g3133 ( 
.A1(n_3127),
.A2(n_3097),
.B1(n_3112),
.B2(n_3096),
.C(n_627),
.Y(n_3133)
);

AOI321xp33_ASAP7_75t_L g3134 ( 
.A1(n_3124),
.A2(n_628),
.A3(n_630),
.B1(n_625),
.B2(n_626),
.C(n_629),
.Y(n_3134)
);

NOR3xp33_ASAP7_75t_L g3135 ( 
.A(n_3120),
.B(n_631),
.C(n_632),
.Y(n_3135)
);

AOI211xp5_ASAP7_75t_L g3136 ( 
.A1(n_3122),
.A2(n_636),
.B(n_633),
.C(n_634),
.Y(n_3136)
);

NOR2x1_ASAP7_75t_L g3137 ( 
.A(n_3121),
.B(n_637),
.Y(n_3137)
);

NOR3xp33_ASAP7_75t_L g3138 ( 
.A(n_3117),
.B(n_639),
.C(n_640),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_3137),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_3128),
.Y(n_3140)
);

INVx1_ASAP7_75t_SL g3141 ( 
.A(n_3130),
.Y(n_3141)
);

INVxp67_ASAP7_75t_L g3142 ( 
.A(n_3133),
.Y(n_3142)
);

AOI22xp33_ASAP7_75t_L g3143 ( 
.A1(n_3135),
.A2(n_645),
.B1(n_642),
.B2(n_644),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_3129),
.Y(n_3144)
);

OA22x2_ASAP7_75t_L g3145 ( 
.A1(n_3132),
.A2(n_648),
.B1(n_646),
.B2(n_647),
.Y(n_3145)
);

OAI21xp5_ASAP7_75t_L g3146 ( 
.A1(n_3138),
.A2(n_649),
.B(n_651),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_L g3147 ( 
.A(n_3136),
.B(n_653),
.Y(n_3147)
);

OAI222xp33_ASAP7_75t_L g3148 ( 
.A1(n_3141),
.A2(n_3131),
.B1(n_3134),
.B2(n_657),
.C1(n_660),
.C2(n_655),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_L g3149 ( 
.A(n_3140),
.B(n_656),
.Y(n_3149)
);

XNOR2xp5_ASAP7_75t_L g3150 ( 
.A(n_3144),
.B(n_659),
.Y(n_3150)
);

NOR4xp25_ASAP7_75t_L g3151 ( 
.A(n_3139),
.B(n_663),
.C(n_661),
.D(n_662),
.Y(n_3151)
);

XNOR2xp5_ASAP7_75t_L g3152 ( 
.A(n_3145),
.B(n_664),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_L g3153 ( 
.A(n_3147),
.B(n_665),
.Y(n_3153)
);

OR4x1_ASAP7_75t_L g3154 ( 
.A(n_3142),
.B(n_669),
.C(n_666),
.D(n_668),
.Y(n_3154)
);

OAI322xp33_ASAP7_75t_L g3155 ( 
.A1(n_3146),
.A2(n_678),
.A3(n_675),
.B1(n_672),
.B2(n_670),
.C1(n_671),
.C2(n_674),
.Y(n_3155)
);

A2O1A1Ixp33_ASAP7_75t_L g3156 ( 
.A1(n_3143),
.A2(n_682),
.B(n_679),
.C(n_680),
.Y(n_3156)
);

AOI22xp5_ASAP7_75t_L g3157 ( 
.A1(n_3152),
.A2(n_686),
.B1(n_683),
.B2(n_685),
.Y(n_3157)
);

OAI22xp33_ASAP7_75t_L g3158 ( 
.A1(n_3149),
.A2(n_691),
.B1(n_687),
.B2(n_689),
.Y(n_3158)
);

OAI22xp5_ASAP7_75t_SL g3159 ( 
.A1(n_3154),
.A2(n_695),
.B1(n_692),
.B2(n_694),
.Y(n_3159)
);

OAI22xp5_ASAP7_75t_SL g3160 ( 
.A1(n_3153),
.A2(n_698),
.B1(n_696),
.B2(n_697),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_3150),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_3156),
.Y(n_3162)
);

AO21x2_ASAP7_75t_L g3163 ( 
.A1(n_3161),
.A2(n_3148),
.B(n_3151),
.Y(n_3163)
);

XNOR2x1_ASAP7_75t_L g3164 ( 
.A(n_3157),
.B(n_3155),
.Y(n_3164)
);

AOI21xp5_ASAP7_75t_L g3165 ( 
.A1(n_3162),
.A2(n_700),
.B(n_701),
.Y(n_3165)
);

OAI21xp5_ASAP7_75t_L g3166 ( 
.A1(n_3164),
.A2(n_3158),
.B(n_3159),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_3163),
.Y(n_3167)
);

INVxp67_ASAP7_75t_SL g3168 ( 
.A(n_3167),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_3166),
.Y(n_3169)
);

OR2x6_ASAP7_75t_L g3170 ( 
.A(n_3169),
.B(n_3165),
.Y(n_3170)
);

AOI21xp33_ASAP7_75t_L g3171 ( 
.A1(n_3170),
.A2(n_3168),
.B(n_3160),
.Y(n_3171)
);

AOI21xp5_ASAP7_75t_L g3172 ( 
.A1(n_3171),
.A2(n_702),
.B(n_704),
.Y(n_3172)
);


endmodule