module real_jpeg_33927_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_0),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g213 ( 
.A(n_0),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_0),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_0),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_1),
.B(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_1),
.B(n_169),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_3),
.A2(n_69),
.B1(n_75),
.B2(n_76),
.Y(n_68)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_3),
.A2(n_75),
.B1(n_276),
.B2(n_278),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_3),
.A2(n_75),
.B1(n_426),
.B2(n_431),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_3),
.A2(n_75),
.B1(n_466),
.B2(n_470),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_4),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_4),
.Y(n_206)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_4),
.Y(n_218)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_4),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_5),
.Y(n_131)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_5),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_6),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_7),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_7),
.Y(n_108)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_7),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_7),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_9),
.A2(n_183),
.B1(n_184),
.B2(n_186),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_9),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_L g225 ( 
.A1(n_9),
.A2(n_105),
.B1(n_183),
.B2(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_9),
.A2(n_183),
.B1(n_290),
.B2(n_293),
.Y(n_289)
);

OAI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_9),
.A2(n_183),
.B1(n_364),
.B2(n_366),
.Y(n_363)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_10),
.Y(n_85)
);

OAI22x1_ASAP7_75t_SL g57 ( 
.A1(n_11),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_11),
.Y(n_61)
);

AO22x2_ASAP7_75t_SL g114 ( 
.A1(n_11),
.A2(n_61),
.B1(n_115),
.B2(n_118),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_11),
.A2(n_61),
.B1(n_215),
.B2(n_219),
.Y(n_214)
);

OAI22x1_ASAP7_75t_L g314 ( 
.A1(n_11),
.A2(n_61),
.B1(n_315),
.B2(n_317),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_12),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_12),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_13),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_13),
.A2(n_28),
.B1(n_103),
.B2(n_105),
.Y(n_102)
);

AOI22x1_ASAP7_75t_SL g153 ( 
.A1(n_13),
.A2(n_28),
.B1(n_154),
.B2(n_157),
.Y(n_153)
);

AO22x1_ASAP7_75t_SL g203 ( 
.A1(n_13),
.A2(n_28),
.B1(n_204),
.B2(n_207),
.Y(n_203)
);

NAND2xp33_ASAP7_75t_SL g240 ( 
.A(n_13),
.B(n_241),
.Y(n_240)
);

OAI32xp33_ASAP7_75t_L g326 ( 
.A1(n_13),
.A2(n_327),
.A3(n_333),
.B1(n_335),
.B2(n_339),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_13),
.B(n_151),
.Y(n_354)
);

OAI21xp33_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_171),
.B(n_548),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_168),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_16),
.B(n_169),
.Y(n_549)
);

OR2x2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_167),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_65),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_18),
.B(n_65),
.Y(n_167)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_45),
.Y(n_19)
);

INVxp33_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_21),
.B(n_409),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_32),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_22),
.B(n_48),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_22),
.A2(n_48),
.B(n_475),
.Y(n_474)
);

OAI21x1_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_28),
.B(n_29),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_27),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_27),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_30),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_28),
.B(n_33),
.Y(n_193)
);

AOI32xp33_ASAP7_75t_L g230 ( 
.A1(n_28),
.A2(n_231),
.A3(n_234),
.B1(n_239),
.B2(n_240),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_28),
.B(n_336),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_28),
.B(n_379),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_28),
.B(n_197),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_29),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_31),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_32),
.B(n_57),
.Y(n_161)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2x1p5_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_34),
.B(n_289),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_34),
.Y(n_475)
);

AO22x2_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_38),
.B1(n_40),
.B2(n_42),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_37),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_37),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_37),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g469 ( 
.A(n_37),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_39),
.Y(n_260)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_39),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_41),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_41),
.Y(n_271)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OA21x2_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_68),
.B(n_79),
.Y(n_67)
);

OA21x2_ASAP7_75t_SL g505 ( 
.A1(n_46),
.A2(n_68),
.B(n_79),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_47),
.B(n_288),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_57),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_48),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_48),
.B(n_289),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_53),
.B2(n_55),
.Y(n_49)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_159),
.C(n_162),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_66),
.B(n_517),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_80),
.C(n_109),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_68),
.A2(n_160),
.B(n_161),
.Y(n_159)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_80),
.B(n_284),
.Y(n_283)
);

MAJx2_ASAP7_75t_L g412 ( 
.A(n_80),
.B(n_284),
.C(n_286),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_80),
.A2(n_110),
.B(n_507),
.Y(n_506)
);

NOR3xp33_ASAP7_75t_L g507 ( 
.A(n_80),
.B(n_112),
.C(n_149),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_80),
.Y(n_514)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_80),
.Y(n_533)
);

OA21x2_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_92),
.B(n_102),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_81),
.B(n_102),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_81),
.B(n_225),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_81),
.B(n_314),
.Y(n_357)
);

INVxp33_ASAP7_75t_L g379 ( 
.A(n_81),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_81),
.B(n_425),
.Y(n_424)
);

AO22x2_ASAP7_75t_L g455 ( 
.A1(n_81),
.A2(n_92),
.B1(n_314),
.B2(n_425),
.Y(n_455)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_93),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_86),
.B1(n_89),
.B2(n_91),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_85),
.Y(n_347)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_87),
.Y(n_220)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_87),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_87),
.Y(n_338)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_88),
.Y(n_202)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_92),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_92),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_92),
.B(n_102),
.Y(n_350)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_97),
.B1(n_98),
.B2(n_100),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_96),
.Y(n_233)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_96),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_101),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_104),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_107),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_108),
.Y(n_228)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_148),
.Y(n_110)
);

NAND2x1_ASAP7_75t_L g462 ( 
.A(n_111),
.B(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_113),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_122),
.Y(n_113)
);

AND2x4_ASAP7_75t_L g191 ( 
.A(n_114),
.B(n_151),
.Y(n_191)
);

NAND2xp33_ASAP7_75t_L g513 ( 
.A(n_114),
.B(n_151),
.Y(n_513)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_117),
.Y(n_185)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_117),
.Y(n_256)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_122),
.B(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

NOR2x1_ASAP7_75t_L g309 ( 
.A(n_123),
.B(n_153),
.Y(n_309)
);

AO21x2_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_132),
.B(n_140),
.Y(n_123)
);

INVxp33_ASAP7_75t_L g239 ( 
.A(n_124),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_127),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_136),
.A2(n_141),
.B1(n_143),
.B2(n_145),
.Y(n_140)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_141),
.Y(n_342)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_142),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_150),
.B(n_181),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_151),
.B(n_182),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_151),
.B(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_153),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_159),
.A2(n_162),
.B1(n_163),
.B2(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_159),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_161),
.B(n_409),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_161),
.B(n_287),
.Y(n_508)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_163),
.B(n_438),
.C(n_439),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_164),
.B(n_438),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_166),
.A2(n_465),
.B(n_513),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_171),
.A2(n_549),
.B(n_550),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_500),
.B(n_543),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_490),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_399),
.B(n_489),
.Y(n_174)
);

AO21x1_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_296),
.B(n_398),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_248),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_177),
.B(n_248),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_222),
.C(n_229),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_178),
.A2(n_179),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_192),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_180),
.A2(n_221),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_190),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_191),
.Y(n_190)
);

NOR2x1p5_ASAP7_75t_SL g451 ( 
.A(n_191),
.B(n_309),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_194),
.B(n_221),
.Y(n_192)
);

NOR2x1_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_194),
.Y(n_221)
);

NAND2xp33_ASAP7_75t_SL g251 ( 
.A(n_193),
.B(n_194),
.Y(n_251)
);

NOR2x1p5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_209),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_195),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_203),
.Y(n_195)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_196),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_196),
.B(n_214),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_196),
.B(n_363),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_201),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_203),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_203),
.B(n_361),
.Y(n_360)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_206),
.Y(n_208)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp33_ASAP7_75t_SL g380 ( 
.A(n_210),
.B(n_362),
.Y(n_380)
);

OAI21xp33_ASAP7_75t_SL g414 ( 
.A1(n_210),
.A2(n_244),
.B(n_275),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_211),
.Y(n_274)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_218),
.Y(n_277)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_222),
.B(n_229),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_223),
.B(n_313),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_224),
.B(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

NOR2xp67_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_243),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_230),
.A2(n_243),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_230),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx6f_ASAP7_75t_SL g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_243),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_243),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_243),
.A2(n_304),
.B1(n_474),
.B2(n_476),
.Y(n_473)
);

AO21x2_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_245),
.B(n_247),
.Y(n_243)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_245),
.Y(n_361)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_282),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_250),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_252),
.B(n_282),
.C(n_442),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_273),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_253),
.B(n_273),
.Y(n_405)
);

OAI31xp33_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_257),
.A3(n_261),
.B(n_265),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_270),
.B(n_272),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx5_ASAP7_75t_L g470 ( 
.A(n_270),
.Y(n_470)
);

INVx8_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B(n_281),
.Y(n_273)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_277),
.Y(n_365)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_281),
.B(n_372),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_281),
.B(n_360),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_286),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_291),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_321),
.B(n_397),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_301),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_298),
.B(n_301),
.Y(n_397)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_306),
.C(n_310),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_303),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_303),
.B(n_393),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_304),
.A2(n_454),
.B1(n_455),
.B2(n_456),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_304),
.B(n_455),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_306),
.A2(n_307),
.B1(n_310),
.B2(n_311),
.Y(n_393)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_312),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_313),
.B(n_424),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_313),
.A2(n_422),
.B(n_424),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_320),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_391),
.B(n_396),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_323),
.A2(n_369),
.B(n_390),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_351),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_324),
.B(n_351),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_348),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_325),
.A2(n_326),
.B1(n_348),
.B2(n_349),
.Y(n_375)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_332),
.Y(n_368)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_343),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_350),
.B(n_357),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_358),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_353),
.A2(n_354),
.B1(n_355),
.B2(n_356),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_353),
.B(n_359),
.C(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_356),
.Y(n_395)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_362),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_363),
.B(n_373),
.Y(n_372)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_366),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

AOI21x1_ASAP7_75t_L g369 ( 
.A1(n_370),
.A2(n_376),
.B(n_389),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_375),
.Y(n_370)
);

NOR2xp67_ASAP7_75t_L g389 ( 
.A(n_371),
.B(n_375),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_372),
.B(n_383),
.Y(n_382)
);

BUFx4f_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_377),
.A2(n_381),
.B(n_388),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_380),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_378),
.B(n_380),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_382),
.B(n_384),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_387),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_394),
.Y(n_391)
);

NOR2xp67_ASAP7_75t_L g396 ( 
.A(n_392),
.B(n_394),
.Y(n_396)
);

NOR3xp33_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_445),
.C(n_482),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_440),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_401),
.B(n_493),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_416),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_402),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_412),
.C(n_413),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_403),
.B(n_444),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_406),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_405),
.B(n_411),
.C(n_420),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_407),
.A2(n_408),
.B1(n_410),
.B2(n_411),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_408),
.Y(n_420)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_410),
.Y(n_411)
);

XOR2x1_ASAP7_75t_SL g444 ( 
.A(n_412),
.B(n_413),
.Y(n_444)
);

XOR2x2_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_415),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_414),
.B(n_415),
.Y(n_439)
);

INVxp33_ASAP7_75t_L g496 ( 
.A(n_416),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_417),
.A2(n_418),
.B1(n_435),
.B2(n_436),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_421),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_419),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_421),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_427),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_435),
.B(n_484),
.C(n_486),
.Y(n_483)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_437),
.B(n_439),
.Y(n_436)
);

OR2x2_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_443),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_441),
.B(n_443),
.Y(n_493)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_445),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_459),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_446),
.B(n_459),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_453),
.C(n_457),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_448),
.B(n_453),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_450),
.Y(n_448)
);

INVxp33_ASAP7_75t_SL g480 ( 
.A(n_449),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_452),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_451),
.Y(n_481)
);

INVxp33_ASAP7_75t_SL g479 ( 
.A(n_452),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_454),
.A2(n_477),
.B(n_527),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_455),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_458),
.B(n_488),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_478),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_472),
.Y(n_460)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_461),
.Y(n_523)
);

XNOR2x1_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_471),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_462),
.B(n_471),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVxp33_ASAP7_75t_SL g522 ( 
.A(n_472),
.Y(n_522)
);

XNOR2x1_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_477),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g476 ( 
.A(n_474),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_474),
.Y(n_528)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_478),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_480),
.C(n_481),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_482),
.A2(n_492),
.B(n_494),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_487),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_483),
.B(n_487),
.Y(n_498)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_491),
.A2(n_497),
.B(n_499),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_496),
.Y(n_494)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_519),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_501),
.A2(n_544),
.B(n_547),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_516),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_502),
.B(n_516),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_508),
.C(n_509),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_504),
.A2(n_508),
.B1(n_515),
.B2(n_542),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_504),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_506),
.Y(n_504)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_508),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_508),
.A2(n_515),
.B1(n_532),
.B2(n_534),
.Y(n_531)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_510),
.B(n_541),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_514),
.C(n_515),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_512),
.B(n_533),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_537),
.Y(n_519)
);

NOR2xp67_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_525),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_521),
.B(n_525),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_523),
.C(n_524),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_526),
.B(n_529),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_526),
.B(n_535),
.C(n_539),
.Y(n_538)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_530),
.A2(n_531),
.B1(n_535),
.B2(n_536),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_531),
.Y(n_539)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_532),
.Y(n_534)
);

INVxp67_ASAP7_75t_SL g535 ( 
.A(n_536),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g544 ( 
.A1(n_537),
.A2(n_545),
.B(n_546),
.Y(n_544)
);

NOR2x1_ASAP7_75t_SL g537 ( 
.A(n_538),
.B(n_540),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_538),
.B(n_540),
.Y(n_546)
);


endmodule