module fake_ariane_3240_n_5976 (n_295, n_356, n_556, n_170, n_190, n_698, n_695, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_176, n_691, n_34, n_404, n_172, n_678, n_651, n_347, n_423, n_183, n_469, n_479, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_610, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_690, n_416, n_283, n_50, n_187, n_525, n_367, n_713, n_649, n_598, n_345, n_374, n_318, n_103, n_244, n_643, n_679, n_226, n_220, n_261, n_682, n_36, n_663, n_370, n_706, n_189, n_72, n_286, n_443, n_586, n_57, n_686, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_607, n_670, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_631, n_23, n_399, n_554, n_520, n_87, n_279, n_702, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_665, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_668, n_339, n_672, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_701, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_703, n_510, n_256, n_326, n_681, n_227, n_48, n_188, n_323, n_550, n_635, n_707, n_330, n_400, n_689, n_694, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_699, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_620, n_228, n_325, n_276, n_93, n_688, n_636, n_427, n_108, n_587, n_497, n_693, n_303, n_671, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_661, n_488, n_667, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_684, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_579, n_459, n_685, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_237, n_175, n_711, n_453, n_74, n_491, n_19, n_40, n_181, n_616, n_617, n_658, n_630, n_705, n_570, n_53, n_260, n_362, n_543, n_310, n_709, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_660, n_464, n_575, n_546, n_297, n_662, n_641, n_503, n_700, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_708, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_680, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_710, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_652, n_451, n_613, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_696, n_674, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_656, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_629, n_664, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_692, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_657, n_513, n_288, n_179, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_659, n_67, n_509, n_583, n_306, n_666, n_313, n_92, n_430, n_626, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_669, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_697, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_704, n_132, n_147, n_204, n_615, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_425, n_431, n_508, n_624, n_118, n_121, n_618, n_411, n_484, n_712, n_353, n_22, n_241, n_29, n_357, n_412, n_687, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_127, n_531, n_675, n_5976);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_698;
input n_695;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_176;
input n_691;
input n_34;
input n_404;
input n_172;
input n_678;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_690;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_713;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_706;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_686;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_702;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_665;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_668;
input n_339;
input n_672;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_701;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_703;
input n_510;
input n_256;
input n_326;
input n_681;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_707;
input n_330;
input n_400;
input n_689;
input n_694;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_699;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_693;
input n_303;
input n_671;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_661;
input n_488;
input n_667;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_685;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_237;
input n_175;
input n_711;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_616;
input n_617;
input n_658;
input n_630;
input n_705;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_709;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_660;
input n_464;
input n_575;
input n_546;
input n_297;
input n_662;
input n_641;
input n_503;
input n_700;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_708;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_710;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_652;
input n_451;
input n_613;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_696;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_692;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_657;
input n_513;
input n_288;
input n_179;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_659;
input n_67;
input n_509;
input n_583;
input n_306;
input n_666;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_669;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_697;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_704;
input n_132;
input n_147;
input n_204;
input n_615;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_425;
input n_431;
input n_508;
input n_624;
input n_118;
input n_121;
input n_618;
input n_411;
input n_484;
input n_712;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;
input n_675;

output n_5976;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_4030;
wire n_4770;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_2679;
wire n_5402;
wire n_2182;
wire n_5553;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_5717;
wire n_2993;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_4962;
wire n_1430;
wire n_2002;
wire n_1238;
wire n_2729;
wire n_4302;
wire n_5791;
wire n_4547;
wire n_5090;
wire n_3765;
wire n_864;
wire n_5302;
wire n_1096;
wire n_1379;
wire n_2376;
wire n_2790;
wire n_2207;
wire n_5712;
wire n_3954;
wire n_4982;
wire n_2042;
wire n_1131;
wire n_5479;
wire n_2646;
wire n_737;
wire n_2653;
wire n_4610;
wire n_3115;
wire n_4028;
wire n_5263;
wire n_5565;
wire n_2482;
wire n_1682;
wire n_958;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_5590;
wire n_2621;
wire n_4853;
wire n_1909;
wire n_5229;
wire n_4260;
wire n_903;
wire n_3348;
wire n_3261;
wire n_1761;
wire n_1690;
wire n_2807;
wire n_1018;
wire n_4512;
wire n_4132;
wire n_1364;
wire n_2390;
wire n_4500;
wire n_2322;
wire n_1107;
wire n_2663;
wire n_5481;
wire n_4824;
wire n_5340;
wire n_3545;
wire n_1428;
wire n_1284;
wire n_4741;
wire n_1241;
wire n_4143;
wire n_4273;
wire n_901;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_1519;
wire n_5896;
wire n_4567;
wire n_786;
wire n_5833;
wire n_3552;
wire n_2950;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_5589;
wire n_3015;
wire n_5744;
wire n_3870;
wire n_3749;
wire n_1676;
wire n_1085;
wire n_5691;
wire n_3482;
wire n_5403;
wire n_823;
wire n_1900;
wire n_4268;
wire n_863;
wire n_3960;
wire n_2433;
wire n_899;
wire n_3975;
wire n_5830;
wire n_2004;
wire n_4018;
wire n_1495;
wire n_3325;
wire n_4227;
wire n_5158;
wire n_5152;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_1924;
wire n_1811;
wire n_3612;
wire n_4505;
wire n_1840;
wire n_5247;
wire n_5464;
wire n_4476;
wire n_844;
wire n_1267;
wire n_2956;
wire n_5210;
wire n_2382;
wire n_1213;
wire n_780;
wire n_5292;
wire n_1918;
wire n_4119;
wire n_4443;
wire n_4000;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_1140;
wire n_3458;
wire n_5843;
wire n_3511;
wire n_2077;
wire n_1121;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_1216;
wire n_4908;
wire n_3754;
wire n_5060;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_5913;
wire n_4530;
wire n_1432;
wire n_2245;
wire n_5614;
wire n_5391;
wire n_5452;
wire n_3359;
wire n_3841;
wire n_5249;
wire n_851;
wire n_3900;
wire n_3413;
wire n_5076;
wire n_3539;
wire n_5757;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_930;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_5046;
wire n_1386;
wire n_3506;
wire n_4827;
wire n_1842;
wire n_4993;
wire n_3678;
wire n_2791;
wire n_1661;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_5968;
wire n_992;
wire n_966;
wire n_3549;
wire n_3914;
wire n_5586;
wire n_1692;
wire n_2611;
wire n_5468;
wire n_3029;
wire n_4745;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_5971;
wire n_5056;
wire n_1178;
wire n_2015;
wire n_5204;
wire n_2877;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_2161;
wire n_746;
wire n_1357;
wire n_1787;
wire n_1389;
wire n_3172;
wire n_2659;
wire n_4033;
wire n_3747;
wire n_4905;
wire n_4508;
wire n_5897;
wire n_4045;
wire n_4894;
wire n_3651;
wire n_1812;
wire n_3614;
wire n_959;
wire n_2257;
wire n_1101;
wire n_1343;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_5778;
wire n_5179;
wire n_2435;
wire n_5680;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_5685;
wire n_5974;
wire n_5723;
wire n_5922;
wire n_5549;
wire n_1087;
wire n_2388;
wire n_2273;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_3700;
wire n_4307;
wire n_2795;
wire n_1841;
wire n_1680;
wire n_2954;
wire n_4438;
wire n_974;
wire n_3814;
wire n_5831;
wire n_4367;
wire n_5134;
wire n_2467;
wire n_4195;
wire n_5091;
wire n_4866;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_5708;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_5454;
wire n_1209;
wire n_4254;
wire n_3438;
wire n_2625;
wire n_5373;
wire n_1578;
wire n_3147;
wire n_3661;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_1568;
wire n_2919;
wire n_3108;
wire n_5788;
wire n_2632;
wire n_5557;
wire n_4314;
wire n_2980;
wire n_5951;
wire n_1728;
wire n_4315;
wire n_5647;
wire n_3239;
wire n_2631;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_4857;
wire n_1651;
wire n_3087;
wire n_4637;
wire n_5523;
wire n_2697;
wire n_1263;
wire n_1817;
wire n_3704;
wire n_4296;
wire n_2677;
wire n_2483;
wire n_5088;
wire n_5773;
wire n_1032;
wire n_1592;
wire n_5392;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_3589;
wire n_1743;
wire n_720;
wire n_1943;
wire n_5138;
wire n_4588;
wire n_5149;
wire n_1163;
wire n_3054;
wire n_4970;
wire n_5280;
wire n_4153;
wire n_1868;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_2373;
wire n_3881;
wire n_5089;
wire n_5775;
wire n_2099;
wire n_3759;
wire n_3323;
wire n_4643;
wire n_2617;
wire n_808;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_1439;
wire n_3466;
wire n_2074;
wire n_5031;
wire n_1665;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_5082;
wire n_4788;
wire n_1414;
wire n_2067;
wire n_4555;
wire n_5230;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_2117;
wire n_1053;
wire n_5796;
wire n_5296;
wire n_5398;
wire n_1906;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_1828;
wire n_1304;
wire n_3335;
wire n_5960;
wire n_3007;
wire n_2267;
wire n_5858;
wire n_1349;
wire n_1061;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_3370;
wire n_874;
wire n_3949;
wire n_2286;
wire n_5192;
wire n_4247;
wire n_5051;
wire n_5336;
wire n_3036;
wire n_2783;
wire n_4583;
wire n_1015;
wire n_1162;
wire n_4292;
wire n_2118;
wire n_1490;
wire n_5552;
wire n_3764;
wire n_1553;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_1086;
wire n_3025;
wire n_3051;
wire n_986;
wire n_2802;
wire n_1104;
wire n_887;
wire n_2125;
wire n_1156;
wire n_4974;
wire n_5123;
wire n_2861;
wire n_4344;
wire n_5242;
wire n_3130;
wire n_1188;
wire n_1498;
wire n_4856;
wire n_2618;
wire n_4216;
wire n_957;
wire n_1242;
wire n_2707;
wire n_5596;
wire n_2849;
wire n_1489;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_5742;
wire n_5127;
wire n_4313;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_1119;
wire n_3713;
wire n_1863;
wire n_5933;
wire n_5536;
wire n_4798;
wire n_1500;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_1189;
wire n_5810;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_1523;
wire n_2190;
wire n_3931;
wire n_2516;
wire n_4991;
wire n_3070;
wire n_1005;
wire n_5818;
wire n_3275;
wire n_5198;
wire n_3245;
wire n_2894;
wire n_2452;
wire n_4182;
wire n_2827;
wire n_3214;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5539;
wire n_5009;
wire n_3710;
wire n_1844;
wire n_1957;
wire n_1953;
wire n_1219;
wire n_5889;
wire n_3944;
wire n_5632;
wire n_4729;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_5613;
wire n_4800;
wire n_1373;
wire n_1540;
wire n_5427;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_5450;
wire n_832;
wire n_744;
wire n_2821;
wire n_3696;
wire n_1331;
wire n_4781;
wire n_1529;
wire n_3531;
wire n_5124;
wire n_4237;
wire n_5297;
wire n_4828;
wire n_3333;
wire n_4652;
wire n_4114;
wire n_1007;
wire n_1580;
wire n_3135;
wire n_4925;
wire n_5719;
wire n_2448;
wire n_2211;
wire n_951;
wire n_5904;
wire n_5318;
wire n_5374;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_722;
wire n_3277;
wire n_4863;
wire n_1766;
wire n_5463;
wire n_1338;
wire n_2978;
wire n_4859;
wire n_4568;
wire n_3617;
wire n_2958;
wire n_1714;
wire n_1044;
wire n_4429;
wire n_5435;
wire n_3340;
wire n_5053;
wire n_5476;
wire n_5483;
wire n_1243;
wire n_5511;
wire n_3486;
wire n_2457;
wire n_2992;
wire n_3197;
wire n_3256;
wire n_1878;
wire n_3646;
wire n_5829;
wire n_2520;
wire n_811;
wire n_791;
wire n_5881;
wire n_3864;
wire n_4694;
wire n_1025;
wire n_4664;
wire n_3450;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_1406;
wire n_5073;
wire n_4306;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_4288;
wire n_3452;
wire n_4098;
wire n_2691;
wire n_5894;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_2991;
wire n_5419;
wire n_1596;
wire n_4289;
wire n_4972;
wire n_2723;
wire n_1476;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_5165;
wire n_2850;
wire n_1874;
wire n_5077;
wire n_3780;
wire n_1657;
wire n_3753;
wire n_1488;
wire n_4846;
wire n_1330;
wire n_906;
wire n_2295;
wire n_5225;
wire n_4076;
wire n_3142;
wire n_3129;
wire n_3495;
wire n_3843;
wire n_4805;
wire n_2606;
wire n_2386;
wire n_5826;
wire n_4822;
wire n_5931;
wire n_1829;
wire n_4635;
wire n_1450;
wire n_5532;
wire n_3740;
wire n_5441;
wire n_2417;
wire n_1815;
wire n_1493;
wire n_2911;
wire n_3313;
wire n_2354;
wire n_4281;
wire n_3945;
wire n_3726;
wire n_4419;
wire n_5405;
wire n_1256;
wire n_5365;
wire n_3560;
wire n_3345;
wire n_5772;
wire n_3421;
wire n_1448;
wire n_1009;
wire n_3548;
wire n_4906;
wire n_4630;
wire n_4829;
wire n_2612;
wire n_5259;
wire n_3236;
wire n_1995;
wire n_1397;
wire n_5921;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_4966;
wire n_2250;
wire n_1117;
wire n_3321;
wire n_1303;
wire n_4188;
wire n_2001;
wire n_2506;
wire n_2413;
wire n_4825;
wire n_2610;
wire n_3715;
wire n_1593;
wire n_2626;
wire n_2892;
wire n_2605;
wire n_2804;
wire n_5884;
wire n_5006;
wire n_4882;
wire n_3206;
wire n_5728;
wire n_1035;
wire n_3475;
wire n_4878;
wire n_2070;
wire n_3842;
wire n_1367;
wire n_4202;
wire n_2044;
wire n_5679;
wire n_3886;
wire n_825;
wire n_732;
wire n_2619;
wire n_1192;
wire n_5141;
wire n_3098;
wire n_4503;
wire n_1291;
wire n_5208;
wire n_5113;
wire n_3987;
wire n_5205;
wire n_4249;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_3386;
wire n_3921;
wire n_2177;
wire n_2766;
wire n_4196;
wire n_1197;
wire n_2613;
wire n_5667;
wire n_1517;
wire n_2647;
wire n_5508;
wire n_5105;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_5879;
wire n_1671;
wire n_5027;
wire n_2343;
wire n_1048;
wire n_775;
wire n_3380;
wire n_5688;
wire n_2826;
wire n_5825;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_5629;
wire n_5759;
wire n_2411;
wire n_4631;
wire n_1504;
wire n_2110;
wire n_5377;
wire n_3822;
wire n_889;
wire n_4355;
wire n_3818;
wire n_5599;
wire n_3587;
wire n_2608;
wire n_1948;
wire n_4155;
wire n_810;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_3497;
wire n_4542;
wire n_5451;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_5460;
wire n_4685;
wire n_3927;
wire n_2068;
wire n_3595;
wire n_1194;
wire n_4060;
wire n_1647;
wire n_1454;
wire n_2459;
wire n_941;
wire n_3396;
wire n_5517;
wire n_5807;
wire n_5426;
wire n_4093;
wire n_5693;
wire n_5695;
wire n_4123;
wire n_4294;
wire n_1521;
wire n_1940;
wire n_3683;
wire n_4452;
wire n_3887;
wire n_3195;
wire n_5587;
wire n_4722;
wire n_3048;
wire n_3339;
wire n_4164;
wire n_4126;
wire n_5030;
wire n_2963;
wire n_5674;
wire n_2561;
wire n_1056;
wire n_5584;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_1749;
wire n_1653;
wire n_4088;
wire n_2669;
wire n_3911;
wire n_3802;
wire n_4366;
wire n_1584;
wire n_848;
wire n_5125;
wire n_4922;
wire n_4733;
wire n_1814;
wire n_2441;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_4935;
wire n_4509;
wire n_2073;
wire n_4004;
wire n_5238;
wire n_750;
wire n_834;
wire n_3630;
wire n_1612;
wire n_800;
wire n_1910;
wire n_5906;
wire n_2189;
wire n_5732;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_2602;
wire n_5780;
wire n_724;
wire n_2931;
wire n_3433;
wire n_5556;
wire n_3597;
wire n_5743;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_5633;
wire n_3786;
wire n_875;
wire n_2828;
wire n_1626;
wire n_5950;
wire n_1335;
wire n_1715;
wire n_4204;
wire n_3553;
wire n_5323;
wire n_3645;
wire n_793;
wire n_5705;
wire n_4996;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_3550;
wire n_5510;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_1805;
wire n_4068;
wire n_5440;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_3610;
wire n_2443;
wire n_5011;
wire n_1554;
wire n_3279;
wire n_5513;
wire n_5875;
wire n_972;
wire n_4262;
wire n_2923;
wire n_2843;
wire n_3714;
wire n_4832;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_5848;
wire n_1679;
wire n_5834;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_5784;
wire n_3125;
wire n_5128;
wire n_2356;
wire n_5618;
wire n_4672;
wire n_2564;
wire n_3558;
wire n_3034;
wire n_3502;
wire n_783;
wire n_4053;
wire n_1127;
wire n_1008;
wire n_3963;
wire n_3091;
wire n_1024;
wire n_5157;
wire n_4496;
wire n_2518;
wire n_936;
wire n_4596;
wire n_5178;
wire n_3105;
wire n_1525;
wire n_4628;
wire n_1775;
wire n_908;
wire n_1036;
wire n_4083;
wire n_1270;
wire n_1272;
wire n_2794;
wire n_2901;
wire n_3940;
wire n_3225;
wire n_3621;
wire n_5529;
wire n_3473;
wire n_3680;
wire n_3565;
wire n_5388;
wire n_5824;
wire n_5354;
wire n_2453;
wire n_3331;
wire n_1788;
wire n_2138;
wire n_3040;
wire n_4230;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_2000;
wire n_5276;
wire n_4037;
wire n_3804;
wire n_4659;
wire n_3211;
wire n_917;
wire n_5196;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2215;
wire n_3847;
wire n_4073;
wire n_1261;
wire n_5763;
wire n_3633;
wire n_857;
wire n_1235;
wire n_2584;
wire n_4001;
wire n_1462;
wire n_5701;
wire n_1064;
wire n_1446;
wire n_1701;
wire n_3111;
wire n_731;
wire n_1813;
wire n_2997;
wire n_1573;
wire n_3258;
wire n_758;
wire n_3691;
wire n_2252;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_5907;
wire n_784;
wire n_4339;
wire n_4690;
wire n_2987;
wire n_1473;
wire n_1076;
wire n_1348;
wire n_5895;
wire n_2651;
wire n_753;
wire n_2733;
wire n_2445;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_2522;
wire n_3632;
wire n_1344;
wire n_4064;
wire n_3351;
wire n_5478;
wire n_1141;
wire n_3457;
wire n_5384;
wire n_840;
wire n_2324;
wire n_5283;
wire n_3454;
wire n_5961;
wire n_2139;
wire n_2521;
wire n_5686;
wire n_2740;
wire n_1991;
wire n_4066;
wire n_4681;
wire n_3303;
wire n_4414;
wire n_2541;
wire n_5094;
wire n_3232;
wire n_1113;
wire n_3768;
wire n_4295;
wire n_1615;
wire n_4100;
wire n_1265;
wire n_2372;
wire n_2105;
wire n_3445;
wire n_1806;
wire n_4087;
wire n_1409;
wire n_1684;
wire n_1148;
wire n_1588;
wire n_1673;
wire n_4473;
wire n_4619;
wire n_5371;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_3018;
wire n_1875;
wire n_2429;
wire n_5286;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_1039;
wire n_5676;
wire n_5949;
wire n_5040;
wire n_1150;
wire n_4266;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_1136;
wire n_1190;
wire n_5885;
wire n_3628;
wire n_4777;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_5399;
wire n_2846;
wire n_3371;
wire n_4918;
wire n_5856;
wire n_3872;
wire n_5760;
wire n_4415;
wire n_5110;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_1777;
wire n_3366;
wire n_5844;
wire n_3441;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_2545;
wire n_2513;
wire n_4408;
wire n_2115;
wire n_2017;
wire n_1810;
wire n_1347;
wire n_4976;
wire n_860;
wire n_3555;
wire n_5938;
wire n_3534;
wire n_4548;
wire n_2670;
wire n_3556;
wire n_896;
wire n_4574;
wire n_2644;
wire n_4557;
wire n_3071;
wire n_1698;
wire n_1337;
wire n_774;
wire n_2148;
wire n_5548;
wire n_1168;
wire n_4663;
wire n_5840;
wire n_3296;
wire n_3762;
wire n_3794;
wire n_4624;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_4686;
wire n_2384;
wire n_1705;
wire n_768;
wire n_3707;
wire n_3895;
wire n_1091;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_5917;
wire n_2058;
wire n_3231;
wire n_1846;
wire n_4161;
wire n_5304;
wire n_5437;
wire n_1581;
wire n_946;
wire n_757;
wire n_2047;
wire n_3058;
wire n_1655;
wire n_3709;
wire n_3398;
wire n_1146;
wire n_5355;
wire n_998;
wire n_3592;
wire n_5321;
wire n_2536;
wire n_1604;
wire n_3399;
wire n_4772;
wire n_5915;
wire n_1368;
wire n_963;
wire n_4120;
wire n_925;
wire n_2880;
wire n_1313;
wire n_1001;
wire n_3722;
wire n_4716;
wire n_4654;
wire n_1115;
wire n_1339;
wire n_1051;
wire n_5116;
wire n_3771;
wire n_719;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_1010;
wire n_2830;
wire n_5500;
wire n_4622;
wire n_4757;
wire n_803;
wire n_1871;
wire n_5669;
wire n_5672;
wire n_4016;
wire n_3334;
wire n_5621;
wire n_2940;
wire n_3427;
wire n_3162;
wire n_5569;
wire n_4591;
wire n_5966;
wire n_5515;
wire n_3083;
wire n_4570;
wire n_2491;
wire n_1931;
wire n_5559;
wire n_2259;
wire n_5337;
wire n_849;
wire n_5059;
wire n_4655;
wire n_1820;
wire n_1233;
wire n_4493;
wire n_1808;
wire n_1635;
wire n_1704;
wire n_4896;
wire n_4851;
wire n_2479;
wire n_886;
wire n_1308;
wire n_1451;
wire n_1487;
wire n_5528;
wire n_5605;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_2484;
wire n_5753;
wire n_5358;
wire n_1469;
wire n_4901;
wire n_3480;
wire n_1355;
wire n_4213;
wire n_4127;
wire n_2500;
wire n_2334;
wire n_5467;
wire n_1169;
wire n_789;
wire n_3181;
wire n_5493;
wire n_1916;
wire n_4602;
wire n_1713;
wire n_1436;
wire n_2818;
wire n_4900;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_3745;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_1515;
wire n_817;
wire n_5901;
wire n_1566;
wire n_2837;
wire n_717;
wire n_952;
wire n_2446;
wire n_4116;
wire n_5360;
wire n_2671;
wire n_2702;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_1138;
wire n_4103;
wire n_2529;
wire n_2374;
wire n_5439;
wire n_1225;
wire n_3154;
wire n_1366;
wire n_3938;
wire n_2278;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_5250;
wire n_4416;
wire n_4439;
wire n_870;
wire n_4985;
wire n_3382;
wire n_3930;
wire n_3808;
wire n_5471;
wire n_2248;
wire n_813;
wire n_4660;
wire n_3081;
wire n_5497;
wire n_5519;
wire n_995;
wire n_2579;
wire n_1961;
wire n_1535;
wire n_2960;
wire n_3270;
wire n_871;
wire n_2844;
wire n_1979;
wire n_829;
wire n_4814;
wire n_2221;
wire n_5502;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_3657;
wire n_5706;
wire n_2634;
wire n_2746;
wire n_5098;
wire n_721;
wire n_1084;
wire n_1276;
wire n_5145;
wire n_2878;
wire n_3830;
wire n_3252;
wire n_5466;
wire n_1528;
wire n_3315;
wire n_3523;
wire n_3999;
wire n_3420;
wire n_3859;
wire n_868;
wire n_5213;
wire n_3474;
wire n_5738;
wire n_2458;
wire n_5592;
wire n_5620;
wire n_3150;
wire n_5491;
wire n_1542;
wire n_4831;
wire n_4782;
wire n_1539;
wire n_2859;
wire n_5216;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_5953;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_5703;
wire n_1636;
wire n_4597;
wire n_4546;
wire n_5187;
wire n_4031;
wire n_5119;
wire n_1254;
wire n_4147;
wire n_1703;
wire n_3073;
wire n_3571;
wire n_4576;
wire n_3297;
wire n_5148;
wire n_3003;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_5330;
wire n_1560;
wire n_2899;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5526;
wire n_5202;
wire n_3817;
wire n_2722;
wire n_3728;
wire n_5107;
wire n_4680;
wire n_5067;
wire n_1012;
wire n_2061;
wire n_2685;
wire n_2512;
wire n_1790;
wire n_2788;
wire n_1443;
wire n_5264;
wire n_2595;
wire n_1465;
wire n_3084;
wire n_4593;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_3554;
wire n_2717;
wire n_1391;
wire n_2981;
wire n_1006;
wire n_4995;
wire n_1159;
wire n_5873;
wire n_4498;
wire n_772;
wire n_1245;
wire n_5741;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_3758;
wire n_5423;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_3777;
wire n_1872;
wire n_1585;
wire n_3767;
wire n_5926;
wire n_5866;
wire n_3692;
wire n_1351;
wire n_3234;
wire n_2216;
wire n_2426;
wire n_4850;
wire n_1260;
wire n_3716;
wire n_2926;
wire n_4937;
wire n_798;
wire n_5574;
wire n_3391;
wire n_5877;
wire n_912;
wire n_4786;
wire n_5203;
wire n_4354;
wire n_4235;
wire n_3159;
wire n_2855;
wire n_794;
wire n_2848;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_1292;
wire n_1026;
wire n_3460;
wire n_1610;
wire n_5155;
wire n_2202;
wire n_2952;
wire n_3530;
wire n_2693;
wire n_5408;
wire n_5812;
wire n_5540;
wire n_5804;
wire n_3240;
wire n_5066;
wire n_931;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_967;
wire n_5130;
wire n_4175;
wire n_1079;
wire n_5200;
wire n_3393;
wire n_2836;
wire n_2864;
wire n_4456;
wire n_1717;
wire n_2172;
wire n_2601;
wire n_2365;
wire n_1880;
wire n_5684;
wire n_1399;
wire n_1855;
wire n_2333;
wire n_3629;
wire n_4948;
wire n_5413;
wire n_1903;
wire n_2147;
wire n_4020;
wire n_5150;
wire n_5111;
wire n_1226;
wire n_2224;
wire n_1970;
wire n_3724;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_3046;
wire n_2921;
wire n_1240;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_5444;
wire n_3257;
wire n_5737;
wire n_3730;
wire n_5615;
wire n_3979;
wire n_5097;
wire n_2695;
wire n_2598;
wire n_3727;
wire n_976;
wire n_4003;
wire n_1832;
wire n_767;
wire n_2302;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_5640;
wire n_3342;
wire n_2895;
wire n_3796;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_5550;
wire n_3375;
wire n_2768;
wire n_3760;
wire n_5661;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_5306;
wire n_5905;
wire n_2728;
wire n_2025;
wire n_3744;
wire n_5457;
wire n_5159;
wire n_4022;
wire n_1020;
wire n_2495;
wire n_1058;
wire n_4336;
wire n_5314;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_1279;
wire n_2511;
wire n_3981;
wire n_2681;
wire n_1689;
wire n_2535;
wire n_1255;
wire n_3031;
wire n_2335;
wire n_5482;
wire n_3215;
wire n_1401;
wire n_3138;
wire n_776;
wire n_2860;
wire n_2041;
wire n_1933;
wire n_4494;
wire n_4201;
wire n_5287;
wire n_4719;
wire n_5651;
wire n_3577;
wire n_4074;
wire n_3994;
wire n_4636;
wire n_4983;
wire n_3185;
wire n_1217;
wire n_2662;
wire n_4386;
wire n_3917;
wire n_1231;
wire n_5623;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_5524;
wire n_926;
wire n_2296;
wire n_5735;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_4225;
wire n_4658;
wire n_4186;
wire n_1501;
wire n_2241;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_2531;
wire n_1570;
wire n_3377;
wire n_1518;
wire n_4907;
wire n_3961;
wire n_5153;
wire n_855;
wire n_2059;
wire n_4713;
wire n_5787;
wire n_1287;
wire n_1611;
wire n_3374;
wire n_4870;
wire n_4818;
wire n_5935;
wire n_4916;
wire n_5967;
wire n_4323;
wire n_5934;
wire n_1899;
wire n_5376;
wire n_3508;
wire n_4129;
wire n_5488;
wire n_1105;
wire n_5727;
wire n_3599;
wire n_5646;
wire n_4480;
wire n_5711;
wire n_3734;
wire n_5832;
wire n_3401;
wire n_983;
wire n_3542;
wire n_3263;
wire n_5891;
wire n_2523;
wire n_1945;
wire n_2418;
wire n_1614;
wire n_1377;
wire n_5328;
wire n_3819;
wire n_3222;
wire n_1740;
wire n_4616;
wire n_5016;
wire n_5470;
wire n_1092;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_1963;
wire n_3868;
wire n_729;
wire n_2218;
wire n_1122;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_5362;
wire n_2754;
wire n_4580;
wire n_1218;
wire n_3611;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_877;
wire n_3995;
wire n_3908;
wire n_1055;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_1089;
wire n_1502;
wire n_3501;
wire n_1478;
wire n_2555;
wire n_3216;
wire n_3568;
wire n_2708;
wire n_735;
wire n_4844;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_845;
wire n_1649;
wire n_2470;
wire n_1297;
wire n_3551;
wire n_1708;
wire n_5037;
wire n_5650;
wire n_5729;
wire n_5581;
wire n_4677;
wire n_5189;
wire n_4525;
wire n_3364;
wire n_2643;
wire n_755;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_4369;
wire n_3826;
wire n_5648;
wire n_2266;
wire n_4324;
wire n_842;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_742;
wire n_5160;
wire n_1719;
wire n_2742;
wire n_769;
wire n_3671;
wire n_2366;
wire n_5762;
wire n_1753;
wire n_5484;
wire n_1372;
wire n_1895;
wire n_4104;
wire n_982;
wire n_3791;
wire n_915;
wire n_2008;
wire n_4989;
wire n_5874;
wire n_3064;
wire n_3199;
wire n_2127;
wire n_3151;
wire n_3016;
wire n_2460;
wire n_1319;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_4528;
wire n_2772;
wire n_1700;
wire n_1332;
wire n_5385;
wire n_1747;
wire n_3990;
wire n_5622;
wire n_1171;
wire n_5635;
wire n_4069;
wire n_3582;
wire n_4280;
wire n_1867;
wire n_5609;
wire n_3993;
wire n_2576;
wire n_3459;
wire n_4811;
wire n_2696;
wire n_5595;
wire n_5256;
wire n_4779;
wire n_5910;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_5380;
wire n_1400;
wire n_3735;
wire n_1527;
wire n_1513;
wire n_3656;
wire n_4524;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_5568;
wire n_5941;
wire n_4891;
wire n_2629;
wire n_3369;
wire n_1257;
wire n_1954;
wire n_3964;
wire n_5364;
wire n_3302;
wire n_5597;
wire n_2486;
wire n_1897;
wire n_5469;
wire n_2137;
wire n_3685;
wire n_4977;
wire n_2492;
wire n_2939;
wire n_3425;
wire n_4876;
wire n_5021;
wire n_1449;
wire n_2900;
wire n_797;
wire n_2912;
wire n_5936;
wire n_1405;
wire n_3813;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_1757;
wire n_1950;
wire n_2264;
wire n_805;
wire n_5928;
wire n_2032;
wire n_2090;
wire n_3124;
wire n_3811;
wire n_4200;
wire n_2249;
wire n_5785;
wire n_3411;
wire n_5222;
wire n_3463;
wire n_2785;
wire n_730;
wire n_4938;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_1856;
wire n_1524;
wire n_2928;
wire n_5505;
wire n_1118;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_1293;
wire n_961;
wire n_726;
wire n_5504;
wire n_878;
wire n_4118;
wire n_3857;
wire n_3110;
wire n_4239;
wire n_3157;
wire n_1180;
wire n_1697;
wire n_2730;
wire n_5129;
wire n_806;
wire n_1350;
wire n_4704;
wire n_2720;
wire n_1561;
wire n_5494;
wire n_5970;
wire n_2405;
wire n_2700;
wire n_1616;
wire n_2416;
wire n_2064;
wire n_3640;
wire n_5663;
wire n_5161;
wire n_1557;
wire n_4744;
wire n_5378;
wire n_5626;
wire n_4706;
wire n_3879;
wire n_2022;
wire n_4343;
wire n_1505;
wire n_2408;
wire n_4764;
wire n_5389;
wire n_4990;
wire n_2986;
wire n_949;
wire n_2454;
wire n_3591;
wire n_2760;
wire n_4919;
wire n_1208;
wire n_3317;
wire n_5653;
wire n_4835;
wire n_1151;
wire n_4420;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_5266;
wire n_4559;
wire n_4742;
wire n_5038;
wire n_3566;
wire n_5800;
wire n_1133;
wire n_883;
wire n_4372;
wire n_5396;
wire n_4097;
wire n_4162;
wire n_5766;
wire n_5293;
wire n_779;
wire n_4790;
wire n_4173;
wire n_5309;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_1269;
wire n_4727;
wire n_1547;
wire n_1438;
wire n_3654;
wire n_5627;
wire n_1047;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_1288;
wire n_2173;
wire n_3982;
wire n_3647;
wire n_1143;
wire n_3973;
wire n_4799;
wire n_5882;
wire n_4534;
wire n_5636;
wire n_4960;
wire n_1153;
wire n_1103;
wire n_5707;
wire n_5594;
wire n_3738;
wire n_894;
wire n_5697;
wire n_1380;
wire n_2020;
wire n_5606;
wire n_2310;
wire n_5911;
wire n_3600;
wire n_1023;
wire n_914;
wire n_5382;
wire n_4327;
wire n_3190;
wire n_3027;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_3733;
wire n_1165;
wire n_3967;
wire n_4370;
wire n_5638;
wire n_4816;
wire n_4091;
wire n_5058;
wire n_1417;
wire n_3096;
wire n_4166;
wire n_2777;
wire n_5356;
wire n_2234;
wire n_1341;
wire n_5849;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_1603;
wire n_5841;
wire n_4478;
wire n_2935;
wire n_4246;
wire n_715;
wire n_1066;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_4061;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_4754;
wire n_1534;
wire n_1290;
wire n_4375;
wire n_2396;
wire n_3368;
wire n_1559;
wire n_3117;
wire n_4684;
wire n_743;
wire n_1546;
wire n_3384;
wire n_5279;
wire n_2592;
wire n_3490;
wire n_962;
wire n_5043;
wire n_4241;
wire n_2751;
wire n_3113;
wire n_1622;
wire n_4183;
wire n_918;
wire n_1968;
wire n_5645;
wire n_5020;
wire n_2842;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_5232;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_1193;
wire n_1345;
wire n_5035;
wire n_3037;
wire n_1336;
wire n_1033;
wire n_5453;
wire n_4333;
wire n_5339;
wire n_5443;
wire n_1166;
wire n_2007;
wire n_3363;
wire n_1158;
wire n_1803;
wire n_872;
wire n_3522;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_5631;
wire n_3481;
wire n_5101;
wire n_2236;
wire n_4457;
wire n_2150;
wire n_1816;
wire n_2803;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_3305;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_3354;
wire n_5608;
wire n_2204;
wire n_1481;
wire n_2040;
wire n_2151;
wire n_2455;
wire n_827;
wire n_3437;
wire n_2231;
wire n_4212;
wire n_4584;
wire n_5702;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_4477;
wire n_5806;
wire n_4110;
wire n_5182;
wire n_1221;
wire n_4217;
wire n_5277;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_1579;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_923;
wire n_1124;
wire n_1326;
wire n_3969;
wire n_2282;
wire n_4605;
wire n_981;
wire n_3873;
wire n_4649;
wire n_5747;
wire n_1204;
wire n_2428;
wire n_994;
wire n_1360;
wire n_2858;
wire n_3076;
wire n_3410;
wire n_5415;
wire n_856;
wire n_4592;
wire n_4999;
wire n_1564;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_1361;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_5687;
wire n_1411;
wire n_1359;
wire n_3536;
wire n_1721;
wire n_3782;
wire n_1317;
wire n_3594;
wire n_5383;
wire n_2385;
wire n_5690;
wire n_1980;
wire n_5740;
wire n_4177;
wire n_2501;
wire n_1385;
wire n_1998;
wire n_5029;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_2985;
wire n_5218;
wire n_2630;
wire n_2028;
wire n_919;
wire n_3114;
wire n_2092;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_2402;
wire n_1458;
wire n_3047;
wire n_3163;
wire n_5361;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_5512;
wire n_2808;
wire n_2344;
wire n_3520;
wire n_2392;
wire n_3272;
wire n_3122;
wire n_5898;
wire n_5923;
wire n_3687;
wire n_2787;
wire n_5617;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_5946;
wire n_1268;
wire n_2676;
wire n_2770;
wire n_4550;
wire n_4347;
wire n_5193;
wire n_4933;
wire n_968;
wire n_4144;
wire n_5514;
wire n_5611;
wire n_2375;
wire n_3278;
wire n_5579;
wire n_4167;
wire n_3608;
wire n_4895;
wire n_1282;
wire n_4726;
wire n_5573;
wire n_5143;
wire n_5836;
wire n_1755;
wire n_5188;
wire n_5049;
wire n_2212;
wire n_5308;
wire n_4434;
wire n_5068;
wire n_5739;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_816;
wire n_1322;
wire n_3829;
wire n_4510;
wire n_5057;
wire n_5425;
wire n_5273;
wire n_5839;
wire n_2469;
wire n_1125;
wire n_2358;
wire n_1710;
wire n_3546;
wire n_2355;
wire n_1390;
wire n_5887;
wire n_3068;
wire n_1629;
wire n_1094;
wire n_5683;
wire n_1510;
wire n_3002;
wire n_1099;
wire n_5248;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_759;
wire n_4156;
wire n_1727;
wire n_3693;
wire n_5880;
wire n_3132;
wire n_5002;
wire n_5487;
wire n_5649;
wire n_5531;
wire n_831;
wire n_3681;
wire n_5666;
wire n_3970;
wire n_778;
wire n_2351;
wire n_1619;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_1152;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_1236;
wire n_4579;
wire n_4776;
wire n_2704;
wire n_1334;
wire n_3729;
wire n_4471;
wire n_4392;
wire n_3103;
wire n_2048;
wire n_3028;
wire n_4691;
wire n_3148;
wire n_3775;
wire n_5682;
wire n_5461;
wire n_3966;
wire n_4397;
wire n_3616;
wire n_4753;
wire n_4803;
wire n_1289;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_5730;
wire n_4165;
wire n_2056;
wire n_5754;
wire n_2852;
wire n_2515;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1941;
wire n_3637;
wire n_1017;
wire n_734;
wire n_4893;
wire n_2240;
wire n_4258;
wire n_5756;
wire n_2917;
wire n_3194;
wire n_2085;
wire n_2432;
wire n_5033;
wire n_1686;
wire n_4232;
wire n_5075;
wire n_2097;
wire n_3461;
wire n_1410;
wire n_939;
wire n_2297;
wire n_4203;
wire n_5789;
wire n_5400;
wire n_1325;
wire n_1223;
wire n_5347;
wire n_2957;
wire n_1983;
wire n_4767;
wire n_4569;
wire n_948;
wire n_3820;
wire n_5144;
wire n_3072;
wire n_2961;
wire n_4468;
wire n_5509;
wire n_1923;
wire n_3848;
wire n_3631;
wire n_5169;
wire n_4885;
wire n_1479;
wire n_4698;
wire n_1031;
wire n_3674;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_5349;
wire n_3763;
wire n_933;
wire n_3499;
wire n_5534;
wire n_1821;
wire n_3910;
wire n_3947;
wire n_2585;
wire n_5183;
wire n_3361;
wire n_2995;
wire n_4533;
wire n_4287;
wire n_3228;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_1186;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_4556;
wire n_2205;
wire n_2183;
wire n_3088;
wire n_1724;
wire n_1707;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_1126;
wire n_5079;
wire n_2761;
wire n_2357;
wire n_4520;
wire n_895;
wire n_1639;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_5751;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_5039;
wire n_1818;
wire n_4265;
wire n_3557;
wire n_1598;
wire n_2269;
wire n_1583;
wire n_4612;
wire n_5375;
wire n_5438;
wire n_1264;
wire n_4149;
wire n_1827;
wire n_4958;
wire n_1752;
wire n_2361;
wire n_4538;
wire n_3030;
wire n_3505;
wire n_5563;
wire n_3075;
wire n_1102;
wire n_2239;
wire n_1296;
wire n_4730;
wire n_4421;
wire n_2464;
wire n_3697;
wire n_882;
wire n_2304;
wire n_2514;
wire n_5932;
wire n_1299;
wire n_3430;
wire n_5919;
wire n_2063;
wire n_3489;
wire n_5012;
wire n_2079;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_3484;
wire n_4971;
wire n_2095;
wire n_5664;
wire n_2738;
wire n_5890;
wire n_2590;
wire n_4661;
wire n_2797;
wire n_3041;
wire n_5823;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_5422;
wire n_5944;
wire n_5246;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_1069;
wire n_4305;
wire n_2037;
wire n_2953;
wire n_2823;
wire n_3684;
wire n_5725;
wire n_5404;
wire n_913;
wire n_1681;
wire n_4834;
wire n_1507;
wire n_5332;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_2346;
wire n_4692;
wire n_1353;
wire n_3268;
wire n_2559;
wire n_5616;
wire n_1383;
wire n_4259;
wire n_5870;
wire n_2030;
wire n_850;
wire n_4299;
wire n_5625;
wire n_2407;
wire n_5367;
wire n_2243;
wire n_5288;
wire n_2694;
wire n_5601;
wire n_3742;
wire n_4965;
wire n_1837;
wire n_4178;
wire n_2006;
wire n_4953;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_5294;
wire n_5570;
wire n_2731;
wire n_3703;
wire n_5411;
wire n_5670;
wire n_1246;
wire n_5265;
wire n_5955;
wire n_2123;
wire n_2238;
wire n_4793;
wire n_4802;
wire n_1196;
wire n_5733;
wire n_3435;
wire n_2380;
wire n_1187;
wire n_4897;
wire n_1298;
wire n_1745;
wire n_4674;
wire n_4796;
wire n_1088;
wire n_766;
wire n_5184;
wire n_2750;
wire n_2547;
wire n_945;
wire n_4575;
wire n_3665;
wire n_3063;
wire n_3281;
wire n_3535;
wire n_5061;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_4589;
wire n_3220;
wire n_4581;
wire n_4625;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_4148;
wire n_3679;
wire n_738;
wire n_5575;
wire n_4968;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_4038;
wire n_3856;
wire n_5316;
wire n_2735;
wire n_953;
wire n_4214;
wire n_1888;
wire n_5290;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_3419;
wire n_989;
wire n_5048;
wire n_2233;
wire n_5363;
wire n_5665;
wire n_795;
wire n_4892;
wire n_1936;
wire n_3890;
wire n_821;
wire n_770;
wire n_5607;
wire n_1514;
wire n_2782;
wire n_3929;
wire n_971;
wire n_4353;
wire n_2201;
wire n_4950;
wire n_1650;
wire n_4176;
wire n_4124;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_5462;
wire n_4488;
wire n_5278;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_5214;
wire n_3756;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_5845;
wire n_4608;
wire n_3948;
wire n_4839;
wire n_1074;
wire n_5969;
wire n_1765;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_2332;
wire n_2391;
wire n_1295;
wire n_2060;
wire n_3883;
wire n_1013;
wire n_4032;
wire n_2571;
wire n_5736;
wire n_4929;
wire n_2874;
wire n_4117;
wire n_3049;
wire n_3634;
wire n_5436;
wire n_2341;
wire n_1654;
wire n_3066;
wire n_2045;
wire n_3913;
wire n_5341;
wire n_2575;
wire n_3739;
wire n_1230;
wire n_5140;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_4541;
wire n_3271;
wire n_3164;
wire n_3861;
wire n_5096;
wire n_2043;
wire n_4171;
wire n_5847;
wire n_4815;
wire n_4665;
wire n_5639;
wire n_4884;
wire n_3580;
wire n_1437;
wire n_4276;
wire n_1378;
wire n_5268;
wire n_5050;
wire n_5240;
wire n_5503;
wire n_1461;
wire n_5718;
wire n_1876;
wire n_1830;
wire n_5001;
wire n_5658;
wire n_1112;
wire n_4174;
wire n_5131;
wire n_5546;
wire n_5174;
wire n_2145;
wire n_4801;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_3119;
wire n_4740;
wire n_1108;
wire n_1274;
wire n_4394;
wire n_5544;
wire n_5660;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_5541;
wire n_5610;
wire n_916;
wire n_2810;
wire n_1884;
wire n_1555;
wire n_762;
wire n_1253;
wire n_1468;
wire n_4378;
wire n_5166;
wire n_2683;
wire n_4180;
wire n_4459;
wire n_3624;
wire n_5808;
wire n_1182;
wire n_4594;
wire n_2748;
wire n_4642;
wire n_1376;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1506;
wire n_3544;
wire n_5300;
wire n_2072;
wire n_3852;
wire n_5233;
wire n_5381;
wire n_5770;
wire n_5710;
wire n_2628;
wire n_1491;
wire n_3219;
wire n_1083;
wire n_5333;
wire n_5799;
wire n_4914;
wire n_3510;
wire n_4587;
wire n_1139;
wire n_3688;
wire n_5008;
wire n_1312;
wire n_3871;
wire n_892;
wire n_3757;
wire n_1567;
wire n_2219;
wire n_2100;
wire n_3666;
wire n_5538;
wire n_990;
wire n_867;
wire n_3479;
wire n_944;
wire n_5499;
wire n_749;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_4285;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_3741;
wire n_5582;
wire n_2567;
wire n_2557;
wire n_1908;
wire n_5675;
wire n_1155;
wire n_2755;
wire n_1071;
wire n_5109;
wire n_909;
wire n_1392;
wire n_2066;
wire n_5281;
wire n_2762;
wire n_964;
wire n_2220;
wire n_4433;
wire n_2829;
wire n_5862;
wire n_1914;
wire n_2253;
wire n_5886;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_1633;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_5285;
wire n_2328;
wire n_2434;
wire n_1234;
wire n_3936;
wire n_5564;
wire n_2261;
wire n_3082;
wire n_5162;
wire n_5442;
wire n_2473;
wire n_5802;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_3867;
wire n_3397;
wire n_1646;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_1237;
wire n_5883;
wire n_1095;
wire n_3078;
wire n_3971;
wire n_5630;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_1531;
wire n_2113;
wire n_1387;
wire n_3711;
wire n_5054;
wire n_3171;
wire n_5929;
wire n_5394;
wire n_4751;
wire n_4242;
wire n_5975;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_1496;
wire n_2812;
wire n_3300;
wire n_5496;
wire n_3104;
wire n_4122;
wire n_2132;
wire n_4522;
wire n_4952;
wire n_4426;
wire n_5956;
wire n_5699;
wire n_4362;
wire n_3267;
wire n_3946;
wire n_5920;
wire n_2112;
wire n_2640;
wire n_5000;
wire n_4634;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2983;
wire n_5211;
wire n_4089;
wire n_3513;
wire n_1173;
wire n_3498;
wire n_5132;
wire n_2350;
wire n_5535;
wire n_1068;
wire n_1198;
wire n_4506;
wire n_4728;
wire n_1886;
wire n_4346;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_3863;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_1365;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_3332;
wire n_2055;
wire n_2998;
wire n_1423;
wire n_4359;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_5176;
wire n_4039;
wire n_5793;
wire n_1798;
wire n_3057;
wire n_1608;
wire n_5761;
wire n_3983;
wire n_3318;
wire n_3385;
wire n_3773;
wire n_3494;
wire n_1278;
wire n_5074;
wire n_3788;
wire n_3939;
wire n_727;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_3260;
wire n_2496;
wire n_3349;
wire n_4348;
wire n_1602;
wire n_3139;
wire n_3801;
wire n_5681;
wire n_2338;
wire n_5261;
wire n_1080;
wire n_3636;
wire n_3653;
wire n_3823;
wire n_3403;
wire n_2057;
wire n_1205;
wire n_2716;
wire n_2944;
wire n_2780;
wire n_3439;
wire n_1120;
wire n_1202;
wire n_4084;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_2774;
wire n_2799;
wire n_5748;
wire n_4393;
wire n_3984;
wire n_1586;
wire n_1431;
wire n_4389;
wire n_1763;
wire n_5641;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_4615;
wire n_3044;
wire n_3492;
wire n_3737;
wire n_5657;
wire n_3579;
wire n_2379;
wire n_1667;
wire n_888;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_1677;
wire n_5244;
wire n_5765;
wire n_5114;
wire n_4551;
wire n_4521;
wire n_2284;
wire n_3005;
wire n_5420;
wire n_2283;
wire n_5206;
wire n_2526;
wire n_1097;
wire n_1711;
wire n_4387;
wire n_3186;
wire n_2508;
wire n_2594;
wire n_1239;
wire n_5298;
wire n_3417;
wire n_890;
wire n_3626;
wire n_4598;
wire n_4464;
wire n_5106;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_1081;
wire n_2119;
wire n_2493;
wire n_5080;
wire n_4565;
wire n_3392;
wire n_1800;
wire n_5081;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_3512;
wire n_1734;
wire n_1860;
wire n_4552;
wire n_2840;
wire n_4482;
wire n_837;
wire n_812;
wire n_4172;
wire n_5957;
wire n_4040;
wire n_3024;
wire n_5567;
wire n_5406;
wire n_4328;
wire n_1854;
wire n_5191;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_2893;
wire n_4940;
wire n_785;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_5867;
wire n_1394;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_873;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_4112;
wire n_5602;
wire n_2035;
wire n_4928;
wire n_2614;
wire n_5428;
wire n_2494;
wire n_1538;
wire n_4865;
wire n_2128;
wire n_4071;
wire n_4436;
wire n_5786;
wire n_5822;
wire n_3586;
wire n_5817;
wire n_4160;
wire n_1668;
wire n_5798;
wire n_4137;
wire n_1078;
wire n_5417;
wire n_4545;
wire n_4758;
wire n_1161;
wire n_4840;
wire n_5713;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_1191;
wire n_4535;
wire n_4385;
wire n_1215;
wire n_3748;
wire n_4731;
wire n_2337;
wire n_1786;
wire n_3732;
wire n_1804;
wire n_4671;
wire n_2272;
wire n_5571;
wire n_4766;
wire n_4558;
wire n_1318;
wire n_1769;
wire n_1632;
wire n_1929;
wire n_4319;
wire n_2929;
wire n_4358;
wire n_1526;
wire n_4874;
wire n_2656;
wire n_4904;
wire n_1997;
wire n_1137;
wire n_1258;
wire n_1733;
wire n_4651;
wire n_943;
wire n_3167;
wire n_4748;
wire n_1807;
wire n_1123;
wire n_2857;
wire n_1784;
wire n_4618;
wire n_3787;
wire n_4025;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_752;
wire n_985;
wire n_5506;
wire n_5475;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_5908;
wire n_1352;
wire n_5431;
wire n_5100;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_5315;
wire n_2633;
wire n_3708;
wire n_5752;
wire n_2907;
wire n_1429;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_5746;
wire n_1154;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_1130;
wire n_3718;
wire n_756;
wire n_3390;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_4666;
wire n_4082;
wire n_3140;
wire n_2320;
wire n_979;
wire n_3976;
wire n_3381;
wire n_2546;
wire n_2813;
wire n_897;
wire n_3736;
wire n_4466;
wire n_891;
wire n_885;
wire n_3955;
wire n_1659;
wire n_5366;
wire n_5322;
wire n_1864;
wire n_5414;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_3336;
wire n_5903;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_5151;
wire n_714;
wire n_3605;
wire n_5307;
wire n_2170;
wire n_4721;
wire n_725;
wire n_1577;
wire n_5003;
wire n_3840;
wire n_2198;
wire n_5369;
wire n_3067;
wire n_3809;
wire n_4921;
wire n_1852;
wire n_801;
wire n_5912;
wire n_5745;
wire n_4377;
wire n_818;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_5803;
wire n_5593;
wire n_5270;
wire n_5853;
wire n_3468;
wire n_5779;
wire n_1877;
wire n_4301;
wire n_5313;
wire n_2133;
wire n_2497;
wire n_879;
wire n_5446;
wire n_4561;
wire n_1541;
wire n_3291;
wire n_1472;
wire n_1050;
wire n_2578;
wire n_1201;
wire n_1185;
wire n_2475;
wire n_4715;
wire n_2715;
wire n_2665;
wire n_4879;
wire n_5044;
wire n_1090;
wire n_3755;
wire n_4536;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_5459;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_4418;
wire n_3341;
wire n_4125;
wire n_5390;
wire n_5351;
wire n_5267;
wire n_1116;
wire n_5024;
wire n_3043;
wire n_2747;
wire n_1511;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_4151;
wire n_2845;
wire n_4412;
wire n_2036;
wire n_843;
wire n_3358;
wire n_2533;
wire n_2003;
wire n_1307;
wire n_4682;
wire n_1128;
wire n_2419;
wire n_2330;
wire n_5078;
wire n_4810;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_1955;
wire n_3289;
wire n_1440;
wire n_1370;
wire n_5005;
wire n_1549;
wire n_5207;
wire n_2658;
wire n_5624;
wire n_3620;
wire n_4601;
wire n_1065;
wire n_4518;
wire n_2767;
wire n_5474;
wire n_3376;
wire n_1362;
wire n_3123;
wire n_5447;
wire n_2692;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_5700;
wire n_5755;
wire n_2862;
wire n_4325;
wire n_1420;
wire n_2645;
wire n_2553;
wire n_4711;
wire n_2749;
wire n_5962;
wire n_4413;
wire n_1210;
wire n_3307;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2833;
wire n_1038;
wire n_3723;
wire n_4135;
wire n_5223;
wire n_5662;
wire n_3880;
wire n_5801;
wire n_3904;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_3405;
wire n_2313;
wire n_1022;
wire n_5465;
wire n_3532;
wire n_5154;
wire n_5721;
wire n_2609;
wire n_1767;
wire n_1040;
wire n_3131;
wire n_4138;
wire n_1973;
wire n_1444;
wire n_820;
wire n_2882;
wire n_2303;
wire n_4384;
wire n_4639;
wire n_1664;
wire n_4577;
wire n_2154;
wire n_1986;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_984;
wire n_5087;
wire n_1552;
wire n_2938;
wire n_2498;
wire n_3992;
wire n_1772;
wire n_1311;
wire n_3106;
wire n_2881;
wire n_3092;
wire n_4270;
wire n_4620;
wire n_5397;
wire n_4924;
wire n_4044;
wire n_2305;
wire n_880;
wire n_5566;
wire n_3304;
wire n_4388;
wire n_3247;
wire n_739;
wire n_1028;
wire n_4271;
wire n_2180;
wire n_4406;
wire n_2809;
wire n_5652;
wire n_975;
wire n_1645;
wire n_5805;
wire n_932;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_3785;
wire n_5492;
wire n_2465;
wire n_5501;
wire n_2972;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_3178;
wire n_2251;
wire n_5758;
wire n_5842;
wire n_3100;
wire n_3721;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_5692;
wire n_4973;
wire n_4792;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_2487;
wire n_5473;
wire n_1834;
wire n_1011;
wire n_2534;
wire n_2941;
wire n_4286;
wire n_3638;
wire n_3576;
wire n_5562;
wire n_4858;
wire n_1445;
wire n_5370;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_5458;
wire n_2387;
wire n_4318;
wire n_5227;
wire n_830;
wire n_5902;
wire n_987;
wire n_2510;
wire n_3570;
wire n_3227;
wire n_5359;
wire n_4673;
wire n_2793;
wire n_5282;
wire n_2639;
wire n_4738;
wire n_2603;
wire n_5386;
wire n_1167;
wire n_4554;
wire n_4526;
wire n_4105;
wire n_3663;
wire n_969;
wire n_1663;
wire n_5952;
wire n_2086;
wire n_1926;
wire n_1630;
wire n_1720;
wire n_2966;
wire n_2409;
wire n_3431;
wire n_3355;
wire n_1738;
wire n_5716;
wire n_3897;
wire n_1735;
wire n_5888;
wire n_4005;
wire n_4181;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_956;
wire n_765;
wire n_4092;
wire n_4875;
wire n_4255;
wire n_2758;
wire n_5036;
wire n_1271;
wire n_2186;
wire n_5790;
wire n_4647;
wire n_3575;
wire n_2471;
wire n_3042;
wire n_1067;
wire n_1323;
wire n_1937;
wire n_4142;
wire n_5118;
wire n_900;
wire n_5485;
wire n_5525;
wire n_3004;
wire n_1551;
wire n_4849;
wire n_5271;
wire n_2039;
wire n_1285;
wire n_733;
wire n_761;
wire n_3838;
wire n_4059;
wire n_5194;
wire n_5445;
wire n_2734;
wire n_5948;
wire n_4499;
wire n_4504;
wire n_3598;
wire n_4917;
wire n_2420;
wire n_3273;
wire n_2918;
wire n_835;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_1792;
wire n_5628;
wire n_5245;
wire n_2062;
wire n_4489;
wire n_822;
wire n_1459;
wire n_2153;
wire n_5329;
wire n_5472;
wire n_839;
wire n_1754;
wire n_4833;
wire n_3394;
wire n_2235;
wire n_5850;
wire n_1575;
wire n_4564;
wire n_1848;
wire n_1172;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_3581;
wire n_5072;
wire n_3778;
wire n_4322;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_2206;
wire n_997;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_5940;
wire n_3001;
wire n_5260;
wire n_4981;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_5372;
wire n_4507;
wire n_4756;
wire n_1576;
wire n_5860;
wire n_2422;
wire n_2933;
wire n_3387;
wire n_3952;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_1059;
wire n_2736;
wire n_3825;
wire n_4198;
wire n_977;
wire n_2339;
wire n_2532;
wire n_4373;
wire n_1866;
wire n_2664;
wire n_4154;
wire n_5859;
wire n_4390;
wire n_1782;
wire n_1558;
wire n_4107;
wire n_2519;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_2360;
wire n_4453;
wire n_723;
wire n_1393;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_809;
wire n_3032;
wire n_5612;
wire n_4886;
wire n_5172;
wire n_881;
wire n_1477;
wire n_1019;
wire n_1982;
wire n_5311;
wire n_910;
wire n_5164;
wire n_4964;
wire n_4700;
wire n_4002;
wire n_1114;
wire n_1742;
wire n_4679;
wire n_3815;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_1273;
wire n_2982;
wire n_5495;
wire n_4483;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_5547;
wire n_4693;
wire n_1043;
wire n_5121;
wire n_4956;
wire n_2869;
wire n_5379;
wire n_4487;
wire n_5878;
wire n_2674;
wire n_5820;
wire n_1737;
wire n_1613;
wire n_3026;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_3244;
wire n_1779;
wire n_2562;
wire n_954;
wire n_3112;
wire n_2051;
wire n_3196;
wire n_5964;
wire n_2673;
wire n_4678;
wire n_1591;
wire n_5301;
wire n_5126;
wire n_2548;
wire n_3488;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_5776;
wire n_2179;
wire n_1280;
wire n_3779;
wire n_1063;
wire n_991;
wire n_2275;
wire n_4606;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_5603;
wire n_938;
wire n_1891;
wire n_5348;
wire n_1000;
wire n_4868;
wire n_4072;
wire n_2792;
wire n_4465;
wire n_2596;
wire n_5217;
wire n_3986;
wire n_5558;
wire n_3725;
wire n_4026;
wire n_4245;
wire n_5520;
wire n_2524;
wire n_3894;
wire n_1702;
wire n_5909;
wire n_4852;
wire n_3202;
wire n_4290;
wire n_4945;
wire n_5750;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1082;
wire n_1725;
wire n_5654;
wire n_2318;
wire n_866;
wire n_2819;
wire n_1722;
wire n_2229;
wire n_1644;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_2255;
wire n_5554;
wire n_1252;
wire n_3045;
wire n_773;
wire n_5135;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_5448;
wire n_2573;
wire n_5837;
wire n_2336;
wire n_5412;
wire n_1662;
wire n_3249;
wire n_3483;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_782;
wire n_2915;
wire n_4869;
wire n_3213;
wire n_5533;
wire n_4047;
wire n_1244;
wire n_1796;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_1574;
wire n_3033;
wire n_893;
wire n_1582;
wire n_1981;
wire n_2824;
wire n_5327;
wire n_4417;
wire n_796;
wire n_1374;
wire n_2089;
wire n_4688;
wire n_4939;
wire n_5900;
wire n_1486;
wire n_3619;
wire n_4013;
wire n_3434;
wire n_4342;
wire n_4903;
wire n_2131;
wire n_3853;
wire n_4382;
wire n_2509;
wire n_4085;
wire n_5486;
wire n_2135;
wire n_4475;
wire n_5432;
wire n_5851;
wire n_1463;
wire n_4626;
wire n_4997;
wire n_5065;
wire n_924;
wire n_781;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_2436;
wire n_3517;
wire n_1706;
wire n_2461;
wire n_3719;
wire n_1214;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_5295;
wire n_1181;
wire n_1999;
wire n_4841;
wire n_4683;
wire n_5173;
wire n_2873;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_5655;
wire n_3383;
wire n_1835;
wire n_5855;
wire n_3965;
wire n_1457;
wire n_3905;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_4600;
wire n_5861;
wire n_1453;
wire n_3943;
wire n_3145;
wire n_5749;
wire n_2908;
wire n_4106;
wire n_2156;
wire n_1184;
wire n_754;
wire n_2323;
wire n_1073;
wire n_4549;
wire n_1277;
wire n_1746;
wire n_1062;
wire n_4702;
wire n_5102;
wire n_4954;
wire n_740;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_3283;
wire n_4331;
wire n_4159;
wire n_3451;
wire n_4734;
wire n_2832;
wire n_1688;
wire n_5827;
wire n_2370;
wire n_1944;
wire n_2914;
wire n_5656;
wire n_1988;
wire n_5678;
wire n_5865;
wire n_1718;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_2539;
wire n_5555;
wire n_2078;
wire n_1145;
wire n_4809;
wire n_787;
wire n_4012;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_5212;
wire n_4760;
wire n_1207;
wire n_3606;
wire n_2232;
wire n_1847;
wire n_5815;
wire n_4320;
wire n_5084;
wire n_5251;
wire n_1314;
wire n_1512;
wire n_5965;
wire n_884;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_5407;
wire n_2988;
wire n_4560;
wire n_3230;
wire n_3793;
wire n_859;
wire n_5042;
wire n_4768;
wire n_1889;
wire n_5368;
wire n_929;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_3607;
wire n_1637;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_5310;
wire n_2769;
wire n_1548;
wire n_4987;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_2739;
wire n_3962;
wire n_4988;
wire n_2902;
wire n_4360;
wire n_1544;
wire n_4540;
wire n_2094;
wire n_5588;
wire n_3854;
wire n_1354;
wire n_2349;
wire n_3652;
wire n_3449;
wire n_1021;
wire n_3089;
wire n_4854;
wire n_1595;
wire n_1142;
wire n_5477;
wire n_2727;
wire n_942;
wire n_5234;
wire n_1416;
wire n_1599;
wire n_5871;
wire n_4747;
wire n_3472;
wire n_2527;
wire n_3126;
wire n_2759;
wire n_5007;
wire n_4881;
wire n_2038;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_1838;
wire n_4357;
wire n_2806;
wire n_4502;
wire n_3191;
wire n_1716;
wire n_5334;
wire n_3562;
wire n_2281;
wire n_5253;
wire n_3588;
wire n_1590;
wire n_3280;
wire n_4115;
wire n_5274;
wire n_5418;
wire n_5019;
wire n_5939;
wire n_1819;
wire n_3095;
wire n_947;
wire n_5792;
wire n_3698;
wire n_4513;
wire n_1179;
wire n_1442;
wire n_4775;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_2499;
wire n_2549;
wire n_804;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_3885;
wire n_955;
wire n_4264;
wire n_5954;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_3839;
wire n_5490;
wire n_5694;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_5489;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_3120;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_4794;
wire n_4843;
wire n_5580;
wire n_5215;
wire n_3937;
wire n_4763;
wire n_1418;
wire n_5795;
wire n_5715;
wire n_4170;
wire n_5561;
wire n_2462;
wire n_2155;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_3604;
wire n_5430;
wire n_824;
wire n_5659;
wire n_4272;
wire n_5195;
wire n_3176;
wire n_3792;
wire n_5720;
wire n_4267;
wire n_2083;
wire n_815;
wire n_5598;
wire n_2753;
wire n_1340;
wire n_3021;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_2898;
wire n_1825;
wire n_3567;
wire n_2682;
wire n_5854;
wire n_5958;
wire n_5585;
wire n_5112;
wire n_5326;
wire n_1627;
wire n_5783;
wire n_2903;
wire n_5303;
wire n_3812;
wire n_3127;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_5530;
wire n_965;
wire n_5809;
wire n_934;
wire n_2213;
wire n_4056;
wire n_4806;
wire n_1674;
wire n_4015;
wire n_2924;
wire n_4445;
wire n_4462;
wire n_5299;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_1042;
wire n_3170;
wire n_2311;
wire n_1455;
wire n_2287;
wire n_836;
wire n_3415;
wire n_3464;
wire n_3414;
wire n_4234;
wire n_760;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_3467;
wire n_5821;
wire n_3179;
wire n_5522;
wire n_4836;
wire n_3889;
wire n_5262;
wire n_3262;
wire n_5319;
wire n_927;
wire n_3699;
wire n_2120;
wire n_1419;
wire n_3816;
wire n_3528;
wire n_4207;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_4725;
wire n_2312;
wire n_1826;
wire n_5943;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_5335;
wire n_1259;
wire n_2801;
wire n_4334;
wire n_1177;
wire n_5284;
wire n_4978;
wire n_5771;
wire n_3246;
wire n_3299;
wire n_980;
wire n_1618;
wire n_1869;
wire n_3623;
wire n_905;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_5516;
wire n_3615;
wire n_1802;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_3200;
wire n_3642;
wire n_2146;
wire n_4274;
wire n_5583;
wire n_3276;
wire n_5433;
wire n_3682;
wire n_5429;
wire n_5698;
wire n_5731;
wire n_4007;
wire n_1456;
wire n_1879;
wire n_2129;
wire n_5857;
wire n_814;
wire n_5120;
wire n_3572;
wire n_2975;
wire n_2399;
wire n_1134;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_2027;
wire n_2932;
wire n_3118;
wire n_5560;
wire n_4441;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_5455;
wire n_1467;
wire n_5209;
wire n_5704;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_5916;
wire n_3705;
wire n_3022;
wire n_1709;
wire n_5099;
wire n_3286;
wire n_5781;
wire n_5619;
wire n_2023;
wire n_3974;
wire n_3443;
wire n_2599;
wire n_3988;
wire n_5022;
wire n_2075;
wire n_1726;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_5353;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_1098;
wire n_3009;
wire n_777;
wire n_5219;
wire n_920;
wire n_3951;
wire n_5518;
wire n_3035;
wire n_4261;
wire n_1132;
wire n_1823;
wire n_5236;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_2254;
wire n_3290;
wire n_1402;
wire n_3957;
wire n_3418;
wire n_1607;
wire n_5673;
wire n_861;
wire n_5814;
wire n_1666;
wire n_5103;
wire n_4648;
wire n_2214;
wire n_2256;
wire n_3326;
wire n_2732;
wire n_1883;
wire n_4094;
wire n_2776;
wire n_3224;
wire n_1969;
wire n_5671;
wire n_2949;
wire n_4269;
wire n_1927;
wire n_1222;
wire n_3803;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_4913;
wire n_2449;
wire n_4428;
wire n_745;
wire n_1572;
wire n_4463;
wire n_5357;
wire n_3648;
wire n_1975;
wire n_5421;
wire n_1388;
wire n_1266;
wire n_4396;
wire n_1990;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_1075;
wire n_1890;
wire n_4034;
wire n_4228;
wire n_1227;
wire n_3166;
wire n_3649;
wire n_3065;
wire n_5045;
wire n_5237;
wire n_3924;
wire n_3997;
wire n_3564;
wire n_862;
wire n_5769;
wire n_2637;
wire n_3795;
wire n_4931;
wire n_2306;
wire n_2071;
wire n_3953;
wire n_4400;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_5434;
wire n_1532;
wire n_1030;
wire n_5181;
wire n_3208;
wire n_5768;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_852;
wire n_2916;
wire n_1060;
wire n_5963;
wire n_4424;
wire n_4351;
wire n_4192;
wire n_1748;
wire n_1301;
wire n_5972;
wire n_3400;
wire n_1466;
wire n_2581;
wire n_5937;
wire n_1783;
wire n_5146;
wire n_4646;
wire n_4221;
wire n_3650;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_4035;
wire n_1480;
wire n_3670;
wire n_2540;
wire n_4190;
wire n_1605;
wire n_3060;
wire n_2984;
wire n_4009;
wire n_2489;
wire n_5013;
wire n_4145;
wire n_5577;
wire n_876;
wire n_5872;
wire n_5017;
wire n_736;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_2106;
wire n_4717;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_854;
wire n_2091;
wire n_4312;
wire n_5424;
wire n_3789;
wire n_1658;
wire n_1072;
wire n_1305;
wire n_4750;
wire n_2348;
wire n_1873;
wire n_2667;
wire n_2725;
wire n_3746;
wire n_4537;
wire n_1046;
wire n_5838;
wire n_3694;
wire n_771;
wire n_5456;
wire n_3893;
wire n_4847;
wire n_5846;
wire n_2307;
wire n_3702;
wire n_5930;
wire n_1984;
wire n_3453;
wire n_1556;
wire n_5345;
wire n_2815;
wire n_4427;
wire n_1824;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_819;
wire n_1971;
wire n_2945;
wire n_1324;
wire n_3543;
wire n_1776;
wire n_3448;
wire n_4279;
wire n_2936;
wire n_3609;
wire n_4330;
wire n_4152;
wire n_5537;
wire n_2698;
wire n_5572;
wire n_4783;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_5409;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_807;
wire n_5142;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_1987;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_802;
wire n_5401;
wire n_4595;
wire n_960;
wire n_2352;
wire n_5201;
wire n_5816;
wire n_790;
wire n_5551;
wire n_5416;
wire n_4404;
wire n_2377;
wire n_2652;
wire n_5498;
wire n_5543;
wire n_4054;
wire n_1286;
wire n_4617;
wire n_1685;
wire n_2477;
wire n_4611;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_5797;
wire n_1052;
wire n_4732;
wire n_2076;
wire n_2203;
wire n_5942;
wire n_5764;
wire n_1426;
wire n_4969;
wire n_5252;
wire n_5777;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_4140;
wire n_5171;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_3309;
wire n_2796;
wire n_858;
wire n_5393;
wire n_4817;
wire n_2136;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_2771;
wire n_2403;
wire n_2947;
wire n_5643;
wire n_928;
wire n_3769;
wire n_1565;
wire n_4437;
wire n_3055;
wire n_4070;
wire n_5346;
wire n_748;
wire n_1045;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_4139;
wire n_4769;
wire n_5868;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_2713;
wire n_1422;
wire n_1965;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_2934;
wire n_5104;
wire n_2210;
wire n_4368;
wire n_5794;
wire n_3141;
wire n_2053;
wire n_5272;
wire n_3476;
wire n_1049;
wire n_4430;
wire n_3238;
wire n_2450;
wire n_5338;
wire n_1356;
wire n_1773;
wire n_3175;
wire n_4544;
wire n_2666;
wire n_5578;
wire n_728;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_3255;
wire n_2588;
wire n_5722;
wire n_5811;
wire n_935;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_911;
wire n_3509;
wire n_1403;
wire n_5395;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_3456;
wire n_4532;
wire n_5863;
wire n_3790;
wire n_907;
wire n_5734;
wire n_847;
wire n_747;
wire n_1135;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_3662;
wire n_5774;
wire n_5199;
wire n_4257;
wire n_4282;
wire n_4341;
wire n_1694;
wire n_1695;
wire n_4027;
wire n_4309;
wire n_4650;
wire n_5480;
wire n_3077;
wire n_4944;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_4994;
wire n_3533;
wire n_5175;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_3409;
wire n_4381;
wire n_3583;
wire n_4316;
wire n_4860;
wire n_4469;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_1157;
wire n_5959;
wire n_3563;
wire n_5945;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_3689;
wire n_1789;
wire n_763;
wire n_2174;
wire n_5668;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_4703;
wire n_1687;
wire n_4934;
wire n_2638;
wire n_2046;
wire n_1756;
wire n_4350;
wire n_1606;
wire n_5600;
wire n_1587;
wire n_2340;
wire n_4804;
wire n_2444;
wire n_4888;
wire n_1014;
wire n_5767;
wire n_1427;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_2199;
wire n_4669;
wire n_5228;
wire n_1100;
wire n_1617;
wire n_2600;
wire n_3436;
wire n_5973;
wire n_1962;
wire n_3806;
wire n_4759;
wire n_5869;
wire n_5914;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_1175;
wire n_4887;
wire n_3751;
wire n_3402;
wire n_1621;
wire n_5186;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_3664;
wire n_4218;
wire n_4687;
wire n_1381;
wire n_3686;
wire n_1183;
wire n_4720;
wire n_2889;
wire n_2141;
wire n_1758;
wire n_1110;
wire n_5604;
wire n_3470;
wire n_5221;
wire n_1407;
wire n_2865;
wire n_5925;
wire n_973;
wire n_5591;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_1176;
wire n_3677;
wire n_1054;
wire n_5387;
wire n_3292;
wire n_3989;
wire n_4644;
wire n_4752;
wire n_4746;
wire n_1057;
wire n_4131;
wire n_5449;
wire n_4215;
wire n_978;
wire n_2488;
wire n_1509;
wire n_828;
wire n_4158;
wire n_3079;
wire n_5190;
wire n_3269;
wire n_5325;
wire n_4231;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_4926;
wire n_2050;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_5876;
wire n_5344;
wire n_2550;
wire n_1536;
wire n_3177;
wire n_4667;
wire n_5813;
wire n_1471;
wire n_3440;
wire n_3658;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1620;
wire n_2542;
wire n_5892;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_788;
wire n_5714;
wire n_2169;
wire n_5634;
wire n_5133;
wire n_5305;
wire n_2175;
wire n_1625;
wire n_5689;
wire n_4578;
wire n_5644;
wire n_3644;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_1922;
wire n_940;
wire n_1537;
wire n_4877;
wire n_2065;
wire n_4470;
wire n_4187;
wire n_1904;
wire n_4998;
wire n_5576;
wire n_2395;
wire n_2868;
wire n_1530;
wire n_4057;
wire n_5852;
wire n_5918;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_898;
wire n_3328;
wire n_2012;
wire n_3182;
wire n_2967;
wire n_5343;
wire n_1093;
wire n_4021;
wire n_3379;
wire n_4379;
wire n_5947;
wire n_2268;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_5835;
wire n_2111;
wire n_3743;
wire n_5542;
wire n_2948;
wire n_5015;
wire n_3099;
wire n_5527;
wire n_2897;
wire n_4812;
wire n_4497;
wire n_2583;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1770;
wire n_1003;
wire n_4472;
wire n_2699;
wire n_5819;
wire n_3901;
wire n_5180;
wire n_1640;
wire n_2973;
wire n_5893;
wire n_2710;
wire n_2505;
wire n_4519;
wire n_5025;
wire n_2397;
wire n_3878;
wire n_4197;
wire n_2721;
wire n_1892;
wire n_2615;
wire n_4787;
wire n_1212;
wire n_4310;
wire n_4566;
wire n_3933;
wire n_5726;
wire n_4371;
wire n_1902;
wire n_5828;
wire n_2784;
wire n_3898;
wire n_4749;
wire n_5924;
wire n_1845;
wire n_921;
wire n_5545;
wire n_2104;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_5083;
wire n_3253;
wire n_2088;
wire n_1275;
wire n_4238;
wire n_904;
wire n_2005;
wire n_1696;
wire n_2108;
wire n_3824;
wire n_2246;
wire n_5899;
wire n_3846;
wire n_5122;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_3845;
wire n_3203;
wire n_4986;
wire n_1316;
wire n_4668;
wire n_950;
wire n_5782;
wire n_4168;
wire n_1369;
wire n_4298;
wire n_4743;
wire n_1781;
wire n_4250;
wire n_3143;
wire n_3690;
wire n_3229;
wire n_5864;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_5637;
wire n_4211;
wire n_3094;
wire n_741;
wire n_5185;
wire n_2964;
wire n_5032;
wire n_865;
wire n_5034;
wire n_3312;
wire n_1041;
wire n_2451;
wire n_2913;
wire n_993;
wire n_1862;
wire n_3752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_2839;
wire n_3237;
wire n_4128;
wire n_4036;
wire n_5269;
wire n_3655;
wire n_2955;
wire n_5709;
wire n_1764;
wire n_4807;
wire n_5115;
wire n_902;
wire n_1723;
wire n_3918;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_4095;
wire n_1310;
wire n_5927;
wire n_4485;
wire n_3593;
wire n_5163;
wire n_1229;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_1896;
wire n_1516;
wire n_4890;
wire n_2485;
wire n_2563;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_5507;
wire n_4573;
wire n_1328;
wire n_4943;
wire n_2875;
wire n_3519;
wire n_2209;
wire n_4042;
wire n_4244;
wire n_1928;
wire n_5642;
wire n_4708;
wire n_4883;
wire n_4553;
wire n_1634;
wire n_1203;
wire n_1699;
wire n_5226;
wire n_2081;
wire n_937;
wire n_1474;
wire n_1631;
wire n_1794;
wire n_5696;
wire n_1375;
wire n_3053;
wire n_5014;
wire n_3772;
wire n_2891;
wire n_4335;
wire n_3128;
wire n_5677;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_1002;
wire n_4516;
wire n_5235;
wire n_1129;
wire n_1464;
wire n_2798;
wire n_3217;
wire n_1249;
wire n_5724;
wire n_3821;
wire n_3201;
wire n_3503;
wire n_1870;
wire n_4467;
wire n_5521;
wire n_2654;
wire n_3935;
wire n_1861;
wire n_1228;
wire n_2319;
wire n_2965;
wire n_4955;
wire n_5410;
wire n_1251;
wire n_1989;
wire n_2689;
wire n_1762;
wire n_3798;
wire n_3080;
wire n_5241;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_4645;
wire n_5331;
wire n_3308;
wire n_841;
wire n_3204;
wire n_4134;
wire n_5018;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;
wire n_5258;

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_396),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_506),
.Y(n_715)
);

CKINVDCx20_ASAP7_75t_R g716 ( 
.A(n_219),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_709),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_710),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_686),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_525),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_107),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_304),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_519),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_201),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_390),
.Y(n_725)
);

INVxp33_ASAP7_75t_SL g726 ( 
.A(n_451),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_649),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_299),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_276),
.Y(n_729)
);

CKINVDCx20_ASAP7_75t_R g730 ( 
.A(n_394),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_358),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_479),
.Y(n_732)
);

CKINVDCx20_ASAP7_75t_R g733 ( 
.A(n_496),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_299),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_556),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_87),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_108),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_665),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_413),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_28),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_368),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_432),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_163),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_540),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_10),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_129),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_625),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_703),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_493),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_704),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_653),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_461),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_594),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_632),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_395),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_610),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_44),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_680),
.Y(n_758)
);

CKINVDCx14_ASAP7_75t_R g759 ( 
.A(n_326),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_17),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_165),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_527),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_380),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_84),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_297),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_350),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_20),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_561),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_78),
.Y(n_769)
);

CKINVDCx14_ASAP7_75t_R g770 ( 
.A(n_215),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_533),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_281),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_377),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_280),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_405),
.Y(n_775)
);

CKINVDCx20_ASAP7_75t_R g776 ( 
.A(n_631),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_360),
.Y(n_777)
);

CKINVDCx20_ASAP7_75t_R g778 ( 
.A(n_611),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_246),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_679),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_158),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_335),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_423),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_157),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_20),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_331),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_104),
.Y(n_787)
);

CKINVDCx20_ASAP7_75t_R g788 ( 
.A(n_471),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_58),
.Y(n_789)
);

CKINVDCx20_ASAP7_75t_R g790 ( 
.A(n_253),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_375),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_302),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_59),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_121),
.Y(n_794)
);

BUFx10_ASAP7_75t_L g795 ( 
.A(n_125),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_608),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_652),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_434),
.Y(n_798)
);

INVx1_ASAP7_75t_SL g799 ( 
.A(n_101),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_226),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_684),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_32),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_259),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_610),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_269),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_494),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_695),
.Y(n_807)
);

BUFx2_ASAP7_75t_L g808 ( 
.A(n_421),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_502),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_139),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_379),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_190),
.Y(n_812)
);

CKINVDCx20_ASAP7_75t_R g813 ( 
.A(n_176),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_303),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_286),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_444),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_477),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_244),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_494),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_206),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_358),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_698),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_422),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_672),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_681),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_420),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_4),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_527),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_19),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_96),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_196),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_638),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_548),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_294),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_650),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_281),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_300),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_526),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_262),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_466),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_327),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_261),
.Y(n_842)
);

INVxp33_ASAP7_75t_SL g843 ( 
.A(n_122),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_306),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_597),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_472),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_333),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_690),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_226),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_170),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_218),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_630),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_223),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_247),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_546),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_476),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_615),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_100),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_439),
.Y(n_859)
);

CKINVDCx20_ASAP7_75t_R g860 ( 
.A(n_162),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_107),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_346),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_464),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_645),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_601),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_691),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_431),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_643),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_332),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_355),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_2),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_250),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_428),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_414),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_1),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_535),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_411),
.Y(n_877)
);

CKINVDCx16_ASAP7_75t_R g878 ( 
.A(n_508),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_103),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_436),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_225),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_190),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_427),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_197),
.Y(n_884)
);

INVxp67_ASAP7_75t_L g885 ( 
.A(n_284),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_662),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_630),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_141),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_334),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_461),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_210),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_682),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_79),
.Y(n_893)
);

CKINVDCx14_ASAP7_75t_R g894 ( 
.A(n_298),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_378),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_295),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_364),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_585),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_238),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_6),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_188),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_198),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_713),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_409),
.Y(n_904)
);

INVx1_ASAP7_75t_SL g905 ( 
.A(n_557),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_409),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_641),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_174),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_43),
.Y(n_909)
);

BUFx2_ASAP7_75t_L g910 ( 
.A(n_116),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_706),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_272),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_132),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_705),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_64),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_559),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_60),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_586),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_108),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_694),
.Y(n_920)
);

BUFx5_ASAP7_75t_L g921 ( 
.A(n_353),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_711),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_656),
.Y(n_923)
);

CKINVDCx20_ASAP7_75t_R g924 ( 
.A(n_306),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_631),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_552),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_291),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_204),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_342),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_13),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_647),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_274),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_465),
.Y(n_933)
);

BUFx10_ASAP7_75t_L g934 ( 
.A(n_572),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_385),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_422),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_387),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_476),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_641),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_442),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_310),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_640),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_276),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_490),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_364),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_683),
.Y(n_946)
);

CKINVDCx16_ASAP7_75t_R g947 ( 
.A(n_94),
.Y(n_947)
);

CKINVDCx20_ASAP7_75t_R g948 ( 
.A(n_151),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_667),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_49),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_121),
.Y(n_951)
);

BUFx10_ASAP7_75t_L g952 ( 
.A(n_522),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_57),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_639),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_290),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_84),
.Y(n_956)
);

CKINVDCx20_ASAP7_75t_R g957 ( 
.A(n_676),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_465),
.Y(n_958)
);

BUFx2_ASAP7_75t_SL g959 ( 
.A(n_343),
.Y(n_959)
);

CKINVDCx16_ASAP7_75t_R g960 ( 
.A(n_248),
.Y(n_960)
);

BUFx10_ASAP7_75t_L g961 ( 
.A(n_671),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_499),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_384),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_242),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_528),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_269),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_371),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_625),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_477),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_708),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_469),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_129),
.Y(n_972)
);

BUFx10_ASAP7_75t_L g973 ( 
.A(n_480),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_104),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_373),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_545),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_349),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_66),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_534),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_144),
.Y(n_980)
);

BUFx5_ASAP7_75t_L g981 ( 
.A(n_372),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_531),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_376),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_530),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_127),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_290),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_503),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_492),
.Y(n_988)
);

BUFx8_ASAP7_75t_SL g989 ( 
.A(n_286),
.Y(n_989)
);

BUFx10_ASAP7_75t_L g990 ( 
.A(n_697),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_642),
.Y(n_991)
);

CKINVDCx20_ASAP7_75t_R g992 ( 
.A(n_674),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_270),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_471),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_655),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_193),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_474),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_701),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_558),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_537),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_21),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_340),
.Y(n_1002)
);

INVx1_ASAP7_75t_SL g1003 ( 
.A(n_39),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_547),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_668),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_144),
.Y(n_1006)
);

CKINVDCx16_ASAP7_75t_R g1007 ( 
.A(n_657),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_646),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_554),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_619),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_593),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_335),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_209),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_10),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_183),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_654),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_242),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_349),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_596),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_532),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_136),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_225),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_637),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_430),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_61),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_570),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_655),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_640),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_45),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_660),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_673),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_101),
.Y(n_1032)
);

CKINVDCx20_ASAP7_75t_R g1033 ( 
.A(n_113),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_582),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_252),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_675),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_259),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_266),
.Y(n_1038)
);

INVxp67_ASAP7_75t_L g1039 ( 
.A(n_439),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_106),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_340),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_528),
.Y(n_1042)
);

CKINVDCx20_ASAP7_75t_R g1043 ( 
.A(n_525),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_323),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_68),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_202),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_496),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_196),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_597),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_44),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_566),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_619),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_488),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_687),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_267),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_336),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_78),
.Y(n_1057)
);

CKINVDCx14_ASAP7_75t_R g1058 ( 
.A(n_623),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_418),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_712),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_359),
.Y(n_1061)
);

INVx1_ASAP7_75t_SL g1062 ( 
.A(n_1),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_643),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_157),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_518),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_586),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_642),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_413),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_266),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_651),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_15),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_592),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_427),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_685),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_96),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_573),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_490),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_24),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_18),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_173),
.Y(n_1080)
);

INVx2_ASAP7_75t_SL g1081 ( 
.A(n_699),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_244),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_689),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_663),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_587),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_43),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_111),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_233),
.Y(n_1088)
);

BUFx10_ASAP7_75t_L g1089 ( 
.A(n_173),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_298),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_250),
.Y(n_1091)
);

CKINVDCx20_ASAP7_75t_R g1092 ( 
.A(n_380),
.Y(n_1092)
);

CKINVDCx14_ASAP7_75t_R g1093 ( 
.A(n_360),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_141),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_31),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_150),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_654),
.Y(n_1097)
);

CKINVDCx20_ASAP7_75t_R g1098 ( 
.A(n_339),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_621),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_440),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_621),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_47),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_301),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_339),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_632),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_601),
.Y(n_1106)
);

BUFx10_ASAP7_75t_L g1107 ( 
.A(n_613),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_379),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_16),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_408),
.Y(n_1110)
);

INVx1_ASAP7_75t_SL g1111 ( 
.A(n_68),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_412),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_273),
.Y(n_1113)
);

BUFx5_ASAP7_75t_L g1114 ( 
.A(n_222),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_172),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_345),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_567),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_605),
.Y(n_1118)
);

CKINVDCx16_ASAP7_75t_R g1119 ( 
.A(n_105),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_62),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_48),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_201),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_135),
.Y(n_1123)
);

INVx1_ASAP7_75t_SL g1124 ( 
.A(n_311),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_664),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_436),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_283),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_219),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_170),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_516),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_628),
.Y(n_1131)
);

BUFx8_ASAP7_75t_SL g1132 ( 
.A(n_90),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_472),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_251),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_551),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_304),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_384),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_237),
.Y(n_1138)
);

CKINVDCx16_ASAP7_75t_R g1139 ( 
.A(n_479),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_49),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_543),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_158),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_65),
.Y(n_1143)
);

CKINVDCx16_ASAP7_75t_R g1144 ( 
.A(n_204),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_430),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_508),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_117),
.Y(n_1147)
);

CKINVDCx16_ASAP7_75t_R g1148 ( 
.A(n_416),
.Y(n_1148)
);

INVx1_ASAP7_75t_SL g1149 ( 
.A(n_628),
.Y(n_1149)
);

CKINVDCx20_ASAP7_75t_R g1150 ( 
.A(n_239),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_396),
.Y(n_1151)
);

INVx2_ASAP7_75t_SL g1152 ( 
.A(n_24),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_557),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_285),
.Y(n_1154)
);

INVx1_ASAP7_75t_SL g1155 ( 
.A(n_210),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_503),
.Y(n_1156)
);

CKINVDCx20_ASAP7_75t_R g1157 ( 
.A(n_639),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_321),
.Y(n_1158)
);

INVxp67_ASAP7_75t_L g1159 ( 
.A(n_277),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_352),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_29),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_584),
.Y(n_1162)
);

CKINVDCx16_ASAP7_75t_R g1163 ( 
.A(n_253),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_392),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_629),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_634),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_132),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_435),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_407),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_315),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_46),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_570),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_SL g1173 ( 
.A(n_536),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_359),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_651),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_5),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_404),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_644),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_317),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_287),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_328),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_275),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_554),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_258),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_692),
.Y(n_1185)
);

CKINVDCx16_ASAP7_75t_R g1186 ( 
.A(n_134),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_300),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_647),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_678),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_658),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_89),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_143),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_589),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_311),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_322),
.Y(n_1195)
);

CKINVDCx20_ASAP7_75t_R g1196 ( 
.A(n_63),
.Y(n_1196)
);

BUFx10_ASAP7_75t_L g1197 ( 
.A(n_636),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_707),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_702),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_453),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_95),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_256),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_262),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_700),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_216),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_445),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_462),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_9),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_562),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_373),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_594),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_34),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_195),
.Y(n_1213)
);

INVx1_ASAP7_75t_SL g1214 ( 
.A(n_576),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_624),
.Y(n_1215)
);

BUFx10_ASAP7_75t_L g1216 ( 
.A(n_192),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_581),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_155),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_541),
.Y(n_1219)
);

CKINVDCx16_ASAP7_75t_R g1220 ( 
.A(n_435),
.Y(n_1220)
);

CKINVDCx20_ASAP7_75t_R g1221 ( 
.A(n_54),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_183),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_341),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_519),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_151),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_656),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_547),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_480),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_389),
.Y(n_1229)
);

INVxp67_ASAP7_75t_L g1230 ( 
.A(n_410),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_693),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_0),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_446),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_629),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_98),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_696),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_115),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_61),
.Y(n_1238)
);

INVx2_ASAP7_75t_SL g1239 ( 
.A(n_272),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_677),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_294),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_561),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_401),
.Y(n_1243)
);

INVx1_ASAP7_75t_SL g1244 ( 
.A(n_81),
.Y(n_1244)
);

INVx2_ASAP7_75t_SL g1245 ( 
.A(n_659),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_648),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_562),
.Y(n_1247)
);

CKINVDCx20_ASAP7_75t_R g1248 ( 
.A(n_271),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_535),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_288),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_450),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_433),
.Y(n_1252)
);

CKINVDCx20_ASAP7_75t_R g1253 ( 
.A(n_688),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_65),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_188),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_575),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_462),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_315),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_137),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_463),
.Y(n_1260)
);

INVxp67_ASAP7_75t_SL g1261 ( 
.A(n_764),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_759),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_764),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_801),
.Y(n_1264)
);

CKINVDCx20_ASAP7_75t_R g1265 ( 
.A(n_1007),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_847),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_847),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_950),
.Y(n_1268)
);

INVxp33_ASAP7_75t_L g1269 ( 
.A(n_828),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_950),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1051),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1051),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1187),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_921),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1187),
.Y(n_1275)
);

INVxp67_ASAP7_75t_SL g1276 ( 
.A(n_1217),
.Y(n_1276)
);

INVxp33_ASAP7_75t_SL g1277 ( 
.A(n_1128),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1217),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_989),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1132),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_808),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_808),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_921),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_910),
.Y(n_1284)
);

INVx1_ASAP7_75t_SL g1285 ( 
.A(n_1173),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_910),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_986),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_986),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_921),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1021),
.Y(n_1290)
);

INVxp67_ASAP7_75t_L g1291 ( 
.A(n_1021),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_1064),
.Y(n_1292)
);

BUFx5_ASAP7_75t_L g1293 ( 
.A(n_718),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1064),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_1007),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_729),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_878),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_947),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_729),
.Y(n_1299)
);

INVxp67_ASAP7_75t_SL g1300 ( 
.A(n_732),
.Y(n_1300)
);

INVxp67_ASAP7_75t_L g1301 ( 
.A(n_959),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_737),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_737),
.Y(n_1303)
);

INVxp33_ASAP7_75t_SL g1304 ( 
.A(n_1231),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_960),
.Y(n_1305)
);

BUFx2_ASAP7_75t_L g1306 ( 
.A(n_770),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_743),
.Y(n_1307)
);

CKINVDCx20_ASAP7_75t_R g1308 ( 
.A(n_1139),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_801),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_743),
.Y(n_1310)
);

NOR2xp67_ASAP7_75t_L g1311 ( 
.A(n_744),
.B(n_0),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_746),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_921),
.Y(n_1313)
);

INVxp67_ASAP7_75t_L g1314 ( 
.A(n_959),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_746),
.Y(n_1315)
);

INVxp67_ASAP7_75t_L g1316 ( 
.A(n_1254),
.Y(n_1316)
);

INVxp67_ASAP7_75t_SL g1317 ( 
.A(n_732),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_747),
.Y(n_1318)
);

INVx1_ASAP7_75t_SL g1319 ( 
.A(n_716),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_747),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_1139),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_894),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_752),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_921),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_1058),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_752),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_921),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_762),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_762),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_921),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_765),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1144),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_765),
.Y(n_1333)
);

INVxp67_ASAP7_75t_L g1334 ( 
.A(n_766),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_766),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_773),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_773),
.Y(n_1337)
);

CKINVDCx16_ASAP7_75t_R g1338 ( 
.A(n_1093),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_801),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_783),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_783),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_785),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_785),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_791),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_791),
.Y(n_1345)
);

INVxp67_ASAP7_75t_SL g1346 ( 
.A(n_732),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_794),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_921),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_794),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_796),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_796),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_797),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_797),
.Y(n_1353)
);

INVxp33_ASAP7_75t_L g1354 ( 
.A(n_787),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_803),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_803),
.Y(n_1356)
);

BUFx5_ASAP7_75t_L g1357 ( 
.A(n_718),
.Y(n_1357)
);

CKINVDCx20_ASAP7_75t_R g1358 ( 
.A(n_1144),
.Y(n_1358)
);

OR2x2_ASAP7_75t_L g1359 ( 
.A(n_1186),
.B(n_2),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_810),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_810),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_820),
.Y(n_1362)
);

CKINVDCx20_ASAP7_75t_R g1363 ( 
.A(n_1186),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_820),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_921),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_848),
.B(n_3),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_981),
.Y(n_1367)
);

INVxp33_ASAP7_75t_SL g1368 ( 
.A(n_714),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_823),
.Y(n_1369)
);

INVxp67_ASAP7_75t_L g1370 ( 
.A(n_823),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_826),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_826),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_795),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_829),
.Y(n_1374)
);

XNOR2xp5_ASAP7_75t_L g1375 ( 
.A(n_720),
.B(n_3),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_829),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_830),
.Y(n_1377)
);

INVxp33_ASAP7_75t_SL g1378 ( 
.A(n_715),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_830),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_834),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_834),
.Y(n_1381)
);

CKINVDCx16_ASAP7_75t_R g1382 ( 
.A(n_1220),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_837),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_837),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_838),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1119),
.Y(n_1386)
);

INVxp67_ASAP7_75t_L g1387 ( 
.A(n_838),
.Y(n_1387)
);

INVxp33_ASAP7_75t_L g1388 ( 
.A(n_787),
.Y(n_1388)
);

INVx1_ASAP7_75t_SL g1389 ( 
.A(n_730),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_961),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_732),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_839),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_848),
.B(n_4),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_839),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_840),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_840),
.Y(n_1396)
);

CKINVDCx20_ASAP7_75t_R g1397 ( 
.A(n_1220),
.Y(n_1397)
);

CKINVDCx14_ASAP7_75t_R g1398 ( 
.A(n_961),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_841),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_841),
.Y(n_1400)
);

INVx2_ASAP7_75t_SL g1401 ( 
.A(n_795),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_842),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_733),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_842),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_853),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_853),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_801),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_855),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_767),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_855),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_857),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_857),
.Y(n_1412)
);

BUFx2_ASAP7_75t_SL g1413 ( 
.A(n_961),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_858),
.Y(n_1414)
);

INVxp33_ASAP7_75t_SL g1415 ( 
.A(n_721),
.Y(n_1415)
);

XOR2xp5_ASAP7_75t_L g1416 ( 
.A(n_774),
.B(n_5),
.Y(n_1416)
);

CKINVDCx16_ASAP7_75t_R g1417 ( 
.A(n_1148),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_858),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_859),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1163),
.Y(n_1420)
);

CKINVDCx20_ASAP7_75t_R g1421 ( 
.A(n_776),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_859),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_863),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_863),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_864),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_864),
.Y(n_1426)
);

INVx1_ASAP7_75t_SL g1427 ( 
.A(n_778),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_865),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_865),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_869),
.Y(n_1430)
);

INVxp67_ASAP7_75t_L g1431 ( 
.A(n_869),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_879),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_879),
.Y(n_1433)
);

INVxp33_ASAP7_75t_L g1434 ( 
.A(n_844),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_884),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_884),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1036),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_888),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_888),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_893),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_957),
.Y(n_1441)
);

INVxp67_ASAP7_75t_L g1442 ( 
.A(n_893),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_901),
.Y(n_1443)
);

INVxp33_ASAP7_75t_L g1444 ( 
.A(n_844),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_901),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_992),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_1253),
.Y(n_1447)
);

INVxp67_ASAP7_75t_L g1448 ( 
.A(n_904),
.Y(n_1448)
);

INVxp33_ASAP7_75t_SL g1449 ( 
.A(n_722),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_904),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_913),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_913),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_961),
.Y(n_1453)
);

CKINVDCx16_ASAP7_75t_R g1454 ( 
.A(n_795),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_915),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_915),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_930),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_930),
.Y(n_1458)
);

INVxp33_ASAP7_75t_L g1459 ( 
.A(n_849),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_931),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1036),
.Y(n_1461)
);

INVxp33_ASAP7_75t_L g1462 ( 
.A(n_849),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_931),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_937),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_937),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_990),
.Y(n_1466)
);

CKINVDCx16_ASAP7_75t_R g1467 ( 
.A(n_795),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_981),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_938),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_938),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_940),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_723),
.Y(n_1472)
);

XOR2xp5_ASAP7_75t_L g1473 ( 
.A(n_788),
.B(n_6),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_866),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_940),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_942),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_942),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_943),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_943),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_954),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_954),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_956),
.Y(n_1482)
);

CKINVDCx16_ASAP7_75t_R g1483 ( 
.A(n_934),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_956),
.Y(n_1484)
);

INVxp33_ASAP7_75t_SL g1485 ( 
.A(n_724),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_965),
.Y(n_1486)
);

INVxp67_ASAP7_75t_L g1487 ( 
.A(n_965),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_968),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_968),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_971),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_971),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_974),
.Y(n_1492)
);

INVxp67_ASAP7_75t_SL g1493 ( 
.A(n_732),
.Y(n_1493)
);

CKINVDCx14_ASAP7_75t_R g1494 ( 
.A(n_990),
.Y(n_1494)
);

INVxp33_ASAP7_75t_SL g1495 ( 
.A(n_725),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_974),
.Y(n_1496)
);

CKINVDCx16_ASAP7_75t_R g1497 ( 
.A(n_934),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_979),
.Y(n_1498)
);

INVxp33_ASAP7_75t_SL g1499 ( 
.A(n_727),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_990),
.Y(n_1500)
);

INVxp67_ASAP7_75t_SL g1501 ( 
.A(n_781),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_979),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_983),
.Y(n_1503)
);

INVxp67_ASAP7_75t_L g1504 ( 
.A(n_983),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_984),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_984),
.Y(n_1506)
);

INVxp33_ASAP7_75t_L g1507 ( 
.A(n_867),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_988),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_988),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_996),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_996),
.Y(n_1511)
);

INVxp67_ASAP7_75t_SL g1512 ( 
.A(n_781),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1002),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_981),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_728),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1002),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1012),
.Y(n_1517)
);

BUFx6f_ASAP7_75t_L g1518 ( 
.A(n_801),
.Y(n_1518)
);

INVxp67_ASAP7_75t_L g1519 ( 
.A(n_1012),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1018),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1018),
.Y(n_1521)
);

CKINVDCx16_ASAP7_75t_R g1522 ( 
.A(n_934),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1022),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1022),
.Y(n_1524)
);

INVxp33_ASAP7_75t_SL g1525 ( 
.A(n_734),
.Y(n_1525)
);

BUFx6f_ASAP7_75t_L g1526 ( 
.A(n_1125),
.Y(n_1526)
);

INVxp67_ASAP7_75t_L g1527 ( 
.A(n_1025),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1025),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1032),
.Y(n_1529)
);

INVxp33_ASAP7_75t_SL g1530 ( 
.A(n_735),
.Y(n_1530)
);

CKINVDCx16_ASAP7_75t_R g1531 ( 
.A(n_934),
.Y(n_1531)
);

CKINVDCx16_ASAP7_75t_R g1532 ( 
.A(n_952),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_990),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_736),
.Y(n_1534)
);

CKINVDCx20_ASAP7_75t_R g1535 ( 
.A(n_790),
.Y(n_1535)
);

CKINVDCx14_ASAP7_75t_R g1536 ( 
.A(n_717),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_739),
.Y(n_1537)
);

CKINVDCx20_ASAP7_75t_R g1538 ( 
.A(n_813),
.Y(n_1538)
);

INVxp33_ASAP7_75t_SL g1539 ( 
.A(n_740),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_741),
.Y(n_1540)
);

INVxp67_ASAP7_75t_SL g1541 ( 
.A(n_781),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1032),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_981),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1065),
.Y(n_1544)
);

CKINVDCx16_ASAP7_75t_R g1545 ( 
.A(n_952),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_742),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1065),
.Y(n_1547)
);

INVxp67_ASAP7_75t_L g1548 ( 
.A(n_1067),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1067),
.Y(n_1549)
);

CKINVDCx20_ASAP7_75t_R g1550 ( 
.A(n_835),
.Y(n_1550)
);

INVxp33_ASAP7_75t_L g1551 ( 
.A(n_867),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1071),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_866),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_745),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1071),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1075),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1075),
.Y(n_1557)
);

INVxp33_ASAP7_75t_SL g1558 ( 
.A(n_751),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1077),
.Y(n_1559)
);

BUFx5_ASAP7_75t_L g1560 ( 
.A(n_949),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1077),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1082),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_981),
.Y(n_1563)
);

INVxp33_ASAP7_75t_SL g1564 ( 
.A(n_753),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_981),
.Y(n_1565)
);

BUFx2_ASAP7_75t_L g1566 ( 
.A(n_754),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1082),
.Y(n_1567)
);

INVx2_ASAP7_75t_SL g1568 ( 
.A(n_952),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1087),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_755),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1087),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_726),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_843),
.Y(n_1573)
);

CKINVDCx16_ASAP7_75t_R g1574 ( 
.A(n_952),
.Y(n_1574)
);

CKINVDCx20_ASAP7_75t_R g1575 ( 
.A(n_860),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_756),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1090),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_757),
.Y(n_1578)
);

INVxp33_ASAP7_75t_L g1579 ( 
.A(n_872),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1090),
.Y(n_1580)
);

INVxp33_ASAP7_75t_SL g1581 ( 
.A(n_760),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1100),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1100),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_981),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1105),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1105),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_981),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1106),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_981),
.Y(n_1589)
);

INVxp33_ASAP7_75t_SL g1590 ( 
.A(n_761),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1106),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1114),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1109),
.Y(n_1593)
);

INVxp67_ASAP7_75t_L g1594 ( 
.A(n_1109),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1114),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_763),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_768),
.Y(n_1597)
);

INVxp67_ASAP7_75t_SL g1598 ( 
.A(n_781),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1113),
.Y(n_1599)
);

BUFx2_ASAP7_75t_L g1600 ( 
.A(n_769),
.Y(n_1600)
);

INVxp67_ASAP7_75t_SL g1601 ( 
.A(n_781),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1113),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1115),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_771),
.Y(n_1604)
);

CKINVDCx20_ASAP7_75t_R g1605 ( 
.A(n_912),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1115),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1116),
.Y(n_1607)
);

CKINVDCx20_ASAP7_75t_R g1608 ( 
.A(n_924),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1116),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1127),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1127),
.Y(n_1611)
);

BUFx3_ASAP7_75t_L g1612 ( 
.A(n_949),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1131),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_772),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1131),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_775),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1114),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1133),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1133),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_777),
.Y(n_1620)
);

CKINVDCx16_ASAP7_75t_R g1621 ( 
.A(n_973),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1137),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1137),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1114),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1138),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1138),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_779),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1140),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1140),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1141),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1141),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1142),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1142),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1145),
.Y(n_1634)
);

INVxp67_ASAP7_75t_SL g1635 ( 
.A(n_800),
.Y(n_1635)
);

CKINVDCx16_ASAP7_75t_R g1636 ( 
.A(n_973),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_782),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1145),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1153),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1153),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1154),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1154),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_784),
.Y(n_1643)
);

BUFx2_ASAP7_75t_SL g1644 ( 
.A(n_1054),
.Y(n_1644)
);

BUFx6f_ASAP7_75t_L g1645 ( 
.A(n_1125),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1160),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1160),
.Y(n_1647)
);

INVxp67_ASAP7_75t_L g1648 ( 
.A(n_1161),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_786),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1161),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1164),
.Y(n_1651)
);

CKINVDCx20_ASAP7_75t_R g1652 ( 
.A(n_948),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1164),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1167),
.Y(n_1654)
);

CKINVDCx20_ASAP7_75t_R g1655 ( 
.A(n_1014),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1167),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_789),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1172),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1172),
.Y(n_1659)
);

INVxp67_ASAP7_75t_L g1660 ( 
.A(n_1174),
.Y(n_1660)
);

INVxp67_ASAP7_75t_SL g1661 ( 
.A(n_800),
.Y(n_1661)
);

CKINVDCx20_ASAP7_75t_R g1662 ( 
.A(n_1033),
.Y(n_1662)
);

INVxp33_ASAP7_75t_L g1663 ( 
.A(n_872),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_792),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1174),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1176),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1176),
.Y(n_1667)
);

CKINVDCx20_ASAP7_75t_R g1668 ( 
.A(n_1043),
.Y(n_1668)
);

INVxp67_ASAP7_75t_SL g1669 ( 
.A(n_800),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_793),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1178),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1178),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1181),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1181),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_798),
.Y(n_1675)
);

INVxp33_ASAP7_75t_L g1676 ( 
.A(n_880),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1183),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1183),
.Y(n_1678)
);

INVxp67_ASAP7_75t_L g1679 ( 
.A(n_1192),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_802),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1192),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1193),
.Y(n_1682)
);

BUFx6f_ASAP7_75t_L g1683 ( 
.A(n_1125),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1193),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1200),
.Y(n_1685)
);

BUFx5_ASAP7_75t_L g1686 ( 
.A(n_970),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_804),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1200),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1201),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1201),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_805),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1205),
.Y(n_1692)
);

INVx3_ASAP7_75t_L g1693 ( 
.A(n_800),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1205),
.Y(n_1694)
);

INVxp67_ASAP7_75t_L g1695 ( 
.A(n_1206),
.Y(n_1695)
);

INVxp67_ASAP7_75t_SL g1696 ( 
.A(n_800),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1206),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_806),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1208),
.Y(n_1699)
);

INVxp67_ASAP7_75t_L g1700 ( 
.A(n_1208),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1212),
.Y(n_1701)
);

CKINVDCx16_ASAP7_75t_R g1702 ( 
.A(n_973),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1212),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_809),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1215),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1215),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1224),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1224),
.Y(n_1708)
);

BUFx6f_ASAP7_75t_L g1709 ( 
.A(n_1125),
.Y(n_1709)
);

INVxp67_ASAP7_75t_SL g1710 ( 
.A(n_891),
.Y(n_1710)
);

BUFx3_ASAP7_75t_L g1711 ( 
.A(n_970),
.Y(n_1711)
);

BUFx2_ASAP7_75t_L g1712 ( 
.A(n_811),
.Y(n_1712)
);

BUFx8_ASAP7_75t_SL g1713 ( 
.A(n_1403),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1398),
.B(n_1083),
.Y(n_1714)
);

BUFx6f_ASAP7_75t_L g1715 ( 
.A(n_1264),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1398),
.B(n_1083),
.Y(n_1716)
);

BUFx6f_ASAP7_75t_L g1717 ( 
.A(n_1264),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1494),
.B(n_1189),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1494),
.B(n_1189),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1306),
.B(n_973),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1644),
.B(n_1198),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1437),
.Y(n_1722)
);

INVx5_ASAP7_75t_L g1723 ( 
.A(n_1264),
.Y(n_1723)
);

INVx5_ASAP7_75t_L g1724 ( 
.A(n_1264),
.Y(n_1724)
);

INVx5_ASAP7_75t_L g1725 ( 
.A(n_1309),
.Y(n_1725)
);

INVxp33_ASAP7_75t_SL g1726 ( 
.A(n_1262),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1536),
.B(n_1198),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1304),
.B(n_1204),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1274),
.Y(n_1729)
);

INVx3_ASAP7_75t_L g1730 ( 
.A(n_1437),
.Y(n_1730)
);

AND2x4_ASAP7_75t_L g1731 ( 
.A(n_1373),
.B(n_1401),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1285),
.B(n_1089),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1338),
.B(n_1089),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1300),
.Y(n_1734)
);

BUFx6f_ASAP7_75t_L g1735 ( 
.A(n_1309),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1317),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1346),
.Y(n_1737)
);

INVx3_ASAP7_75t_L g1738 ( 
.A(n_1461),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1493),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1536),
.B(n_1204),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1274),
.Y(n_1741)
);

INVx3_ASAP7_75t_L g1742 ( 
.A(n_1461),
.Y(n_1742)
);

BUFx3_ASAP7_75t_L g1743 ( 
.A(n_1391),
.Y(n_1743)
);

BUFx2_ASAP7_75t_L g1744 ( 
.A(n_1297),
.Y(n_1744)
);

INVx4_ASAP7_75t_L g1745 ( 
.A(n_1390),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_1441),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1283),
.Y(n_1747)
);

AND2x4_ASAP7_75t_L g1748 ( 
.A(n_1568),
.B(n_744),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1413),
.B(n_1236),
.Y(n_1749)
);

INVx3_ASAP7_75t_L g1750 ( 
.A(n_1391),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1261),
.B(n_1236),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1276),
.B(n_1054),
.Y(n_1752)
);

INVx5_ASAP7_75t_L g1753 ( 
.A(n_1309),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1390),
.B(n_1081),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1283),
.Y(n_1755)
);

AND2x6_ASAP7_75t_L g1756 ( 
.A(n_1474),
.B(n_892),
.Y(n_1756)
);

NOR2x1_ASAP7_75t_L g1757 ( 
.A(n_1474),
.B(n_892),
.Y(n_1757)
);

BUFx3_ASAP7_75t_L g1758 ( 
.A(n_1693),
.Y(n_1758)
);

BUFx6f_ASAP7_75t_L g1759 ( 
.A(n_1309),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1453),
.B(n_1081),
.Y(n_1760)
);

INVx3_ASAP7_75t_L g1761 ( 
.A(n_1693),
.Y(n_1761)
);

BUFx3_ASAP7_75t_L g1762 ( 
.A(n_1289),
.Y(n_1762)
);

BUFx6f_ASAP7_75t_L g1763 ( 
.A(n_1339),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1453),
.B(n_1114),
.Y(n_1764)
);

INVx5_ASAP7_75t_L g1765 ( 
.A(n_1339),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1289),
.Y(n_1766)
);

INVx5_ASAP7_75t_L g1767 ( 
.A(n_1339),
.Y(n_1767)
);

AND2x4_ASAP7_75t_L g1768 ( 
.A(n_1472),
.B(n_749),
.Y(n_1768)
);

BUFx8_ASAP7_75t_SL g1769 ( 
.A(n_1403),
.Y(n_1769)
);

BUFx6f_ASAP7_75t_L g1770 ( 
.A(n_1339),
.Y(n_1770)
);

BUFx6f_ASAP7_75t_L g1771 ( 
.A(n_1407),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1313),
.Y(n_1772)
);

INVx5_ASAP7_75t_L g1773 ( 
.A(n_1407),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1466),
.B(n_1114),
.Y(n_1774)
);

BUFx6f_ASAP7_75t_L g1775 ( 
.A(n_1407),
.Y(n_1775)
);

BUFx12f_ASAP7_75t_L g1776 ( 
.A(n_1279),
.Y(n_1776)
);

INVx4_ASAP7_75t_L g1777 ( 
.A(n_1466),
.Y(n_1777)
);

INVx3_ASAP7_75t_L g1778 ( 
.A(n_1553),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1354),
.B(n_1388),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1313),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1500),
.B(n_1114),
.Y(n_1781)
);

BUFx12f_ASAP7_75t_L g1782 ( 
.A(n_1280),
.Y(n_1782)
);

INVx5_ASAP7_75t_L g1783 ( 
.A(n_1407),
.Y(n_1783)
);

INVx5_ASAP7_75t_L g1784 ( 
.A(n_1518),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1354),
.B(n_1089),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1500),
.B(n_1114),
.Y(n_1786)
);

CKINVDCx16_ASAP7_75t_R g1787 ( 
.A(n_1454),
.Y(n_1787)
);

BUFx6f_ASAP7_75t_L g1788 ( 
.A(n_1518),
.Y(n_1788)
);

INVx5_ASAP7_75t_L g1789 ( 
.A(n_1518),
.Y(n_1789)
);

BUFx2_ASAP7_75t_L g1790 ( 
.A(n_1298),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1501),
.Y(n_1791)
);

BUFx8_ASAP7_75t_SL g1792 ( 
.A(n_1409),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1533),
.B(n_1114),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1533),
.B(n_998),
.Y(n_1794)
);

BUFx6f_ASAP7_75t_L g1795 ( 
.A(n_1518),
.Y(n_1795)
);

INVx5_ASAP7_75t_L g1796 ( 
.A(n_1526),
.Y(n_1796)
);

BUFx8_ASAP7_75t_SL g1797 ( 
.A(n_1409),
.Y(n_1797)
);

AND2x6_ASAP7_75t_L g1798 ( 
.A(n_1553),
.B(n_998),
.Y(n_1798)
);

BUFx12f_ASAP7_75t_L g1799 ( 
.A(n_1262),
.Y(n_1799)
);

BUFx6f_ASAP7_75t_L g1800 ( 
.A(n_1526),
.Y(n_1800)
);

BUFx2_ASAP7_75t_L g1801 ( 
.A(n_1305),
.Y(n_1801)
);

INVx4_ASAP7_75t_L g1802 ( 
.A(n_1526),
.Y(n_1802)
);

BUFx3_ASAP7_75t_L g1803 ( 
.A(n_1324),
.Y(n_1803)
);

BUFx8_ASAP7_75t_SL g1804 ( 
.A(n_1421),
.Y(n_1804)
);

INVx6_ASAP7_75t_L g1805 ( 
.A(n_1612),
.Y(n_1805)
);

BUFx3_ASAP7_75t_L g1806 ( 
.A(n_1324),
.Y(n_1806)
);

AND2x4_ASAP7_75t_L g1807 ( 
.A(n_1566),
.B(n_749),
.Y(n_1807)
);

BUFx3_ASAP7_75t_L g1808 ( 
.A(n_1327),
.Y(n_1808)
);

INVx3_ASAP7_75t_L g1809 ( 
.A(n_1612),
.Y(n_1809)
);

CKINVDCx16_ASAP7_75t_R g1810 ( 
.A(n_1467),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1512),
.Y(n_1811)
);

BUFx6f_ASAP7_75t_L g1812 ( 
.A(n_1526),
.Y(n_1812)
);

BUFx6f_ASAP7_75t_L g1813 ( 
.A(n_1645),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1541),
.B(n_719),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1327),
.Y(n_1815)
);

BUFx2_ASAP7_75t_L g1816 ( 
.A(n_1386),
.Y(n_1816)
);

BUFx12f_ASAP7_75t_L g1817 ( 
.A(n_1322),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1598),
.Y(n_1818)
);

AND2x4_ASAP7_75t_L g1819 ( 
.A(n_1600),
.B(n_845),
.Y(n_1819)
);

INVx5_ASAP7_75t_L g1820 ( 
.A(n_1645),
.Y(n_1820)
);

CKINVDCx11_ASAP7_75t_R g1821 ( 
.A(n_1265),
.Y(n_1821)
);

INVx4_ASAP7_75t_L g1822 ( 
.A(n_1645),
.Y(n_1822)
);

INVx5_ASAP7_75t_L g1823 ( 
.A(n_1645),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_SL g1824 ( 
.A(n_1304),
.B(n_891),
.Y(n_1824)
);

INVx3_ASAP7_75t_L g1825 ( 
.A(n_1711),
.Y(n_1825)
);

INVx4_ASAP7_75t_L g1826 ( 
.A(n_1683),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_L g1827 ( 
.A(n_1301),
.B(n_891),
.Y(n_1827)
);

INVx5_ASAP7_75t_L g1828 ( 
.A(n_1683),
.Y(n_1828)
);

AND2x4_ASAP7_75t_L g1829 ( 
.A(n_1712),
.B(n_845),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1281),
.B(n_887),
.Y(n_1830)
);

INVx5_ASAP7_75t_L g1831 ( 
.A(n_1683),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_SL g1832 ( 
.A(n_1382),
.B(n_1089),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1388),
.B(n_1107),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1601),
.B(n_738),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1330),
.Y(n_1835)
);

AND2x4_ASAP7_75t_L g1836 ( 
.A(n_1282),
.B(n_887),
.Y(n_1836)
);

NOR2x1_ASAP7_75t_L g1837 ( 
.A(n_1711),
.B(n_1125),
.Y(n_1837)
);

AND2x4_ASAP7_75t_L g1838 ( 
.A(n_1284),
.B(n_900),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1635),
.B(n_748),
.Y(n_1839)
);

AND2x4_ASAP7_75t_L g1840 ( 
.A(n_1287),
.B(n_900),
.Y(n_1840)
);

NOR2xp33_ASAP7_75t_SL g1841 ( 
.A(n_1483),
.B(n_1107),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1661),
.B(n_750),
.Y(n_1842)
);

BUFx6f_ASAP7_75t_L g1843 ( 
.A(n_1683),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1669),
.B(n_758),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1330),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1434),
.B(n_1107),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1348),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1348),
.Y(n_1848)
);

BUFx3_ASAP7_75t_L g1849 ( 
.A(n_1365),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1696),
.B(n_1710),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1293),
.B(n_780),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1365),
.Y(n_1852)
);

INVx3_ASAP7_75t_L g1853 ( 
.A(n_1263),
.Y(n_1853)
);

BUFx6f_ASAP7_75t_L g1854 ( 
.A(n_1709),
.Y(n_1854)
);

BUFx6f_ASAP7_75t_L g1855 ( 
.A(n_1709),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1293),
.B(n_807),
.Y(n_1856)
);

INVx3_ASAP7_75t_L g1857 ( 
.A(n_1266),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1296),
.Y(n_1858)
);

BUFx3_ASAP7_75t_L g1859 ( 
.A(n_1367),
.Y(n_1859)
);

BUFx3_ASAP7_75t_L g1860 ( 
.A(n_1367),
.Y(n_1860)
);

BUFx6f_ASAP7_75t_L g1861 ( 
.A(n_1709),
.Y(n_1861)
);

HB1xp67_ASAP7_75t_L g1862 ( 
.A(n_1332),
.Y(n_1862)
);

INVx2_ASAP7_75t_SL g1863 ( 
.A(n_1578),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1293),
.B(n_822),
.Y(n_1864)
);

BUFx6f_ASAP7_75t_L g1865 ( 
.A(n_1709),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1293),
.B(n_824),
.Y(n_1866)
);

BUFx6f_ASAP7_75t_L g1867 ( 
.A(n_1468),
.Y(n_1867)
);

INVx5_ASAP7_75t_L g1868 ( 
.A(n_1468),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1293),
.B(n_825),
.Y(n_1869)
);

NOR2xp33_ASAP7_75t_SL g1870 ( 
.A(n_1497),
.B(n_1522),
.Y(n_1870)
);

INVx5_ASAP7_75t_L g1871 ( 
.A(n_1514),
.Y(n_1871)
);

HB1xp67_ASAP7_75t_L g1872 ( 
.A(n_1420),
.Y(n_1872)
);

BUFx12f_ASAP7_75t_L g1873 ( 
.A(n_1322),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1514),
.Y(n_1874)
);

INVx5_ASAP7_75t_L g1875 ( 
.A(n_1543),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1299),
.Y(n_1876)
);

INVx2_ASAP7_75t_SL g1877 ( 
.A(n_1596),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1293),
.B(n_886),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1302),
.Y(n_1879)
);

AND2x4_ASAP7_75t_L g1880 ( 
.A(n_1288),
.B(n_1152),
.Y(n_1880)
);

INVx4_ASAP7_75t_L g1881 ( 
.A(n_1604),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1303),
.Y(n_1882)
);

INVx5_ASAP7_75t_L g1883 ( 
.A(n_1543),
.Y(n_1883)
);

AND2x4_ASAP7_75t_L g1884 ( 
.A(n_1290),
.B(n_1152),
.Y(n_1884)
);

BUFx8_ASAP7_75t_L g1885 ( 
.A(n_1286),
.Y(n_1885)
);

AND2x4_ASAP7_75t_L g1886 ( 
.A(n_1294),
.B(n_1239),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1434),
.B(n_1107),
.Y(n_1887)
);

INVx5_ASAP7_75t_L g1888 ( 
.A(n_1563),
.Y(n_1888)
);

HB1xp67_ASAP7_75t_L g1889 ( 
.A(n_1292),
.Y(n_1889)
);

AND2x6_ASAP7_75t_L g1890 ( 
.A(n_1563),
.B(n_1255),
.Y(n_1890)
);

AND2x4_ASAP7_75t_L g1891 ( 
.A(n_1314),
.B(n_1239),
.Y(n_1891)
);

BUFx6f_ASAP7_75t_L g1892 ( 
.A(n_1565),
.Y(n_1892)
);

NOR2xp33_ASAP7_75t_L g1893 ( 
.A(n_1444),
.B(n_891),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1307),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1565),
.Y(n_1895)
);

INVx5_ASAP7_75t_L g1896 ( 
.A(n_1584),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1291),
.B(n_1254),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1444),
.B(n_1197),
.Y(n_1898)
);

BUFx2_ASAP7_75t_L g1899 ( 
.A(n_1265),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1293),
.B(n_903),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1584),
.Y(n_1901)
);

BUFx6f_ASAP7_75t_L g1902 ( 
.A(n_1587),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1357),
.B(n_911),
.Y(n_1903)
);

AND2x4_ASAP7_75t_L g1904 ( 
.A(n_1515),
.B(n_1245),
.Y(n_1904)
);

BUFx2_ASAP7_75t_L g1905 ( 
.A(n_1295),
.Y(n_1905)
);

BUFx12f_ASAP7_75t_L g1906 ( 
.A(n_1325),
.Y(n_1906)
);

BUFx6f_ASAP7_75t_L g1907 ( 
.A(n_1587),
.Y(n_1907)
);

AND2x4_ASAP7_75t_L g1908 ( 
.A(n_1554),
.B(n_1245),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1589),
.Y(n_1909)
);

INVx5_ASAP7_75t_L g1910 ( 
.A(n_1589),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1357),
.B(n_914),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1310),
.Y(n_1912)
);

NAND2x1_ASAP7_75t_L g1913 ( 
.A(n_1267),
.B(n_891),
.Y(n_1913)
);

INVx3_ASAP7_75t_L g1914 ( 
.A(n_1268),
.Y(n_1914)
);

BUFx6f_ASAP7_75t_L g1915 ( 
.A(n_1592),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1592),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1357),
.B(n_920),
.Y(n_1917)
);

BUFx8_ASAP7_75t_SL g1918 ( 
.A(n_1421),
.Y(n_1918)
);

BUFx6f_ASAP7_75t_L g1919 ( 
.A(n_1595),
.Y(n_1919)
);

NOR2xp33_ASAP7_75t_SL g1920 ( 
.A(n_1531),
.B(n_1197),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1312),
.Y(n_1921)
);

INVx5_ASAP7_75t_L g1922 ( 
.A(n_1595),
.Y(n_1922)
);

INVxp67_ASAP7_75t_L g1923 ( 
.A(n_1576),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1357),
.B(n_922),
.Y(n_1924)
);

NOR2xp33_ASAP7_75t_L g1925 ( 
.A(n_1459),
.B(n_902),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1417),
.Y(n_1926)
);

BUFx12f_ASAP7_75t_L g1927 ( 
.A(n_1325),
.Y(n_1927)
);

BUFx6f_ASAP7_75t_L g1928 ( 
.A(n_1617),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1617),
.Y(n_1929)
);

BUFx2_ASAP7_75t_L g1930 ( 
.A(n_1295),
.Y(n_1930)
);

INVx5_ASAP7_75t_L g1931 ( 
.A(n_1624),
.Y(n_1931)
);

BUFx6f_ASAP7_75t_L g1932 ( 
.A(n_1624),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1357),
.B(n_946),
.Y(n_1933)
);

INVx5_ASAP7_75t_L g1934 ( 
.A(n_1532),
.Y(n_1934)
);

HB1xp67_ASAP7_75t_L g1935 ( 
.A(n_1614),
.Y(n_1935)
);

BUFx12f_ASAP7_75t_L g1936 ( 
.A(n_1446),
.Y(n_1936)
);

BUFx6f_ASAP7_75t_L g1937 ( 
.A(n_1315),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1459),
.B(n_902),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1357),
.Y(n_1939)
);

AND2x4_ASAP7_75t_L g1940 ( 
.A(n_1597),
.B(n_880),
.Y(n_1940)
);

INVx2_ASAP7_75t_SL g1941 ( 
.A(n_1620),
.Y(n_1941)
);

BUFx3_ASAP7_75t_L g1942 ( 
.A(n_1270),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_SL g1943 ( 
.A(n_1311),
.B(n_902),
.Y(n_1943)
);

INVx5_ASAP7_75t_L g1944 ( 
.A(n_1545),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1357),
.B(n_1560),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1560),
.B(n_1005),
.Y(n_1946)
);

INVx5_ASAP7_75t_L g1947 ( 
.A(n_1574),
.Y(n_1947)
);

INVx3_ASAP7_75t_L g1948 ( 
.A(n_1271),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1462),
.B(n_1197),
.Y(n_1949)
);

INVx3_ASAP7_75t_L g1950 ( 
.A(n_1272),
.Y(n_1950)
);

INVx5_ASAP7_75t_L g1951 ( 
.A(n_1621),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1560),
.Y(n_1952)
);

BUFx12f_ASAP7_75t_L g1953 ( 
.A(n_1447),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1560),
.B(n_1030),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1318),
.Y(n_1955)
);

BUFx6f_ASAP7_75t_L g1956 ( 
.A(n_1320),
.Y(n_1956)
);

INVx4_ASAP7_75t_L g1957 ( 
.A(n_1627),
.Y(n_1957)
);

HB1xp67_ASAP7_75t_L g1958 ( 
.A(n_1637),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1462),
.B(n_1197),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1560),
.B(n_1686),
.Y(n_1960)
);

BUFx3_ASAP7_75t_L g1961 ( 
.A(n_1273),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1507),
.B(n_1216),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1560),
.B(n_1031),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1507),
.B(n_1216),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1551),
.B(n_1216),
.Y(n_1965)
);

BUFx12f_ASAP7_75t_L g1966 ( 
.A(n_1643),
.Y(n_1966)
);

BUFx12f_ASAP7_75t_L g1967 ( 
.A(n_1649),
.Y(n_1967)
);

NOR2xp33_ASAP7_75t_L g1968 ( 
.A(n_1551),
.B(n_902),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1323),
.Y(n_1969)
);

INVx4_ASAP7_75t_L g1970 ( 
.A(n_1675),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1579),
.B(n_1216),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1326),
.Y(n_1972)
);

BUFx6f_ASAP7_75t_L g1973 ( 
.A(n_1328),
.Y(n_1973)
);

BUFx3_ASAP7_75t_L g1974 ( 
.A(n_1275),
.Y(n_1974)
);

HB1xp67_ASAP7_75t_L g1975 ( 
.A(n_1698),
.Y(n_1975)
);

INVx4_ASAP7_75t_L g1976 ( 
.A(n_1534),
.Y(n_1976)
);

BUFx6f_ASAP7_75t_L g1977 ( 
.A(n_1329),
.Y(n_1977)
);

BUFx8_ASAP7_75t_SL g1978 ( 
.A(n_1535),
.Y(n_1978)
);

BUFx6f_ASAP7_75t_L g1979 ( 
.A(n_1331),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_SL g1980 ( 
.A(n_1636),
.B(n_1157),
.Y(n_1980)
);

BUFx12f_ASAP7_75t_L g1981 ( 
.A(n_1534),
.Y(n_1981)
);

BUFx6f_ASAP7_75t_L g1982 ( 
.A(n_1333),
.Y(n_1982)
);

AND2x6_ASAP7_75t_L g1983 ( 
.A(n_1366),
.B(n_1255),
.Y(n_1983)
);

BUFx6f_ASAP7_75t_L g1984 ( 
.A(n_1335),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1560),
.B(n_1060),
.Y(n_1985)
);

BUFx3_ASAP7_75t_L g1986 ( 
.A(n_1278),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1336),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1579),
.B(n_909),
.Y(n_1988)
);

INVx4_ASAP7_75t_L g1989 ( 
.A(n_1537),
.Y(n_1989)
);

NAND2xp33_ASAP7_75t_L g1990 ( 
.A(n_1686),
.B(n_902),
.Y(n_1990)
);

BUFx12f_ASAP7_75t_L g1991 ( 
.A(n_1537),
.Y(n_1991)
);

BUFx6f_ASAP7_75t_L g1992 ( 
.A(n_1337),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1686),
.B(n_1074),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1663),
.B(n_909),
.Y(n_1994)
);

CKINVDCx5p33_ASAP7_75t_R g1995 ( 
.A(n_1319),
.Y(n_1995)
);

INVx5_ASAP7_75t_L g1996 ( 
.A(n_1702),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1340),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1341),
.Y(n_1998)
);

INVx3_ASAP7_75t_L g1999 ( 
.A(n_1342),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1663),
.B(n_967),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_SL g2001 ( 
.A(n_1366),
.B(n_918),
.Y(n_2001)
);

BUFx6f_ASAP7_75t_L g2002 ( 
.A(n_1343),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1686),
.B(n_1084),
.Y(n_2003)
);

AND2x4_ASAP7_75t_L g2004 ( 
.A(n_1616),
.B(n_967),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1676),
.B(n_980),
.Y(n_2005)
);

INVx2_ASAP7_75t_SL g2006 ( 
.A(n_1540),
.Y(n_2006)
);

CKINVDCx5p33_ASAP7_75t_R g2007 ( 
.A(n_1389),
.Y(n_2007)
);

INVx5_ASAP7_75t_L g2008 ( 
.A(n_1686),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1676),
.B(n_980),
.Y(n_2009)
);

AND2x4_ASAP7_75t_L g2010 ( 
.A(n_1657),
.B(n_991),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1686),
.B(n_1185),
.Y(n_2011)
);

BUFx6f_ASAP7_75t_L g2012 ( 
.A(n_1344),
.Y(n_2012)
);

NOR2xp33_ASAP7_75t_L g2013 ( 
.A(n_1670),
.B(n_918),
.Y(n_2013)
);

NOR2xp33_ASAP7_75t_L g2014 ( 
.A(n_1680),
.B(n_918),
.Y(n_2014)
);

INVx5_ASAP7_75t_L g2015 ( 
.A(n_1686),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1345),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1316),
.B(n_1199),
.Y(n_2017)
);

AND2x4_ASAP7_75t_L g2018 ( 
.A(n_1334),
.B(n_991),
.Y(n_2018)
);

BUFx12f_ASAP7_75t_L g2019 ( 
.A(n_1540),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_SL g2020 ( 
.A(n_1393),
.B(n_918),
.Y(n_2020)
);

NOR2xp33_ASAP7_75t_SL g2021 ( 
.A(n_1368),
.B(n_1080),
.Y(n_2021)
);

AND2x4_ASAP7_75t_L g2022 ( 
.A(n_1370),
.B(n_1016),
.Y(n_2022)
);

INVxp67_ASAP7_75t_L g2023 ( 
.A(n_1546),
.Y(n_2023)
);

INVx5_ASAP7_75t_L g2024 ( 
.A(n_1393),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1347),
.Y(n_2025)
);

INVx5_ASAP7_75t_L g2026 ( 
.A(n_1387),
.Y(n_2026)
);

INVx2_ASAP7_75t_SL g2027 ( 
.A(n_1546),
.Y(n_2027)
);

INVx5_ASAP7_75t_L g2028 ( 
.A(n_1431),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1349),
.Y(n_2029)
);

NOR2xp33_ASAP7_75t_L g2030 ( 
.A(n_1368),
.B(n_918),
.Y(n_2030)
);

INVx5_ASAP7_75t_L g2031 ( 
.A(n_1442),
.Y(n_2031)
);

NOR2xp33_ASAP7_75t_L g2032 ( 
.A(n_1378),
.B(n_1180),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1350),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1269),
.B(n_1016),
.Y(n_2034)
);

INVx3_ASAP7_75t_L g2035 ( 
.A(n_1351),
.Y(n_2035)
);

AND2x4_ASAP7_75t_L g2036 ( 
.A(n_1448),
.B(n_1059),
.Y(n_2036)
);

INVx5_ASAP7_75t_L g2037 ( 
.A(n_1487),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1504),
.B(n_1240),
.Y(n_2038)
);

BUFx6f_ASAP7_75t_L g2039 ( 
.A(n_1352),
.Y(n_2039)
);

AND2x4_ASAP7_75t_L g2040 ( 
.A(n_1519),
.B(n_1059),
.Y(n_2040)
);

INVx2_ASAP7_75t_SL g2041 ( 
.A(n_1570),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1527),
.B(n_1548),
.Y(n_2042)
);

BUFx6f_ASAP7_75t_L g2043 ( 
.A(n_1353),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1269),
.B(n_1096),
.Y(n_2044)
);

AND2x6_ASAP7_75t_L g2045 ( 
.A(n_1708),
.B(n_1096),
.Y(n_2045)
);

INVx5_ASAP7_75t_L g2046 ( 
.A(n_1594),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1355),
.Y(n_2047)
);

BUFx6f_ASAP7_75t_L g2048 ( 
.A(n_1356),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1360),
.Y(n_2049)
);

CKINVDCx5p33_ASAP7_75t_R g2050 ( 
.A(n_1427),
.Y(n_2050)
);

INVx3_ASAP7_75t_L g2051 ( 
.A(n_1361),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1570),
.B(n_1664),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1362),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1364),
.Y(n_2054)
);

AND2x6_ASAP7_75t_L g2055 ( 
.A(n_1707),
.B(n_1099),
.Y(n_2055)
);

INVx3_ASAP7_75t_L g2056 ( 
.A(n_1369),
.Y(n_2056)
);

AND2x4_ASAP7_75t_L g2057 ( 
.A(n_1638),
.B(n_1099),
.Y(n_2057)
);

BUFx12f_ASAP7_75t_L g2058 ( 
.A(n_1664),
.Y(n_2058)
);

INVx5_ASAP7_75t_L g2059 ( 
.A(n_1648),
.Y(n_2059)
);

BUFx6f_ASAP7_75t_L g2060 ( 
.A(n_1371),
.Y(n_2060)
);

BUFx6f_ASAP7_75t_L g2061 ( 
.A(n_1372),
.Y(n_2061)
);

INVx5_ASAP7_75t_L g2062 ( 
.A(n_1660),
.Y(n_2062)
);

HB1xp67_ASAP7_75t_L g2063 ( 
.A(n_1687),
.Y(n_2063)
);

INVx5_ASAP7_75t_L g2064 ( 
.A(n_1679),
.Y(n_2064)
);

AND2x4_ASAP7_75t_L g2065 ( 
.A(n_1695),
.B(n_1118),
.Y(n_2065)
);

BUFx6f_ASAP7_75t_L g2066 ( 
.A(n_1374),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1687),
.B(n_1691),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_1691),
.B(n_1704),
.Y(n_2068)
);

INVx3_ASAP7_75t_L g2069 ( 
.A(n_1376),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1700),
.B(n_1180),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_SL g2071 ( 
.A(n_1704),
.B(n_1180),
.Y(n_2071)
);

NOR2xp33_ASAP7_75t_L g2072 ( 
.A(n_1378),
.B(n_1180),
.Y(n_2072)
);

INVx5_ASAP7_75t_L g2073 ( 
.A(n_1377),
.Y(n_2073)
);

BUFx6f_ASAP7_75t_L g2074 ( 
.A(n_1379),
.Y(n_2074)
);

BUFx6f_ASAP7_75t_L g2075 ( 
.A(n_1380),
.Y(n_2075)
);

BUFx12f_ASAP7_75t_L g2076 ( 
.A(n_1572),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1381),
.Y(n_2077)
);

AND2x4_ASAP7_75t_L g2078 ( 
.A(n_1383),
.B(n_1118),
.Y(n_2078)
);

BUFx2_ASAP7_75t_L g2079 ( 
.A(n_1308),
.Y(n_2079)
);

OR2x6_ASAP7_75t_L g2080 ( 
.A(n_1359),
.B(n_731),
.Y(n_2080)
);

AND2x4_ASAP7_75t_L g2081 ( 
.A(n_1384),
.B(n_1134),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2016),
.Y(n_2082)
);

BUFx2_ASAP7_75t_L g2083 ( 
.A(n_1926),
.Y(n_2083)
);

CKINVDCx5p33_ASAP7_75t_R g2084 ( 
.A(n_1966),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1778),
.B(n_1415),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2016),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1729),
.Y(n_2087)
);

AND2x4_ASAP7_75t_L g2088 ( 
.A(n_1722),
.B(n_1685),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1729),
.Y(n_2089)
);

INVx4_ASAP7_75t_L g2090 ( 
.A(n_2008),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2025),
.Y(n_2091)
);

HB1xp67_ASAP7_75t_L g2092 ( 
.A(n_1862),
.Y(n_2092)
);

NOR2xp33_ASAP7_75t_L g2093 ( 
.A(n_1794),
.B(n_1415),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2025),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2029),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_1741),
.Y(n_2096)
);

BUFx3_ASAP7_75t_L g2097 ( 
.A(n_1762),
.Y(n_2097)
);

INVx3_ASAP7_75t_L g2098 ( 
.A(n_1743),
.Y(n_2098)
);

INVx3_ASAP7_75t_L g2099 ( 
.A(n_1743),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2029),
.Y(n_2100)
);

BUFx6f_ASAP7_75t_L g2101 ( 
.A(n_1867),
.Y(n_2101)
);

AND2x4_ASAP7_75t_L g2102 ( 
.A(n_1722),
.B(n_1689),
.Y(n_2102)
);

BUFx6f_ASAP7_75t_L g2103 ( 
.A(n_1867),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2033),
.Y(n_2104)
);

NOR2xp67_ASAP7_75t_L g2105 ( 
.A(n_1934),
.B(n_1573),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1741),
.Y(n_2106)
);

OA21x2_ASAP7_75t_L g2107 ( 
.A1(n_1747),
.A2(n_1392),
.B(n_1385),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1747),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2033),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_1778),
.B(n_1449),
.Y(n_2110)
);

AND2x4_ASAP7_75t_L g2111 ( 
.A(n_1730),
.B(n_1697),
.Y(n_2111)
);

INVx3_ASAP7_75t_L g2112 ( 
.A(n_1758),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2053),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_1779),
.B(n_1308),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_1755),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2053),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1755),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2077),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1766),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2077),
.Y(n_2120)
);

BUFx6f_ASAP7_75t_L g2121 ( 
.A(n_1867),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1809),
.B(n_1449),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_SL g2123 ( 
.A(n_2024),
.B(n_1485),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1750),
.Y(n_2124)
);

CKINVDCx5p33_ASAP7_75t_R g2125 ( 
.A(n_1966),
.Y(n_2125)
);

NAND3xp33_ASAP7_75t_L g2126 ( 
.A(n_1728),
.B(n_814),
.C(n_812),
.Y(n_2126)
);

BUFx3_ASAP7_75t_L g2127 ( 
.A(n_1762),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1750),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1761),
.Y(n_2129)
);

INVx3_ASAP7_75t_L g2130 ( 
.A(n_1758),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_SL g2131 ( 
.A(n_2024),
.B(n_1485),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_1809),
.B(n_1495),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1761),
.Y(n_2133)
);

HB1xp67_ASAP7_75t_L g2134 ( 
.A(n_1862),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_1785),
.B(n_1321),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1937),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1937),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1937),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_1833),
.B(n_1321),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1937),
.Y(n_2140)
);

NOR2xp33_ASAP7_75t_L g2141 ( 
.A(n_1730),
.B(n_1495),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1956),
.Y(n_2142)
);

HB1xp67_ASAP7_75t_L g2143 ( 
.A(n_1872),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_1846),
.B(n_1358),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_1956),
.Y(n_2145)
);

INVx3_ASAP7_75t_L g2146 ( 
.A(n_1956),
.Y(n_2146)
);

INVx5_ASAP7_75t_L g2147 ( 
.A(n_1890),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1956),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_1887),
.B(n_1358),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1973),
.Y(n_2150)
);

NAND2x1_ASAP7_75t_L g2151 ( 
.A(n_1805),
.B(n_1180),
.Y(n_2151)
);

INVx4_ASAP7_75t_L g2152 ( 
.A(n_2008),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1973),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_SL g2154 ( 
.A(n_2024),
.B(n_1745),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1973),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_1766),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1973),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_1772),
.Y(n_2158)
);

OA21x2_ASAP7_75t_L g2159 ( 
.A1(n_1772),
.A2(n_1815),
.B(n_1780),
.Y(n_2159)
);

AND2x4_ASAP7_75t_L g2160 ( 
.A(n_1738),
.B(n_1681),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_1780),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_1898),
.B(n_1363),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1815),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_1949),
.B(n_1363),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1835),
.Y(n_2165)
);

BUFx6f_ASAP7_75t_L g2166 ( 
.A(n_1867),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1977),
.Y(n_2167)
);

HB1xp67_ASAP7_75t_L g2168 ( 
.A(n_1872),
.Y(n_2168)
);

BUFx6f_ASAP7_75t_L g2169 ( 
.A(n_1892),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_1835),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_1959),
.B(n_1397),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1845),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_1845),
.Y(n_2173)
);

NAND2x1p5_ASAP7_75t_L g2174 ( 
.A(n_1934),
.B(n_1394),
.Y(n_2174)
);

AOI22xp5_ASAP7_75t_L g2175 ( 
.A1(n_1728),
.A2(n_1277),
.B1(n_1525),
.B2(n_1499),
.Y(n_2175)
);

AND2x4_ASAP7_75t_L g2176 ( 
.A(n_1738),
.B(n_1742),
.Y(n_2176)
);

HB1xp67_ASAP7_75t_L g2177 ( 
.A(n_1889),
.Y(n_2177)
);

INVx3_ASAP7_75t_L g2178 ( 
.A(n_1977),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1977),
.Y(n_2179)
);

INVx3_ASAP7_75t_L g2180 ( 
.A(n_1803),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1977),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1979),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1979),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1979),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1979),
.Y(n_2185)
);

OAI21x1_ASAP7_75t_L g2186 ( 
.A1(n_1945),
.A2(n_1960),
.B(n_1952),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_SL g2187 ( 
.A(n_2024),
.B(n_1499),
.Y(n_2187)
);

NAND2xp33_ASAP7_75t_L g2188 ( 
.A(n_1983),
.B(n_1226),
.Y(n_2188)
);

AND2x4_ASAP7_75t_L g2189 ( 
.A(n_1742),
.B(n_1690),
.Y(n_2189)
);

AND2x4_ASAP7_75t_L g2190 ( 
.A(n_1825),
.B(n_1692),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1982),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1982),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_1847),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_1825),
.B(n_1525),
.Y(n_2194)
);

NOR2xp33_ASAP7_75t_L g2195 ( 
.A(n_1714),
.B(n_1530),
.Y(n_2195)
);

INVx3_ASAP7_75t_L g2196 ( 
.A(n_1803),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_1962),
.B(n_1397),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_1964),
.B(n_1395),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1982),
.Y(n_2199)
);

OAI21x1_ASAP7_75t_L g2200 ( 
.A1(n_1939),
.A2(n_1399),
.B(n_1396),
.Y(n_2200)
);

BUFx2_ASAP7_75t_L g2201 ( 
.A(n_1926),
.Y(n_2201)
);

OR2x6_ASAP7_75t_L g2202 ( 
.A(n_1776),
.B(n_1405),
.Y(n_2202)
);

BUFx6f_ASAP7_75t_L g2203 ( 
.A(n_1892),
.Y(n_2203)
);

HB1xp67_ASAP7_75t_L g2204 ( 
.A(n_1889),
.Y(n_2204)
);

INVx3_ASAP7_75t_L g2205 ( 
.A(n_1806),
.Y(n_2205)
);

HB1xp67_ASAP7_75t_L g2206 ( 
.A(n_2042),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_1716),
.B(n_1530),
.Y(n_2207)
);

BUFx2_ASAP7_75t_L g2208 ( 
.A(n_2050),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_1847),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_1848),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1982),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_1718),
.B(n_1539),
.Y(n_2212)
);

BUFx3_ASAP7_75t_L g2213 ( 
.A(n_1806),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_1719),
.B(n_1539),
.Y(n_2214)
);

BUFx6f_ASAP7_75t_L g2215 ( 
.A(n_1892),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_1965),
.B(n_1400),
.Y(n_2216)
);

BUFx3_ASAP7_75t_L g2217 ( 
.A(n_1808),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1984),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1984),
.Y(n_2219)
);

NOR2xp33_ASAP7_75t_L g2220 ( 
.A(n_1734),
.B(n_1558),
.Y(n_2220)
);

BUFx6f_ASAP7_75t_L g2221 ( 
.A(n_1892),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1984),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_2030),
.B(n_2032),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1984),
.Y(n_2224)
);

BUFx2_ASAP7_75t_L g2225 ( 
.A(n_2050),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_1848),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1992),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_SL g2228 ( 
.A(n_1745),
.B(n_1777),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_1852),
.Y(n_2229)
);

AND2x6_ASAP7_75t_L g2230 ( 
.A(n_1733),
.B(n_1134),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_1852),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_SL g2232 ( 
.A(n_1777),
.B(n_1558),
.Y(n_2232)
);

NOR2xp33_ASAP7_75t_SL g2233 ( 
.A(n_1841),
.B(n_1564),
.Y(n_2233)
);

BUFx6f_ASAP7_75t_L g2234 ( 
.A(n_1902),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_1874),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_2030),
.B(n_1564),
.Y(n_2236)
);

BUFx6f_ASAP7_75t_L g2237 ( 
.A(n_1902),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_1992),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1992),
.Y(n_2239)
);

AND2x2_ASAP7_75t_L g2240 ( 
.A(n_1971),
.B(n_1402),
.Y(n_2240)
);

INVx6_ASAP7_75t_L g2241 ( 
.A(n_1805),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_1874),
.Y(n_2242)
);

INVx5_ASAP7_75t_L g2243 ( 
.A(n_1890),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_1895),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_1895),
.Y(n_2245)
);

INVx3_ASAP7_75t_L g2246 ( 
.A(n_1992),
.Y(n_2246)
);

NOR2xp33_ASAP7_75t_L g2247 ( 
.A(n_1736),
.B(n_1581),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_2032),
.B(n_2072),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2002),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2002),
.Y(n_2250)
);

INVxp67_ASAP7_75t_L g2251 ( 
.A(n_1732),
.Y(n_2251)
);

AND2x2_ASAP7_75t_L g2252 ( 
.A(n_1988),
.B(n_1404),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_1901),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2002),
.Y(n_2254)
);

INVx2_ASAP7_75t_L g2255 ( 
.A(n_1901),
.Y(n_2255)
);

BUFx8_ASAP7_75t_L g2256 ( 
.A(n_1776),
.Y(n_2256)
);

AOI22xp5_ASAP7_75t_L g2257 ( 
.A1(n_1824),
.A2(n_1277),
.B1(n_1590),
.B2(n_1581),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2072),
.B(n_1737),
.Y(n_2258)
);

INVx3_ASAP7_75t_L g2259 ( 
.A(n_2002),
.Y(n_2259)
);

INVx3_ASAP7_75t_L g2260 ( 
.A(n_2012),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_1739),
.B(n_1590),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2012),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2012),
.Y(n_2263)
);

OA21x2_ASAP7_75t_L g2264 ( 
.A1(n_1909),
.A2(n_1408),
.B(n_1406),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2012),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2039),
.Y(n_2266)
);

OAI22xp5_ASAP7_75t_SL g2267 ( 
.A1(n_2080),
.A2(n_1416),
.B1(n_1473),
.B2(n_1535),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_1791),
.B(n_1410),
.Y(n_2268)
);

INVx3_ASAP7_75t_L g2269 ( 
.A(n_2039),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2039),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2039),
.Y(n_2271)
);

INVx6_ASAP7_75t_L g2272 ( 
.A(n_1805),
.Y(n_2272)
);

NOR2xp33_ASAP7_75t_L g2273 ( 
.A(n_1811),
.B(n_1671),
.Y(n_2273)
);

INVx3_ASAP7_75t_L g2274 ( 
.A(n_2043),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2043),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2043),
.Y(n_2276)
);

OAI22xp5_ASAP7_75t_SL g2277 ( 
.A1(n_2080),
.A2(n_1538),
.B1(n_1575),
.B2(n_1550),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_1909),
.Y(n_2278)
);

INVxp67_ASAP7_75t_L g2279 ( 
.A(n_1995),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_1994),
.B(n_2000),
.Y(n_2280)
);

BUFx6f_ASAP7_75t_L g2281 ( 
.A(n_1902),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_2005),
.B(n_1411),
.Y(n_2282)
);

INVxp67_ASAP7_75t_L g2283 ( 
.A(n_2007),
.Y(n_2283)
);

OAI21x1_ASAP7_75t_L g2284 ( 
.A1(n_1939),
.A2(n_1414),
.B(n_1412),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_1916),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_1916),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_2009),
.B(n_1418),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2043),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_SL g2289 ( 
.A(n_1976),
.B(n_1226),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2048),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2048),
.Y(n_2291)
);

INVx3_ASAP7_75t_L g2292 ( 
.A(n_1808),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_1818),
.B(n_1419),
.Y(n_2293)
);

HB1xp67_ASAP7_75t_L g2294 ( 
.A(n_1746),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2048),
.Y(n_2295)
);

INVx3_ASAP7_75t_L g2296 ( 
.A(n_1849),
.Y(n_2296)
);

BUFx6f_ASAP7_75t_L g2297 ( 
.A(n_1902),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2048),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_1929),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_1749),
.B(n_1422),
.Y(n_2300)
);

BUFx6f_ASAP7_75t_L g2301 ( 
.A(n_1907),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2060),
.Y(n_2302)
);

BUFx6f_ASAP7_75t_L g2303 ( 
.A(n_1907),
.Y(n_2303)
);

BUFx6f_ASAP7_75t_L g2304 ( 
.A(n_1907),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_1929),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_1827),
.B(n_1423),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2060),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_1827),
.B(n_1850),
.Y(n_2308)
);

HB1xp67_ASAP7_75t_L g2309 ( 
.A(n_1768),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_1849),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2060),
.Y(n_2311)
);

AND2x4_ASAP7_75t_L g2312 ( 
.A(n_1942),
.B(n_1688),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_1859),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2060),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2061),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_1893),
.B(n_1424),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_1859),
.Y(n_2317)
);

BUFx8_ASAP7_75t_L g2318 ( 
.A(n_1782),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2061),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2061),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_1893),
.B(n_1925),
.Y(n_2321)
);

HB1xp67_ASAP7_75t_L g2322 ( 
.A(n_1768),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2061),
.Y(n_2323)
);

AND2x4_ASAP7_75t_L g2324 ( 
.A(n_1942),
.B(n_1699),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2066),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2066),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2066),
.Y(n_2327)
);

OAI21x1_ASAP7_75t_L g2328 ( 
.A1(n_1952),
.A2(n_1426),
.B(n_1425),
.Y(n_2328)
);

NOR2xp33_ASAP7_75t_L g2329 ( 
.A(n_1727),
.B(n_1705),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2066),
.Y(n_2330)
);

INVx3_ASAP7_75t_L g2331 ( 
.A(n_2074),
.Y(n_2331)
);

OAI21x1_ASAP7_75t_L g2332 ( 
.A1(n_1764),
.A2(n_1429),
.B(n_1428),
.Y(n_2332)
);

BUFx6f_ASAP7_75t_L g2333 ( 
.A(n_1907),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_1860),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2074),
.Y(n_2335)
);

INVx4_ASAP7_75t_L g2336 ( 
.A(n_2008),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_2034),
.B(n_1430),
.Y(n_2337)
);

INVxp67_ASAP7_75t_L g2338 ( 
.A(n_2021),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2074),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2074),
.Y(n_2340)
);

CKINVDCx16_ASAP7_75t_R g2341 ( 
.A(n_1787),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_2044),
.B(n_1432),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2075),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2075),
.Y(n_2344)
);

BUFx2_ASAP7_75t_L g2345 ( 
.A(n_2076),
.Y(n_2345)
);

BUFx6f_ASAP7_75t_L g2346 ( 
.A(n_1915),
.Y(n_2346)
);

AND3x2_ASAP7_75t_L g2347 ( 
.A(n_1920),
.B(n_885),
.C(n_833),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2075),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_1925),
.B(n_1433),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_1860),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2075),
.Y(n_2351)
);

BUFx6f_ASAP7_75t_L g2352 ( 
.A(n_1915),
.Y(n_2352)
);

INVx4_ASAP7_75t_L g2353 ( 
.A(n_2008),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_1961),
.Y(n_2354)
);

BUFx6f_ASAP7_75t_L g2355 ( 
.A(n_1915),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_1915),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_1961),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_1974),
.Y(n_2358)
);

AND2x6_ASAP7_75t_L g2359 ( 
.A(n_1720),
.B(n_1165),
.Y(n_2359)
);

BUFx12f_ASAP7_75t_L g2360 ( 
.A(n_1782),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_1938),
.B(n_1435),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_1938),
.B(n_1436),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_1974),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_1986),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_1986),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_1968),
.B(n_1438),
.Y(n_2366)
);

CKINVDCx5p33_ASAP7_75t_R g2367 ( 
.A(n_1967),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_1923),
.B(n_1439),
.Y(n_2368)
);

NOR2xp33_ASAP7_75t_L g2369 ( 
.A(n_1740),
.B(n_1682),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_1919),
.Y(n_2370)
);

OAI21x1_ASAP7_75t_L g2371 ( 
.A1(n_1774),
.A2(n_1443),
.B(n_1440),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_1858),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_1876),
.Y(n_2373)
);

BUFx2_ASAP7_75t_L g2374 ( 
.A(n_2076),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_1919),
.Y(n_2375)
);

BUFx6f_ASAP7_75t_L g2376 ( 
.A(n_1919),
.Y(n_2376)
);

INVx3_ASAP7_75t_L g2377 ( 
.A(n_1802),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_1879),
.Y(n_2378)
);

BUFx6f_ASAP7_75t_L g2379 ( 
.A(n_1919),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_1882),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_1968),
.B(n_1445),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_1928),
.Y(n_2382)
);

AND2x4_ASAP7_75t_L g2383 ( 
.A(n_2071),
.B(n_1703),
.Y(n_2383)
);

BUFx6f_ASAP7_75t_L g2384 ( 
.A(n_1928),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_1894),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_1928),
.Y(n_2386)
);

HB1xp67_ASAP7_75t_L g2387 ( 
.A(n_1807),
.Y(n_2387)
);

HB1xp67_ASAP7_75t_L g2388 ( 
.A(n_1807),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_1928),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_1912),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_1932),
.Y(n_2391)
);

HB1xp67_ASAP7_75t_L g2392 ( 
.A(n_1819),
.Y(n_2392)
);

AND2x4_ASAP7_75t_L g2393 ( 
.A(n_2071),
.B(n_1706),
.Y(n_2393)
);

BUFx6f_ASAP7_75t_L g2394 ( 
.A(n_1932),
.Y(n_2394)
);

INVx1_ASAP7_75t_SL g2395 ( 
.A(n_1899),
.Y(n_2395)
);

CKINVDCx5p33_ASAP7_75t_R g2396 ( 
.A(n_1967),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_1921),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_1955),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_1969),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_1754),
.B(n_1450),
.Y(n_2400)
);

NOR2xp33_ASAP7_75t_L g2401 ( 
.A(n_1760),
.B(n_1658),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_1972),
.Y(n_2402)
);

AOI22xp5_ASAP7_75t_L g2403 ( 
.A1(n_1824),
.A2(n_905),
.B1(n_1003),
.B2(n_799),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_1983),
.B(n_1451),
.Y(n_2404)
);

AOI22xp5_ASAP7_75t_L g2405 ( 
.A1(n_1983),
.A2(n_1111),
.B1(n_1124),
.B2(n_1062),
.Y(n_2405)
);

CKINVDCx8_ASAP7_75t_R g2406 ( 
.A(n_1810),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_1987),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_1997),
.Y(n_2408)
);

BUFx6f_ASAP7_75t_L g2409 ( 
.A(n_1932),
.Y(n_2409)
);

BUFx6f_ASAP7_75t_L g2410 ( 
.A(n_1932),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_1983),
.B(n_1452),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_1998),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_1715),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2047),
.Y(n_2414)
);

AND2x2_ASAP7_75t_L g2415 ( 
.A(n_1923),
.B(n_1455),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_1983),
.B(n_1814),
.Y(n_2416)
);

AOI22xp5_ASAP7_75t_L g2417 ( 
.A1(n_1731),
.A2(n_1149),
.B1(n_1214),
.B2(n_1155),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_1715),
.Y(n_2418)
);

HB1xp67_ASAP7_75t_L g2419 ( 
.A(n_1819),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_1715),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_1715),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2052),
.B(n_1456),
.Y(n_2422)
);

AND2x6_ASAP7_75t_L g2423 ( 
.A(n_1757),
.B(n_1165),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_1717),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2049),
.Y(n_2425)
);

BUFx6f_ASAP7_75t_L g2426 ( 
.A(n_1913),
.Y(n_2426)
);

AND2x2_ASAP7_75t_L g2427 ( 
.A(n_2067),
.B(n_1457),
.Y(n_2427)
);

AND2x2_ASAP7_75t_L g2428 ( 
.A(n_2068),
.B(n_1458),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2054),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_1999),
.Y(n_2430)
);

BUFx6f_ASAP7_75t_L g2431 ( 
.A(n_1717),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_1999),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2035),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2035),
.Y(n_2434)
);

BUFx6f_ASAP7_75t_L g2435 ( 
.A(n_1717),
.Y(n_2435)
);

INVxp67_ASAP7_75t_L g2436 ( 
.A(n_1744),
.Y(n_2436)
);

NAND2xp33_ASAP7_75t_L g2437 ( 
.A(n_1863),
.B(n_1226),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_1717),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2051),
.Y(n_2439)
);

CKINVDCx20_ASAP7_75t_R g2440 ( 
.A(n_1713),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2051),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2056),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_1735),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2056),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_1735),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2069),
.Y(n_2446)
);

AND2x2_ASAP7_75t_L g2447 ( 
.A(n_1790),
.B(n_1801),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_1816),
.B(n_1460),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2069),
.Y(n_2449)
);

BUFx6f_ASAP7_75t_L g2450 ( 
.A(n_1735),
.Y(n_2450)
);

AND2x6_ASAP7_75t_L g2451 ( 
.A(n_1731),
.B(n_1188),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_1735),
.Y(n_2452)
);

INVx1_ASAP7_75t_SL g2453 ( 
.A(n_1905),
.Y(n_2453)
);

CKINVDCx20_ASAP7_75t_R g2454 ( 
.A(n_1713),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_1853),
.Y(n_2455)
);

AND2x4_ASAP7_75t_L g2456 ( 
.A(n_1748),
.B(n_1665),
.Y(n_2456)
);

BUFx6f_ASAP7_75t_L g2457 ( 
.A(n_1759),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_1853),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_1759),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_1834),
.B(n_1463),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_1857),
.Y(n_2461)
);

AND2x4_ASAP7_75t_L g2462 ( 
.A(n_1748),
.B(n_1666),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_1759),
.Y(n_2463)
);

NOR2xp33_ASAP7_75t_L g2464 ( 
.A(n_1839),
.B(n_1667),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_L g2465 ( 
.A(n_1842),
.B(n_1464),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_1759),
.Y(n_2466)
);

CKINVDCx11_ASAP7_75t_R g2467 ( 
.A(n_1981),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_1857),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_1914),
.Y(n_2469)
);

OA21x2_ASAP7_75t_L g2470 ( 
.A1(n_2001),
.A2(n_1469),
.B(n_1465),
.Y(n_2470)
);

BUFx6f_ASAP7_75t_L g2471 ( 
.A(n_1763),
.Y(n_2471)
);

INVx3_ASAP7_75t_L g2472 ( 
.A(n_1802),
.Y(n_2472)
);

OR2x2_ASAP7_75t_L g2473 ( 
.A(n_1897),
.B(n_1375),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_1914),
.Y(n_2474)
);

BUFx6f_ASAP7_75t_L g2475 ( 
.A(n_1763),
.Y(n_2475)
);

BUFx6f_ASAP7_75t_L g2476 ( 
.A(n_1763),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_1948),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_1948),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_1763),
.Y(n_2479)
);

AND2x2_ASAP7_75t_L g2480 ( 
.A(n_1934),
.B(n_1470),
.Y(n_2480)
);

BUFx3_ASAP7_75t_L g2481 ( 
.A(n_1868),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_1950),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_1950),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_1770),
.Y(n_2484)
);

INVx3_ASAP7_75t_L g2485 ( 
.A(n_1822),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_1837),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2070),
.Y(n_2487)
);

BUFx8_ASAP7_75t_L g2488 ( 
.A(n_1936),
.Y(n_2488)
);

OA21x2_ASAP7_75t_L g2489 ( 
.A1(n_2001),
.A2(n_1475),
.B(n_1471),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2078),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2078),
.Y(n_2491)
);

AND2x4_ASAP7_75t_L g2492 ( 
.A(n_1721),
.B(n_1694),
.Y(n_2492)
);

BUFx6f_ASAP7_75t_L g2493 ( 
.A(n_1770),
.Y(n_2493)
);

HB1xp67_ASAP7_75t_L g2494 ( 
.A(n_1829),
.Y(n_2494)
);

NAND2xp33_ASAP7_75t_L g2495 ( 
.A(n_1877),
.B(n_1226),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_1770),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2081),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2081),
.Y(n_2498)
);

AND2x2_ASAP7_75t_L g2499 ( 
.A(n_1934),
.B(n_1476),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_1751),
.Y(n_2500)
);

OAI21x1_ASAP7_75t_L g2501 ( 
.A1(n_1781),
.A2(n_1478),
.B(n_1477),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2073),
.Y(n_2502)
);

AND2x2_ASAP7_75t_L g2503 ( 
.A(n_2280),
.B(n_2023),
.Y(n_2503)
);

NOR2xp33_ASAP7_75t_L g2504 ( 
.A(n_2207),
.B(n_2023),
.Y(n_2504)
);

NAND3xp33_ASAP7_75t_L g2505 ( 
.A(n_2175),
.B(n_2093),
.C(n_2195),
.Y(n_2505)
);

INVx4_ASAP7_75t_L g2506 ( 
.A(n_2147),
.Y(n_2506)
);

AOI22xp33_ASAP7_75t_L g2507 ( 
.A1(n_2383),
.A2(n_2080),
.B1(n_2020),
.B2(n_1829),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2159),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_2159),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2107),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_SL g2511 ( 
.A(n_2195),
.B(n_1881),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_2198),
.B(n_2063),
.Y(n_2512)
);

BUFx6f_ASAP7_75t_L g2513 ( 
.A(n_2101),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2372),
.Y(n_2514)
);

INVx2_ASAP7_75t_SL g2515 ( 
.A(n_2422),
.Y(n_2515)
);

AOI22xp33_ASAP7_75t_L g2516 ( 
.A1(n_2383),
.A2(n_2020),
.B1(n_1908),
.B2(n_1904),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_2223),
.B(n_1976),
.Y(n_2517)
);

AND2x2_ASAP7_75t_L g2518 ( 
.A(n_2216),
.B(n_2063),
.Y(n_2518)
);

INVx2_ASAP7_75t_L g2519 ( 
.A(n_2159),
.Y(n_2519)
);

INVxp33_ASAP7_75t_SL g2520 ( 
.A(n_2084),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2373),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2087),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_2087),
.Y(n_2523)
);

AO21x2_ASAP7_75t_L g2524 ( 
.A1(n_2332),
.A2(n_1793),
.B(n_1786),
.Y(n_2524)
);

INVx2_ASAP7_75t_L g2525 ( 
.A(n_2089),
.Y(n_2525)
);

INVx2_ASAP7_75t_SL g2526 ( 
.A(n_2427),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2378),
.Y(n_2527)
);

INVx3_ASAP7_75t_L g2528 ( 
.A(n_2107),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2107),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2264),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2089),
.Y(n_2531)
);

NAND2xp33_ASAP7_75t_L g2532 ( 
.A(n_2248),
.B(n_1941),
.Y(n_2532)
);

INVx2_ASAP7_75t_SL g2533 ( 
.A(n_2428),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2380),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2385),
.Y(n_2535)
);

HB1xp67_ASAP7_75t_L g2536 ( 
.A(n_2395),
.Y(n_2536)
);

BUFx10_ASAP7_75t_L g2537 ( 
.A(n_2084),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2390),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_2096),
.Y(n_2539)
);

NOR2xp33_ASAP7_75t_L g2540 ( 
.A(n_2212),
.B(n_1726),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_SL g2541 ( 
.A(n_2214),
.B(n_1881),
.Y(n_2541)
);

NOR2xp33_ASAP7_75t_L g2542 ( 
.A(n_2236),
.B(n_1726),
.Y(n_2542)
);

INVx2_ASAP7_75t_SL g2543 ( 
.A(n_2448),
.Y(n_2543)
);

INVxp67_ASAP7_75t_SL g2544 ( 
.A(n_2097),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_L g2545 ( 
.A(n_2401),
.B(n_1989),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2096),
.Y(n_2546)
);

BUFx6f_ASAP7_75t_L g2547 ( 
.A(n_2101),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2106),
.Y(n_2548)
);

NOR2xp33_ASAP7_75t_L g2549 ( 
.A(n_2093),
.B(n_1989),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2106),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2108),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_SL g2552 ( 
.A(n_2141),
.B(n_1957),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2108),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_2115),
.Y(n_2554)
);

CKINVDCx20_ASAP7_75t_R g2555 ( 
.A(n_2341),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_SL g2556 ( 
.A(n_2141),
.B(n_1957),
.Y(n_2556)
);

INVx8_ASAP7_75t_L g2557 ( 
.A(n_2230),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_2115),
.Y(n_2558)
);

INVx2_ASAP7_75t_L g2559 ( 
.A(n_2117),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_SL g2560 ( 
.A(n_2233),
.B(n_1970),
.Y(n_2560)
);

INVx2_ASAP7_75t_L g2561 ( 
.A(n_2117),
.Y(n_2561)
);

NAND3xp33_ASAP7_75t_L g2562 ( 
.A(n_2220),
.B(n_2247),
.C(n_2206),
.Y(n_2562)
);

INVx8_ASAP7_75t_L g2563 ( 
.A(n_2230),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2397),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2398),
.Y(n_2565)
);

CKINVDCx5p33_ASAP7_75t_R g2566 ( 
.A(n_2125),
.Y(n_2566)
);

NOR2xp33_ASAP7_75t_L g2567 ( 
.A(n_2251),
.B(n_2006),
.Y(n_2567)
);

INVx5_ASAP7_75t_L g2568 ( 
.A(n_2090),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_SL g2569 ( 
.A(n_2105),
.B(n_1970),
.Y(n_2569)
);

OAI22xp33_ASAP7_75t_L g2570 ( 
.A1(n_2257),
.A2(n_1832),
.B1(n_1991),
.B2(n_1981),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2119),
.Y(n_2571)
);

INVx2_ASAP7_75t_L g2572 ( 
.A(n_2119),
.Y(n_2572)
);

BUFx10_ASAP7_75t_L g2573 ( 
.A(n_2125),
.Y(n_2573)
);

INVx2_ASAP7_75t_L g2574 ( 
.A(n_2156),
.Y(n_2574)
);

AND2x2_ASAP7_75t_L g2575 ( 
.A(n_2240),
.B(n_1935),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_2156),
.Y(n_2576)
);

AO21x2_ASAP7_75t_L g2577 ( 
.A1(n_2332),
.A2(n_2501),
.B(n_2371),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_2158),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_L g2579 ( 
.A(n_2401),
.B(n_1752),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2264),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_SL g2581 ( 
.A(n_2085),
.B(n_2027),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_2158),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_2161),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2264),
.Y(n_2584)
);

INVx2_ASAP7_75t_SL g2585 ( 
.A(n_2176),
.Y(n_2585)
);

INVx2_ASAP7_75t_L g2586 ( 
.A(n_2161),
.Y(n_2586)
);

INVx8_ASAP7_75t_L g2587 ( 
.A(n_2230),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2163),
.Y(n_2588)
);

INVx2_ASAP7_75t_SL g2589 ( 
.A(n_2176),
.Y(n_2589)
);

CKINVDCx5p33_ASAP7_75t_R g2590 ( 
.A(n_2367),
.Y(n_2590)
);

OAI22xp33_ASAP7_75t_L g2591 ( 
.A1(n_2405),
.A2(n_2019),
.B1(n_2058),
.B2(n_1991),
.Y(n_2591)
);

HB1xp67_ASAP7_75t_L g2592 ( 
.A(n_2453),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_2163),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2165),
.Y(n_2594)
);

INVx2_ASAP7_75t_L g2595 ( 
.A(n_2165),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2329),
.B(n_2041),
.Y(n_2596)
);

INVx2_ASAP7_75t_L g2597 ( 
.A(n_2170),
.Y(n_2597)
);

BUFx2_ASAP7_75t_L g2598 ( 
.A(n_2083),
.Y(n_2598)
);

NAND2xp33_ASAP7_75t_L g2599 ( 
.A(n_2451),
.B(n_1935),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2329),
.B(n_2013),
.Y(n_2600)
);

AOI22xp33_ASAP7_75t_L g2601 ( 
.A1(n_2383),
.A2(n_1908),
.B1(n_1904),
.B2(n_1940),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_SL g2602 ( 
.A(n_2110),
.B(n_1958),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_2170),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2172),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2172),
.Y(n_2605)
);

INVx2_ASAP7_75t_SL g2606 ( 
.A(n_2176),
.Y(n_2606)
);

INVx8_ASAP7_75t_L g2607 ( 
.A(n_2230),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2173),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2369),
.B(n_2013),
.Y(n_2609)
);

NAND3xp33_ASAP7_75t_L g2610 ( 
.A(n_2220),
.B(n_2247),
.C(n_2206),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_2173),
.Y(n_2611)
);

OR2x2_ASAP7_75t_L g2612 ( 
.A(n_2208),
.B(n_1930),
.Y(n_2612)
);

NAND3xp33_ASAP7_75t_L g2613 ( 
.A(n_2369),
.B(n_1975),
.C(n_1958),
.Y(n_2613)
);

CKINVDCx20_ASAP7_75t_R g2614 ( 
.A(n_2440),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2399),
.Y(n_2615)
);

BUFx3_ASAP7_75t_L g2616 ( 
.A(n_2241),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2193),
.Y(n_2617)
);

AND2x2_ASAP7_75t_L g2618 ( 
.A(n_2368),
.B(n_1975),
.Y(n_2618)
);

INVx2_ASAP7_75t_L g2619 ( 
.A(n_2193),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2402),
.Y(n_2620)
);

INVx2_ASAP7_75t_L g2621 ( 
.A(n_2209),
.Y(n_2621)
);

NAND2xp33_ASAP7_75t_L g2622 ( 
.A(n_2451),
.B(n_1851),
.Y(n_2622)
);

BUFx6f_ASAP7_75t_L g2623 ( 
.A(n_2101),
.Y(n_2623)
);

NOR2xp33_ASAP7_75t_L g2624 ( 
.A(n_2279),
.B(n_1870),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2407),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2209),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2408),
.Y(n_2627)
);

INVx2_ASAP7_75t_L g2628 ( 
.A(n_2210),
.Y(n_2628)
);

INVx3_ASAP7_75t_L g2629 ( 
.A(n_2180),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2210),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_SL g2631 ( 
.A(n_2122),
.B(n_1944),
.Y(n_2631)
);

INVx2_ASAP7_75t_L g2632 ( 
.A(n_2226),
.Y(n_2632)
);

INVx2_ASAP7_75t_L g2633 ( 
.A(n_2226),
.Y(n_2633)
);

INVx2_ASAP7_75t_L g2634 ( 
.A(n_2229),
.Y(n_2634)
);

INVx3_ASAP7_75t_L g2635 ( 
.A(n_2180),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2412),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2229),
.Y(n_2637)
);

NOR2xp33_ASAP7_75t_L g2638 ( 
.A(n_2283),
.B(n_1944),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2414),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2425),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2429),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2082),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2086),
.Y(n_2643)
);

INVx1_ASAP7_75t_SL g2644 ( 
.A(n_2225),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2500),
.B(n_2014),
.Y(n_2645)
);

BUFx6f_ASAP7_75t_L g2646 ( 
.A(n_2101),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2091),
.Y(n_2647)
);

AND2x2_ASAP7_75t_L g2648 ( 
.A(n_2415),
.B(n_1940),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2094),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2095),
.Y(n_2650)
);

AOI22xp33_ASAP7_75t_L g2651 ( 
.A1(n_2393),
.A2(n_2010),
.B1(n_2004),
.B2(n_1798),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_SL g2652 ( 
.A(n_2132),
.B(n_1944),
.Y(n_2652)
);

INVx2_ASAP7_75t_L g2653 ( 
.A(n_2231),
.Y(n_2653)
);

AOI22xp5_ASAP7_75t_L g2654 ( 
.A1(n_2451),
.A2(n_1943),
.B1(n_2014),
.B2(n_1891),
.Y(n_2654)
);

BUFx6f_ASAP7_75t_L g2655 ( 
.A(n_2103),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_SL g2656 ( 
.A(n_2194),
.B(n_1944),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2100),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2104),
.Y(n_2658)
);

AOI21x1_ASAP7_75t_L g2659 ( 
.A1(n_2416),
.A2(n_1864),
.B(n_1856),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2109),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2113),
.Y(n_2661)
);

CKINVDCx11_ASAP7_75t_R g2662 ( 
.A(n_2440),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2116),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2464),
.B(n_2017),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2118),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2120),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2088),
.Y(n_2667)
);

INVx2_ASAP7_75t_SL g2668 ( 
.A(n_2097),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2088),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_SL g2670 ( 
.A(n_2261),
.B(n_1947),
.Y(n_2670)
);

INVx2_ASAP7_75t_L g2671 ( 
.A(n_2231),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_SL g2672 ( 
.A(n_2232),
.B(n_1947),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_2235),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_SL g2674 ( 
.A(n_2232),
.B(n_1947),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_SL g2675 ( 
.A(n_2174),
.B(n_1947),
.Y(n_2675)
);

AND2x2_ASAP7_75t_L g2676 ( 
.A(n_2337),
.B(n_2004),
.Y(n_2676)
);

INVx2_ASAP7_75t_SL g2677 ( 
.A(n_2127),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2235),
.Y(n_2678)
);

AO21x2_ASAP7_75t_L g2679 ( 
.A1(n_2371),
.A2(n_1869),
.B(n_1866),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_SL g2680 ( 
.A(n_2174),
.B(n_1951),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2242),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_L g2682 ( 
.A(n_2464),
.B(n_2038),
.Y(n_2682)
);

INVx3_ASAP7_75t_L g2683 ( 
.A(n_2180),
.Y(n_2683)
);

NAND2xp33_ASAP7_75t_L g2684 ( 
.A(n_2451),
.B(n_1878),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2242),
.Y(n_2685)
);

CKINVDCx6p67_ASAP7_75t_R g2686 ( 
.A(n_2360),
.Y(n_2686)
);

INVx2_ASAP7_75t_L g2687 ( 
.A(n_2244),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_SL g2688 ( 
.A(n_2492),
.B(n_1951),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2088),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2244),
.Y(n_2690)
);

BUFx8_ASAP7_75t_SL g2691 ( 
.A(n_2454),
.Y(n_2691)
);

INVx2_ASAP7_75t_L g2692 ( 
.A(n_2245),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2102),
.Y(n_2693)
);

INVx2_ASAP7_75t_L g2694 ( 
.A(n_2245),
.Y(n_2694)
);

INVx2_ASAP7_75t_L g2695 ( 
.A(n_2253),
.Y(n_2695)
);

INVx2_ASAP7_75t_L g2696 ( 
.A(n_2253),
.Y(n_2696)
);

INVx2_ASAP7_75t_L g2697 ( 
.A(n_2255),
.Y(n_2697)
);

INVx3_ASAP7_75t_L g2698 ( 
.A(n_2196),
.Y(n_2698)
);

AND2x2_ASAP7_75t_L g2699 ( 
.A(n_2342),
.B(n_2010),
.Y(n_2699)
);

INVx2_ASAP7_75t_L g2700 ( 
.A(n_2255),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_2278),
.Y(n_2701)
);

OAI22xp33_ASAP7_75t_L g2702 ( 
.A1(n_2403),
.A2(n_2309),
.B1(n_2387),
.B2(n_2322),
.Y(n_2702)
);

INVx2_ASAP7_75t_L g2703 ( 
.A(n_2278),
.Y(n_2703)
);

INVxp67_ASAP7_75t_L g2704 ( 
.A(n_2447),
.Y(n_2704)
);

NOR2xp33_ASAP7_75t_L g2705 ( 
.A(n_2436),
.B(n_2123),
.Y(n_2705)
);

OR2x6_ASAP7_75t_L g2706 ( 
.A(n_2202),
.B(n_1936),
.Y(n_2706)
);

INVx2_ASAP7_75t_L g2707 ( 
.A(n_2285),
.Y(n_2707)
);

NAND3xp33_ASAP7_75t_L g2708 ( 
.A(n_2092),
.B(n_1996),
.C(n_1951),
.Y(n_2708)
);

NOR2xp33_ASAP7_75t_L g2709 ( 
.A(n_2123),
.B(n_1951),
.Y(n_2709)
);

INVx2_ASAP7_75t_L g2710 ( 
.A(n_2285),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2286),
.Y(n_2711)
);

NOR2xp33_ASAP7_75t_L g2712 ( 
.A(n_2131),
.B(n_1996),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2258),
.B(n_1891),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2286),
.Y(n_2714)
);

INVx3_ASAP7_75t_L g2715 ( 
.A(n_2196),
.Y(n_2715)
);

INVx2_ASAP7_75t_L g2716 ( 
.A(n_2299),
.Y(n_2716)
);

AOI22xp33_ASAP7_75t_L g2717 ( 
.A1(n_2393),
.A2(n_1798),
.B1(n_1756),
.B2(n_2045),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_L g2718 ( 
.A(n_2492),
.B(n_2400),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2299),
.Y(n_2719)
);

OR2x2_ASAP7_75t_L g2720 ( 
.A(n_2177),
.B(n_2079),
.Y(n_2720)
);

INVx5_ASAP7_75t_L g2721 ( 
.A(n_2090),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2102),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2102),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_SL g2724 ( 
.A(n_2492),
.B(n_1996),
.Y(n_2724)
);

INVx5_ASAP7_75t_L g2725 ( 
.A(n_2090),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_SL g2726 ( 
.A(n_2456),
.B(n_1996),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2305),
.Y(n_2727)
);

AND2x2_ASAP7_75t_L g2728 ( 
.A(n_2252),
.B(n_2018),
.Y(n_2728)
);

NAND3xp33_ASAP7_75t_L g2729 ( 
.A(n_2092),
.B(n_2028),
.C(n_2026),
.Y(n_2729)
);

INVx2_ASAP7_75t_L g2730 ( 
.A(n_2305),
.Y(n_2730)
);

BUFx6f_ASAP7_75t_L g2731 ( 
.A(n_2103),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2200),
.Y(n_2732)
);

INVx2_ASAP7_75t_L g2733 ( 
.A(n_2200),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2111),
.Y(n_2734)
);

INVx2_ASAP7_75t_L g2735 ( 
.A(n_2284),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2393),
.B(n_1844),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2111),
.Y(n_2737)
);

INVx2_ASAP7_75t_L g2738 ( 
.A(n_2284),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2308),
.B(n_2026),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2111),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2160),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_L g2742 ( 
.A(n_2321),
.B(n_2026),
.Y(n_2742)
);

INVx2_ASAP7_75t_SL g2743 ( 
.A(n_2127),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2328),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_SL g2745 ( 
.A(n_2456),
.B(n_2026),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2328),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2160),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_SL g2748 ( 
.A(n_2456),
.B(n_2028),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2460),
.B(n_2465),
.Y(n_2749)
);

AND2x2_ASAP7_75t_L g2750 ( 
.A(n_2282),
.B(n_2018),
.Y(n_2750)
);

BUFx3_ASAP7_75t_L g2751 ( 
.A(n_2241),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2160),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2310),
.Y(n_2753)
);

INVx2_ASAP7_75t_L g2754 ( 
.A(n_2310),
.Y(n_2754)
);

INVx2_ASAP7_75t_L g2755 ( 
.A(n_2313),
.Y(n_2755)
);

INVx5_ASAP7_75t_L g2756 ( 
.A(n_2152),
.Y(n_2756)
);

HB1xp67_ASAP7_75t_L g2757 ( 
.A(n_2201),
.Y(n_2757)
);

INVxp33_ASAP7_75t_L g2758 ( 
.A(n_2143),
.Y(n_2758)
);

INVx2_ASAP7_75t_L g2759 ( 
.A(n_2313),
.Y(n_2759)
);

NAND2xp33_ASAP7_75t_R g2760 ( 
.A(n_2367),
.B(n_2396),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2487),
.B(n_2190),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2317),
.Y(n_2762)
);

NOR2xp33_ASAP7_75t_L g2763 ( 
.A(n_2131),
.B(n_1799),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_2317),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2334),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2334),
.Y(n_2766)
);

AND2x2_ASAP7_75t_L g2767 ( 
.A(n_2287),
.B(n_2022),
.Y(n_2767)
);

INVx2_ASAP7_75t_L g2768 ( 
.A(n_2350),
.Y(n_2768)
);

INVx2_ASAP7_75t_SL g2769 ( 
.A(n_2213),
.Y(n_2769)
);

BUFx6f_ASAP7_75t_L g2770 ( 
.A(n_2103),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2350),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_L g2772 ( 
.A(n_2190),
.B(n_2028),
.Y(n_2772)
);

INVx2_ASAP7_75t_L g2773 ( 
.A(n_2196),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2470),
.Y(n_2774)
);

BUFx10_ASAP7_75t_L g2775 ( 
.A(n_2396),
.Y(n_2775)
);

HB1xp67_ASAP7_75t_L g2776 ( 
.A(n_2143),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2205),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2205),
.Y(n_2778)
);

AO21x2_ASAP7_75t_L g2779 ( 
.A1(n_2501),
.A2(n_2186),
.B(n_2404),
.Y(n_2779)
);

HB1xp67_ASAP7_75t_L g2780 ( 
.A(n_2168),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_2205),
.Y(n_2781)
);

INVx2_ASAP7_75t_L g2782 ( 
.A(n_2292),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_SL g2783 ( 
.A(n_2462),
.B(n_2480),
.Y(n_2783)
);

OAI22xp5_ASAP7_75t_L g2784 ( 
.A1(n_2228),
.A2(n_1039),
.B1(n_1159),
.B2(n_896),
.Y(n_2784)
);

INVx2_ASAP7_75t_L g2785 ( 
.A(n_2292),
.Y(n_2785)
);

BUFx3_ASAP7_75t_L g2786 ( 
.A(n_2241),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2470),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2190),
.B(n_2028),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_L g2789 ( 
.A(n_2300),
.B(n_2031),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2292),
.Y(n_2790)
);

INVx2_ASAP7_75t_L g2791 ( 
.A(n_2296),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_SL g2792 ( 
.A(n_2462),
.B(n_2499),
.Y(n_2792)
);

INVx2_ASAP7_75t_L g2793 ( 
.A(n_2296),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2470),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2489),
.Y(n_2795)
);

NOR2x1p5_ASAP7_75t_L g2796 ( 
.A(n_2360),
.B(n_2019),
.Y(n_2796)
);

AND2x2_ASAP7_75t_L g2797 ( 
.A(n_2309),
.B(n_2022),
.Y(n_2797)
);

AND2x2_ASAP7_75t_L g2798 ( 
.A(n_2322),
.B(n_2036),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2189),
.Y(n_2799)
);

INVx2_ASAP7_75t_L g2800 ( 
.A(n_2296),
.Y(n_2800)
);

INVx2_ASAP7_75t_L g2801 ( 
.A(n_2356),
.Y(n_2801)
);

INVx2_ASAP7_75t_L g2802 ( 
.A(n_2356),
.Y(n_2802)
);

OR2x6_ASAP7_75t_L g2803 ( 
.A(n_2202),
.B(n_1953),
.Y(n_2803)
);

INVx3_ASAP7_75t_L g2804 ( 
.A(n_2370),
.Y(n_2804)
);

INVxp33_ASAP7_75t_L g2805 ( 
.A(n_2168),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2370),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_2375),
.Y(n_2807)
);

AND2x2_ASAP7_75t_L g2808 ( 
.A(n_2387),
.B(n_2036),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2189),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2189),
.B(n_2031),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2430),
.Y(n_2811)
);

NAND2xp33_ASAP7_75t_SL g2812 ( 
.A(n_2294),
.B(n_2228),
.Y(n_2812)
);

INVx3_ASAP7_75t_L g2813 ( 
.A(n_2375),
.Y(n_2813)
);

NOR2xp33_ASAP7_75t_L g2814 ( 
.A(n_2187),
.B(n_1799),
.Y(n_2814)
);

OAI22xp5_ASAP7_75t_L g2815 ( 
.A1(n_2187),
.A2(n_1230),
.B1(n_816),
.B2(n_817),
.Y(n_2815)
);

AND2x2_ASAP7_75t_L g2816 ( 
.A(n_2388),
.B(n_2040),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2382),
.Y(n_2817)
);

INVx2_ASAP7_75t_L g2818 ( 
.A(n_2382),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_SL g2819 ( 
.A(n_2462),
.B(n_2031),
.Y(n_2819)
);

INVxp33_ASAP7_75t_SL g2820 ( 
.A(n_2294),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2386),
.Y(n_2821)
);

INVx2_ASAP7_75t_L g2822 ( 
.A(n_2386),
.Y(n_2822)
);

NOR2xp33_ASAP7_75t_L g2823 ( 
.A(n_2338),
.B(n_1817),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_SL g2824 ( 
.A(n_2126),
.B(n_2031),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2432),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_SL g2826 ( 
.A(n_2312),
.B(n_2037),
.Y(n_2826)
);

INVx2_ASAP7_75t_L g2827 ( 
.A(n_2389),
.Y(n_2827)
);

INVx3_ASAP7_75t_L g2828 ( 
.A(n_2389),
.Y(n_2828)
);

INVx2_ASAP7_75t_L g2829 ( 
.A(n_2391),
.Y(n_2829)
);

INVx3_ASAP7_75t_L g2830 ( 
.A(n_2391),
.Y(n_2830)
);

AND2x2_ASAP7_75t_L g2831 ( 
.A(n_2388),
.B(n_2040),
.Y(n_2831)
);

INVx2_ASAP7_75t_L g2832 ( 
.A(n_2103),
.Y(n_2832)
);

INVx8_ASAP7_75t_L g2833 ( 
.A(n_2230),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2433),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2434),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_L g2836 ( 
.A(n_2316),
.B(n_2037),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2439),
.Y(n_2837)
);

OR2x2_ASAP7_75t_L g2838 ( 
.A(n_2177),
.B(n_2057),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2349),
.B(n_2037),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2441),
.Y(n_2840)
);

INVx2_ASAP7_75t_SL g2841 ( 
.A(n_2213),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2121),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_2121),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2442),
.Y(n_2844)
);

INVx3_ASAP7_75t_L g2845 ( 
.A(n_2121),
.Y(n_2845)
);

INVx2_ASAP7_75t_L g2846 ( 
.A(n_2121),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2444),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2166),
.Y(n_2848)
);

INVx5_ASAP7_75t_L g2849 ( 
.A(n_2152),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2446),
.Y(n_2850)
);

INVx3_ASAP7_75t_L g2851 ( 
.A(n_2166),
.Y(n_2851)
);

AOI21x1_ASAP7_75t_L g2852 ( 
.A1(n_2411),
.A2(n_1903),
.B(n_1900),
.Y(n_2852)
);

INVx4_ASAP7_75t_L g2853 ( 
.A(n_2147),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_L g2854 ( 
.A(n_2361),
.B(n_2037),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_SL g2855 ( 
.A(n_2312),
.B(n_2046),
.Y(n_2855)
);

AND2x6_ASAP7_75t_L g2856 ( 
.A(n_2486),
.B(n_2057),
.Y(n_2856)
);

INVx2_ASAP7_75t_L g2857 ( 
.A(n_2166),
.Y(n_2857)
);

INVx2_ASAP7_75t_L g2858 ( 
.A(n_2166),
.Y(n_2858)
);

INVxp33_ASAP7_75t_L g2859 ( 
.A(n_2204),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2489),
.Y(n_2860)
);

INVx2_ASAP7_75t_L g2861 ( 
.A(n_2169),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2489),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_SL g2863 ( 
.A(n_2312),
.B(n_2046),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2136),
.Y(n_2864)
);

INVx4_ASAP7_75t_L g2865 ( 
.A(n_2147),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2137),
.Y(n_2866)
);

INVx2_ASAP7_75t_SL g2867 ( 
.A(n_2217),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2362),
.B(n_2366),
.Y(n_2868)
);

INVx3_ASAP7_75t_L g2869 ( 
.A(n_2169),
.Y(n_2869)
);

INVx2_ASAP7_75t_L g2870 ( 
.A(n_2169),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2138),
.Y(n_2871)
);

INVx2_ASAP7_75t_L g2872 ( 
.A(n_2169),
.Y(n_2872)
);

BUFx10_ASAP7_75t_L g2873 ( 
.A(n_2347),
.Y(n_2873)
);

BUFx6f_ASAP7_75t_SL g2874 ( 
.A(n_2202),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2140),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2381),
.B(n_2046),
.Y(n_2876)
);

BUFx6f_ASAP7_75t_L g2877 ( 
.A(n_2203),
.Y(n_2877)
);

CKINVDCx5p33_ASAP7_75t_R g2878 ( 
.A(n_2467),
.Y(n_2878)
);

INVx2_ASAP7_75t_L g2879 ( 
.A(n_2203),
.Y(n_2879)
);

BUFx2_ASAP7_75t_L g2880 ( 
.A(n_2204),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2203),
.Y(n_2881)
);

NOR2xp33_ASAP7_75t_L g2882 ( 
.A(n_2392),
.B(n_1817),
.Y(n_2882)
);

INVx2_ASAP7_75t_L g2883 ( 
.A(n_2203),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2215),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2142),
.Y(n_2885)
);

INVx1_ASAP7_75t_SL g2886 ( 
.A(n_2114),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_SL g2887 ( 
.A(n_2324),
.B(n_2046),
.Y(n_2887)
);

NOR2x1p5_ASAP7_75t_L g2888 ( 
.A(n_2473),
.B(n_2058),
.Y(n_2888)
);

INVx2_ASAP7_75t_L g2889 ( 
.A(n_2215),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2145),
.Y(n_2890)
);

NOR2x1p5_ASAP7_75t_L g2891 ( 
.A(n_2135),
.B(n_1873),
.Y(n_2891)
);

INVx2_ASAP7_75t_L g2892 ( 
.A(n_2215),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2148),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2150),
.Y(n_2894)
);

NAND2xp33_ASAP7_75t_L g2895 ( 
.A(n_2451),
.B(n_1911),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_SL g2896 ( 
.A(n_2324),
.B(n_2059),
.Y(n_2896)
);

AOI22xp33_ASAP7_75t_L g2897 ( 
.A1(n_2392),
.A2(n_1798),
.B1(n_1756),
.B2(n_2045),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_SL g2898 ( 
.A(n_2324),
.B(n_2059),
.Y(n_2898)
);

NOR2xp33_ASAP7_75t_L g2899 ( 
.A(n_2419),
.B(n_1873),
.Y(n_2899)
);

INVx2_ASAP7_75t_L g2900 ( 
.A(n_2215),
.Y(n_2900)
);

INVx3_ASAP7_75t_L g2901 ( 
.A(n_2221),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2221),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2153),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_SL g2904 ( 
.A(n_2419),
.B(n_2059),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2155),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2221),
.Y(n_2906)
);

INVx2_ASAP7_75t_SL g2907 ( 
.A(n_2217),
.Y(n_2907)
);

INVx1_ASAP7_75t_SL g2908 ( 
.A(n_2134),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2157),
.Y(n_2909)
);

INVx2_ASAP7_75t_SL g2910 ( 
.A(n_2272),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2167),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_2221),
.Y(n_2912)
);

AOI22xp5_ASAP7_75t_L g2913 ( 
.A1(n_2359),
.A2(n_1943),
.B1(n_1798),
.B2(n_1756),
.Y(n_2913)
);

INVx2_ASAP7_75t_L g2914 ( 
.A(n_2234),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2179),
.Y(n_2915)
);

BUFx2_ASAP7_75t_L g2916 ( 
.A(n_2134),
.Y(n_2916)
);

OR2x2_ASAP7_75t_L g2917 ( 
.A(n_2494),
.B(n_2065),
.Y(n_2917)
);

OR2x2_ASAP7_75t_L g2918 ( 
.A(n_2494),
.B(n_2065),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_SL g2919 ( 
.A(n_2417),
.B(n_2059),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2181),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2182),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_SL g2922 ( 
.A(n_2098),
.B(n_2062),
.Y(n_2922)
);

INVx2_ASAP7_75t_L g2923 ( 
.A(n_2234),
.Y(n_2923)
);

CKINVDCx20_ASAP7_75t_R g2924 ( 
.A(n_2454),
.Y(n_2924)
);

NAND2xp5_ASAP7_75t_SL g2925 ( 
.A(n_2098),
.B(n_2062),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2449),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2455),
.Y(n_2927)
);

INVx3_ASAP7_75t_L g2928 ( 
.A(n_2234),
.Y(n_2928)
);

INVx2_ASAP7_75t_SL g2929 ( 
.A(n_2272),
.Y(n_2929)
);

INVx3_ASAP7_75t_L g2930 ( 
.A(n_2234),
.Y(n_2930)
);

INVxp67_ASAP7_75t_L g2931 ( 
.A(n_2139),
.Y(n_2931)
);

INVx5_ASAP7_75t_L g2932 ( 
.A(n_2152),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_2237),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_L g2934 ( 
.A(n_2306),
.B(n_2062),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_SL g2935 ( 
.A(n_2099),
.B(n_2062),
.Y(n_2935)
);

INVx8_ASAP7_75t_L g2936 ( 
.A(n_2359),
.Y(n_2936)
);

INVx2_ASAP7_75t_L g2937 ( 
.A(n_2237),
.Y(n_2937)
);

BUFx6f_ASAP7_75t_L g2938 ( 
.A(n_2513),
.Y(n_2938)
);

XNOR2x2_ASAP7_75t_L g2939 ( 
.A(n_2505),
.B(n_2144),
.Y(n_2939)
);

AND2x2_ASAP7_75t_L g2940 ( 
.A(n_2618),
.B(n_2149),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2514),
.Y(n_2941)
);

XNOR2xp5_ASAP7_75t_L g2942 ( 
.A(n_2555),
.B(n_1538),
.Y(n_2942)
);

XNOR2xp5_ASAP7_75t_L g2943 ( 
.A(n_2555),
.B(n_1550),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2521),
.Y(n_2944)
);

NOR2xp33_ASAP7_75t_L g2945 ( 
.A(n_2542),
.B(n_2162),
.Y(n_2945)
);

CKINVDCx5p33_ASAP7_75t_R g2946 ( 
.A(n_2760),
.Y(n_2946)
);

INVxp67_ASAP7_75t_SL g2947 ( 
.A(n_2510),
.Y(n_2947)
);

INVxp33_ASAP7_75t_SL g2948 ( 
.A(n_2566),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2522),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2527),
.Y(n_2950)
);

AND2x2_ASAP7_75t_L g2951 ( 
.A(n_2618),
.B(n_2164),
.Y(n_2951)
);

AND2x4_ASAP7_75t_L g2952 ( 
.A(n_2891),
.B(n_2490),
.Y(n_2952)
);

INVx2_ASAP7_75t_L g2953 ( 
.A(n_2522),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2534),
.Y(n_2954)
);

BUFx2_ASAP7_75t_L g2955 ( 
.A(n_2598),
.Y(n_2955)
);

INVxp67_ASAP7_75t_SL g2956 ( 
.A(n_2510),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2535),
.Y(n_2957)
);

NOR2x1p5_ASAP7_75t_L g2958 ( 
.A(n_2566),
.B(n_1906),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2538),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2564),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2565),
.Y(n_2961)
);

CKINVDCx5p33_ASAP7_75t_R g2962 ( 
.A(n_2691),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2615),
.Y(n_2963)
);

AOI21xp5_ASAP7_75t_L g2964 ( 
.A1(n_2749),
.A2(n_2609),
.B(n_2600),
.Y(n_2964)
);

BUFx3_ASAP7_75t_L g2965 ( 
.A(n_2598),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2620),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2625),
.Y(n_2967)
);

BUFx6f_ASAP7_75t_L g2968 ( 
.A(n_2513),
.Y(n_2968)
);

NOR2xp33_ASAP7_75t_L g2969 ( 
.A(n_2504),
.B(n_2171),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2627),
.Y(n_2970)
);

INVx1_ASAP7_75t_SL g2971 ( 
.A(n_2644),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2636),
.Y(n_2972)
);

AND2x2_ASAP7_75t_L g2973 ( 
.A(n_2512),
.B(n_2197),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_2523),
.Y(n_2974)
);

XNOR2xp5_ASAP7_75t_L g2975 ( 
.A(n_2614),
.B(n_1575),
.Y(n_2975)
);

NOR2xp33_ASAP7_75t_L g2976 ( 
.A(n_2549),
.B(n_2354),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2639),
.Y(n_2977)
);

INVxp33_ASAP7_75t_SL g2978 ( 
.A(n_2590),
.Y(n_2978)
);

XOR2xp5_ASAP7_75t_L g2979 ( 
.A(n_2590),
.B(n_1608),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2640),
.Y(n_2980)
);

AND2x2_ASAP7_75t_L g2981 ( 
.A(n_2512),
.B(n_2345),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2641),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2762),
.Y(n_2983)
);

XOR2xp5_ASAP7_75t_L g2984 ( 
.A(n_2520),
.B(n_1608),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2762),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2765),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2765),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2642),
.Y(n_2988)
);

INVx2_ASAP7_75t_L g2989 ( 
.A(n_2523),
.Y(n_2989)
);

NAND2xp33_ASAP7_75t_R g2990 ( 
.A(n_2520),
.B(n_2374),
.Y(n_2990)
);

INVxp67_ASAP7_75t_L g2991 ( 
.A(n_2536),
.Y(n_2991)
);

NOR2xp33_ASAP7_75t_L g2992 ( 
.A(n_2540),
.B(n_2357),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_L g2993 ( 
.A(n_2579),
.B(n_2359),
.Y(n_2993)
);

BUFx6f_ASAP7_75t_L g2994 ( 
.A(n_2513),
.Y(n_2994)
);

INVx2_ASAP7_75t_L g2995 ( 
.A(n_2525),
.Y(n_2995)
);

AND2x2_ASAP7_75t_L g2996 ( 
.A(n_2518),
.B(n_1980),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2643),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2647),
.Y(n_2998)
);

INVxp33_ASAP7_75t_L g2999 ( 
.A(n_2592),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2649),
.Y(n_3000)
);

INVx2_ASAP7_75t_SL g3001 ( 
.A(n_2757),
.Y(n_3001)
);

AND2x2_ASAP7_75t_L g3002 ( 
.A(n_2518),
.B(n_2406),
.Y(n_3002)
);

INVxp33_ASAP7_75t_L g3003 ( 
.A(n_2612),
.Y(n_3003)
);

NOR2xp33_ASAP7_75t_L g3004 ( 
.A(n_2562),
.B(n_2358),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2650),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2657),
.Y(n_3006)
);

INVx1_ASAP7_75t_SL g3007 ( 
.A(n_2880),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2658),
.Y(n_3008)
);

INVxp33_ASAP7_75t_L g3009 ( 
.A(n_2612),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2660),
.Y(n_3010)
);

NOR2xp33_ASAP7_75t_L g3011 ( 
.A(n_2610),
.B(n_2363),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_L g3012 ( 
.A(n_2664),
.B(n_2682),
.Y(n_3012)
);

CKINVDCx20_ASAP7_75t_R g3013 ( 
.A(n_2691),
.Y(n_3013)
);

AND2x4_ASAP7_75t_L g3014 ( 
.A(n_2515),
.B(n_2491),
.Y(n_3014)
);

BUFx2_ASAP7_75t_R g3015 ( 
.A(n_2878),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_L g3016 ( 
.A(n_2868),
.B(n_2359),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2661),
.Y(n_3017)
);

INVx2_ASAP7_75t_L g3018 ( 
.A(n_2525),
.Y(n_3018)
);

NOR2xp33_ASAP7_75t_L g3019 ( 
.A(n_2596),
.B(n_2364),
.Y(n_3019)
);

AND2x6_ASAP7_75t_L g3020 ( 
.A(n_2529),
.B(n_2498),
.Y(n_3020)
);

NOR2xp33_ASAP7_75t_L g3021 ( 
.A(n_2517),
.B(n_2365),
.Y(n_3021)
);

BUFx6f_ASAP7_75t_L g3022 ( 
.A(n_2513),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2663),
.Y(n_3023)
);

NOR2xp33_ASAP7_75t_L g3024 ( 
.A(n_2545),
.B(n_2099),
.Y(n_3024)
);

INVxp33_ASAP7_75t_L g3025 ( 
.A(n_2720),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2665),
.Y(n_3026)
);

XOR2x2_ASAP7_75t_L g3027 ( 
.A(n_2624),
.B(n_2277),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2718),
.B(n_2645),
.Y(n_3028)
);

INVxp33_ASAP7_75t_L g3029 ( 
.A(n_2720),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2666),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_2736),
.B(n_2359),
.Y(n_3031)
);

AND2x2_ASAP7_75t_L g3032 ( 
.A(n_2575),
.B(n_2406),
.Y(n_3032)
);

BUFx5_ASAP7_75t_L g3033 ( 
.A(n_2732),
.Y(n_3033)
);

XOR2xp5_ASAP7_75t_L g3034 ( 
.A(n_2614),
.B(n_1652),
.Y(n_3034)
);

AND2x4_ASAP7_75t_L g3035 ( 
.A(n_2515),
.B(n_2497),
.Y(n_3035)
);

AND2x4_ASAP7_75t_L g3036 ( 
.A(n_2526),
.B(n_2112),
.Y(n_3036)
);

AND2x4_ASAP7_75t_L g3037 ( 
.A(n_2526),
.B(n_2112),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2811),
.Y(n_3038)
);

CKINVDCx20_ASAP7_75t_R g3039 ( 
.A(n_2662),
.Y(n_3039)
);

INVx1_ASAP7_75t_SL g3040 ( 
.A(n_2880),
.Y(n_3040)
);

INVx2_ASAP7_75t_L g3041 ( 
.A(n_2531),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2825),
.Y(n_3042)
);

CKINVDCx20_ASAP7_75t_R g3043 ( 
.A(n_2662),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2834),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2835),
.Y(n_3045)
);

AND2x6_ASAP7_75t_L g3046 ( 
.A(n_2529),
.B(n_2237),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2837),
.Y(n_3047)
);

BUFx6f_ASAP7_75t_L g3048 ( 
.A(n_2513),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2713),
.B(n_2503),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2840),
.Y(n_3050)
);

NOR2xp67_ASAP7_75t_L g3051 ( 
.A(n_2613),
.B(n_1953),
.Y(n_3051)
);

XOR2xp5_ASAP7_75t_L g3052 ( 
.A(n_2924),
.B(n_1652),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2844),
.Y(n_3053)
);

NOR2xp33_ASAP7_75t_L g3054 ( 
.A(n_2503),
.B(n_2130),
.Y(n_3054)
);

INVx2_ASAP7_75t_SL g3055 ( 
.A(n_2916),
.Y(n_3055)
);

NOR2xp33_ASAP7_75t_L g3056 ( 
.A(n_2543),
.B(n_2130),
.Y(n_3056)
);

AND2x2_ASAP7_75t_L g3057 ( 
.A(n_2575),
.B(n_1655),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_L g3058 ( 
.A(n_2648),
.B(n_2273),
.Y(n_3058)
);

CKINVDCx20_ASAP7_75t_R g3059 ( 
.A(n_2924),
.Y(n_3059)
);

INVx1_ASAP7_75t_SL g3060 ( 
.A(n_2916),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2847),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2850),
.Y(n_3062)
);

CKINVDCx20_ASAP7_75t_R g3063 ( 
.A(n_2686),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2926),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2927),
.Y(n_3065)
);

NOR2xp33_ASAP7_75t_L g3066 ( 
.A(n_2543),
.B(n_2458),
.Y(n_3066)
);

AND2x2_ASAP7_75t_L g3067 ( 
.A(n_2648),
.B(n_1655),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2667),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2669),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2531),
.Y(n_3070)
);

INVxp33_ASAP7_75t_L g3071 ( 
.A(n_2776),
.Y(n_3071)
);

BUFx3_ASAP7_75t_L g3072 ( 
.A(n_2686),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2689),
.Y(n_3073)
);

CKINVDCx20_ASAP7_75t_R g3074 ( 
.A(n_2878),
.Y(n_3074)
);

XOR2xp5_ASAP7_75t_L g3075 ( 
.A(n_2820),
.B(n_1662),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2693),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2722),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2723),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_L g3079 ( 
.A(n_2629),
.B(n_2273),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2734),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2737),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2740),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2741),
.Y(n_3083)
);

AND2x2_ASAP7_75t_L g3084 ( 
.A(n_2676),
.B(n_1662),
.Y(n_3084)
);

CKINVDCx5p33_ASAP7_75t_R g3085 ( 
.A(n_2537),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2747),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2752),
.Y(n_3087)
);

CKINVDCx20_ASAP7_75t_R g3088 ( 
.A(n_2537),
.Y(n_3088)
);

INVxp33_ASAP7_75t_SL g3089 ( 
.A(n_2882),
.Y(n_3089)
);

CKINVDCx20_ASAP7_75t_R g3090 ( 
.A(n_2537),
.Y(n_3090)
);

NOR2xp67_ASAP7_75t_L g3091 ( 
.A(n_2823),
.B(n_1906),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2799),
.Y(n_3092)
);

NOR2xp33_ASAP7_75t_L g3093 ( 
.A(n_2705),
.B(n_2461),
.Y(n_3093)
);

BUFx3_ASAP7_75t_L g3094 ( 
.A(n_2573),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2809),
.Y(n_3095)
);

NOR2xp33_ASAP7_75t_L g3096 ( 
.A(n_2602),
.B(n_2468),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2594),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2594),
.Y(n_3098)
);

INVxp67_ASAP7_75t_SL g3099 ( 
.A(n_2530),
.Y(n_3099)
);

AND2x4_ASAP7_75t_L g3100 ( 
.A(n_2533),
.B(n_2706),
.Y(n_3100)
);

AND2x2_ASAP7_75t_L g3101 ( 
.A(n_2676),
.B(n_1668),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_L g3102 ( 
.A(n_2629),
.B(n_2469),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2604),
.Y(n_3103)
);

INVx2_ASAP7_75t_L g3104 ( 
.A(n_2539),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_2604),
.Y(n_3105)
);

CKINVDCx20_ASAP7_75t_R g3106 ( 
.A(n_2573),
.Y(n_3106)
);

CKINVDCx5p33_ASAP7_75t_R g3107 ( 
.A(n_2573),
.Y(n_3107)
);

AND2x6_ASAP7_75t_L g3108 ( 
.A(n_2530),
.B(n_2237),
.Y(n_3108)
);

AND2x2_ASAP7_75t_L g3109 ( 
.A(n_2699),
.B(n_1668),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2605),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2605),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_2608),
.Y(n_3112)
);

INVx2_ASAP7_75t_L g3113 ( 
.A(n_2539),
.Y(n_3113)
);

NOR2xp33_ASAP7_75t_L g3114 ( 
.A(n_2820),
.B(n_2908),
.Y(n_3114)
);

CKINVDCx20_ASAP7_75t_R g3115 ( 
.A(n_2775),
.Y(n_3115)
);

OR2x2_ASAP7_75t_L g3116 ( 
.A(n_2886),
.B(n_2267),
.Y(n_3116)
);

AND2x4_ASAP7_75t_L g3117 ( 
.A(n_2533),
.B(n_2474),
.Y(n_3117)
);

INVx2_ASAP7_75t_L g3118 ( 
.A(n_2546),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2608),
.Y(n_3119)
);

NAND2xp33_ASAP7_75t_SL g3120 ( 
.A(n_2511),
.B(n_2154),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2678),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2678),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_2711),
.Y(n_3123)
);

XOR2xp5_ASAP7_75t_L g3124 ( 
.A(n_2570),
.B(n_1605),
.Y(n_3124)
);

INVx2_ASAP7_75t_L g3125 ( 
.A(n_2546),
.Y(n_3125)
);

XOR2xp5_ASAP7_75t_L g3126 ( 
.A(n_2591),
.B(n_1605),
.Y(n_3126)
);

INVx2_ASAP7_75t_L g3127 ( 
.A(n_2548),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_2711),
.Y(n_3128)
);

NOR2xp33_ASAP7_75t_L g3129 ( 
.A(n_2931),
.B(n_2477),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_2727),
.Y(n_3130)
);

XOR2xp5_ASAP7_75t_L g3131 ( 
.A(n_2708),
.B(n_2256),
.Y(n_3131)
);

NOR2xp33_ASAP7_75t_L g3132 ( 
.A(n_2704),
.B(n_2478),
.Y(n_3132)
);

AND2x2_ASAP7_75t_L g3133 ( 
.A(n_2699),
.B(n_1830),
.Y(n_3133)
);

AND2x2_ASAP7_75t_L g3134 ( 
.A(n_2728),
.B(n_2750),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2727),
.Y(n_3135)
);

OR2x2_ASAP7_75t_L g3136 ( 
.A(n_2780),
.B(n_2268),
.Y(n_3136)
);

BUFx6f_ASAP7_75t_L g3137 ( 
.A(n_2547),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2864),
.Y(n_3138)
);

OR2x2_ASAP7_75t_L g3139 ( 
.A(n_2838),
.B(n_2293),
.Y(n_3139)
);

XOR2xp5_ASAP7_75t_L g3140 ( 
.A(n_2859),
.B(n_2256),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2864),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_2866),
.Y(n_3142)
);

NOR2xp67_ASAP7_75t_L g3143 ( 
.A(n_2763),
.B(n_1927),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2866),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2871),
.Y(n_3145)
);

INVx1_ASAP7_75t_L g3146 ( 
.A(n_2871),
.Y(n_3146)
);

INVx2_ASAP7_75t_SL g3147 ( 
.A(n_2873),
.Y(n_3147)
);

INVx2_ASAP7_75t_L g3148 ( 
.A(n_2548),
.Y(n_3148)
);

BUFx3_ASAP7_75t_L g3149 ( 
.A(n_2775),
.Y(n_3149)
);

NAND2xp5_ASAP7_75t_L g3150 ( 
.A(n_2629),
.B(n_2482),
.Y(n_3150)
);

AND2x2_ASAP7_75t_L g3151 ( 
.A(n_2728),
.B(n_1830),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_2875),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2875),
.Y(n_3153)
);

AOI21xp5_ASAP7_75t_L g3154 ( 
.A1(n_2742),
.A2(n_2186),
.B(n_2154),
.Y(n_3154)
);

AOI21xp5_ASAP7_75t_L g3155 ( 
.A1(n_2739),
.A2(n_1924),
.B(n_1917),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_2885),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2885),
.Y(n_3157)
);

NOR2xp33_ASAP7_75t_L g3158 ( 
.A(n_2758),
.B(n_2483),
.Y(n_3158)
);

NOR2xp33_ASAP7_75t_SL g3159 ( 
.A(n_2557),
.B(n_2563),
.Y(n_3159)
);

INVx1_ASAP7_75t_SL g3160 ( 
.A(n_2838),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2890),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2890),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_2893),
.Y(n_3163)
);

INVxp67_ASAP7_75t_L g3164 ( 
.A(n_2750),
.Y(n_3164)
);

INVx1_ASAP7_75t_SL g3165 ( 
.A(n_2917),
.Y(n_3165)
);

INVx2_ASAP7_75t_L g3166 ( 
.A(n_2550),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2893),
.Y(n_3167)
);

BUFx3_ASAP7_75t_L g3168 ( 
.A(n_2775),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_2894),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2894),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2903),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_2550),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2903),
.Y(n_3173)
);

CKINVDCx20_ASAP7_75t_R g3174 ( 
.A(n_2706),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2905),
.Y(n_3175)
);

INVx2_ASAP7_75t_L g3176 ( 
.A(n_2551),
.Y(n_3176)
);

AND2x2_ASAP7_75t_L g3177 ( 
.A(n_2767),
.B(n_1836),
.Y(n_3177)
);

CKINVDCx5p33_ASAP7_75t_R g3178 ( 
.A(n_2874),
.Y(n_3178)
);

INVxp33_ASAP7_75t_L g3179 ( 
.A(n_2899),
.Y(n_3179)
);

INVx2_ASAP7_75t_L g3180 ( 
.A(n_2551),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_2905),
.Y(n_3181)
);

NOR2xp33_ASAP7_75t_L g3182 ( 
.A(n_2758),
.B(n_1821),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_2909),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_L g3184 ( 
.A(n_2635),
.B(n_2683),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_2909),
.Y(n_3185)
);

INVxp33_ASAP7_75t_L g3186 ( 
.A(n_2859),
.Y(n_3186)
);

INVxp33_ASAP7_75t_L g3187 ( 
.A(n_2805),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2911),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2911),
.Y(n_3189)
);

CKINVDCx16_ASAP7_75t_R g3190 ( 
.A(n_2706),
.Y(n_3190)
);

AOI21x1_ASAP7_75t_L g3191 ( 
.A1(n_2732),
.A2(n_2659),
.B(n_2852),
.Y(n_3191)
);

AND2x2_ASAP7_75t_L g3192 ( 
.A(n_2767),
.B(n_1836),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_2915),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_2915),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_2920),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2920),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_2921),
.Y(n_3197)
);

NAND2xp33_ASAP7_75t_R g3198 ( 
.A(n_2706),
.B(n_2803),
.Y(n_3198)
);

AND2x4_ASAP7_75t_L g3199 ( 
.A(n_2803),
.B(n_2347),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_2921),
.Y(n_3200)
);

XNOR2xp5_ASAP7_75t_L g3201 ( 
.A(n_2888),
.B(n_2796),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_2761),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_2753),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_2635),
.B(n_2146),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_2753),
.Y(n_3205)
);

XOR2x2_ASAP7_75t_L g3206 ( 
.A(n_2814),
.B(n_1769),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_2754),
.Y(n_3207)
);

CKINVDCx20_ASAP7_75t_R g3208 ( 
.A(n_2803),
.Y(n_3208)
);

BUFx3_ASAP7_75t_L g3209 ( 
.A(n_2803),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_2754),
.Y(n_3210)
);

AND2x4_ASAP7_75t_L g3211 ( 
.A(n_2616),
.B(n_2124),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_2755),
.Y(n_3212)
);

INVx2_ASAP7_75t_L g3213 ( 
.A(n_2553),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_L g3214 ( 
.A(n_2635),
.B(n_2146),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_2755),
.Y(n_3215)
);

INVx4_ASAP7_75t_SL g3216 ( 
.A(n_2856),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_2759),
.Y(n_3217)
);

INVxp33_ASAP7_75t_L g3218 ( 
.A(n_2805),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_2759),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_2764),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_2764),
.Y(n_3221)
);

AND2x2_ASAP7_75t_L g3222 ( 
.A(n_2797),
.B(n_1838),
.Y(n_3222)
);

BUFx12f_ASAP7_75t_L g3223 ( 
.A(n_2873),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_2766),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_L g3225 ( 
.A(n_2683),
.B(n_2178),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_2766),
.Y(n_3226)
);

NOR2xp33_ASAP7_75t_L g3227 ( 
.A(n_2702),
.B(n_2272),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_2768),
.Y(n_3228)
);

NAND2xp5_ASAP7_75t_SL g3229 ( 
.A(n_2668),
.B(n_2064),
.Y(n_3229)
);

NOR2xp33_ASAP7_75t_L g3230 ( 
.A(n_2783),
.B(n_2128),
.Y(n_3230)
);

INVxp67_ASAP7_75t_L g3231 ( 
.A(n_2797),
.Y(n_3231)
);

INVxp33_ASAP7_75t_L g3232 ( 
.A(n_2567),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_2768),
.Y(n_3233)
);

XNOR2xp5_ASAP7_75t_L g3234 ( 
.A(n_2601),
.B(n_1769),
.Y(n_3234)
);

CKINVDCx5p33_ASAP7_75t_R g3235 ( 
.A(n_2874),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_L g3236 ( 
.A(n_2683),
.B(n_2178),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_2771),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_2771),
.Y(n_3238)
);

NOR2xp67_ASAP7_75t_L g3239 ( 
.A(n_2638),
.B(n_1927),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_2553),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_2554),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_2554),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_2558),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_2558),
.Y(n_3244)
);

CKINVDCx20_ASAP7_75t_R g3245 ( 
.A(n_2873),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_2559),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_2559),
.Y(n_3247)
);

CKINVDCx5p33_ASAP7_75t_R g3248 ( 
.A(n_2874),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_2561),
.Y(n_3249)
);

NOR2xp33_ASAP7_75t_L g3250 ( 
.A(n_2792),
.B(n_2129),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_2698),
.B(n_2246),
.Y(n_3251)
);

CKINVDCx20_ASAP7_75t_R g3252 ( 
.A(n_2616),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_2561),
.Y(n_3253)
);

AND2x2_ASAP7_75t_L g3254 ( 
.A(n_2798),
.B(n_1838),
.Y(n_3254)
);

AND2x2_ASAP7_75t_L g3255 ( 
.A(n_2798),
.B(n_1840),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_2571),
.Y(n_3256)
);

NAND2x1p5_ASAP7_75t_L g3257 ( 
.A(n_2585),
.B(n_2147),
.Y(n_3257)
);

AND2x2_ASAP7_75t_L g3258 ( 
.A(n_2808),
.B(n_1840),
.Y(n_3258)
);

XNOR2xp5_ASAP7_75t_L g3259 ( 
.A(n_2560),
.B(n_1792),
.Y(n_3259)
);

AND2x2_ASAP7_75t_L g3260 ( 
.A(n_2808),
.B(n_1880),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_2571),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_2572),
.Y(n_3262)
);

XOR2xp5_ASAP7_75t_L g3263 ( 
.A(n_2917),
.B(n_2256),
.Y(n_3263)
);

INVxp67_ASAP7_75t_SL g3264 ( 
.A(n_2580),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_2572),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_2574),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_2574),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_2576),
.Y(n_3268)
);

HB1xp67_ASAP7_75t_L g3269 ( 
.A(n_2918),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_2576),
.Y(n_3270)
);

CKINVDCx14_ASAP7_75t_R g3271 ( 
.A(n_2816),
.Y(n_3271)
);

AND2x2_ASAP7_75t_L g3272 ( 
.A(n_2816),
.B(n_1880),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_2578),
.Y(n_3273)
);

AND2x4_ASAP7_75t_L g3274 ( 
.A(n_2751),
.B(n_2133),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_2578),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_2582),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_2582),
.Y(n_3277)
);

INVx2_ASAP7_75t_L g3278 ( 
.A(n_2583),
.Y(n_3278)
);

AND2x4_ASAP7_75t_L g3279 ( 
.A(n_2751),
.B(n_2246),
.Y(n_3279)
);

AND2x2_ASAP7_75t_L g3280 ( 
.A(n_2831),
.B(n_1884),
.Y(n_3280)
);

NOR2xp67_ASAP7_75t_L g3281 ( 
.A(n_2729),
.B(n_2064),
.Y(n_3281)
);

NOR2xp33_ASAP7_75t_L g3282 ( 
.A(n_2585),
.B(n_2289),
.Y(n_3282)
);

AND2x2_ASAP7_75t_L g3283 ( 
.A(n_2831),
.B(n_1884),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_2583),
.Y(n_3284)
);

BUFx3_ASAP7_75t_L g3285 ( 
.A(n_2786),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_SL g3286 ( 
.A(n_2668),
.B(n_2064),
.Y(n_3286)
);

BUFx6f_ASAP7_75t_SL g3287 ( 
.A(n_2786),
.Y(n_3287)
);

CKINVDCx20_ASAP7_75t_R g3288 ( 
.A(n_2812),
.Y(n_3288)
);

INVx2_ASAP7_75t_L g3289 ( 
.A(n_2586),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_2586),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_2588),
.Y(n_3291)
);

AND2x2_ASAP7_75t_L g3292 ( 
.A(n_2918),
.B(n_1886),
.Y(n_3292)
);

AND2x2_ASAP7_75t_L g3293 ( 
.A(n_2516),
.B(n_1886),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_2588),
.Y(n_3294)
);

BUFx6f_ASAP7_75t_L g3295 ( 
.A(n_2547),
.Y(n_3295)
);

NOR2xp33_ASAP7_75t_L g3296 ( 
.A(n_2589),
.B(n_2289),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_L g3297 ( 
.A(n_2698),
.B(n_2259),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_2593),
.Y(n_3298)
);

AND2x2_ASAP7_75t_L g3299 ( 
.A(n_2507),
.B(n_2064),
.Y(n_3299)
);

XOR2xp5_ASAP7_75t_L g3300 ( 
.A(n_2654),
.B(n_2318),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_2593),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_2595),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_2595),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_2597),
.Y(n_3304)
);

AND2x2_ASAP7_75t_L g3305 ( 
.A(n_2651),
.B(n_2467),
.Y(n_3305)
);

INVx2_ASAP7_75t_L g3306 ( 
.A(n_2597),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_2603),
.Y(n_3307)
);

INVx1_ASAP7_75t_L g3308 ( 
.A(n_2603),
.Y(n_3308)
);

INVx2_ASAP7_75t_L g3309 ( 
.A(n_2611),
.Y(n_3309)
);

NOR2xp33_ASAP7_75t_L g3310 ( 
.A(n_2589),
.B(n_2606),
.Y(n_3310)
);

AND2x4_ASAP7_75t_L g3311 ( 
.A(n_2606),
.B(n_2259),
.Y(n_3311)
);

INVx2_ASAP7_75t_SL g3312 ( 
.A(n_2910),
.Y(n_3312)
);

NOR2xp33_ASAP7_75t_L g3313 ( 
.A(n_2581),
.B(n_2260),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_2611),
.Y(n_3314)
);

INVx2_ASAP7_75t_L g3315 ( 
.A(n_2617),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_2617),
.Y(n_3316)
);

INVx2_ASAP7_75t_SL g3317 ( 
.A(n_2910),
.Y(n_3317)
);

INVx2_ASAP7_75t_L g3318 ( 
.A(n_2619),
.Y(n_3318)
);

NOR2xp33_ASAP7_75t_L g3319 ( 
.A(n_2552),
.B(n_2260),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_2619),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_2621),
.Y(n_3321)
);

NAND2x1p5_ASAP7_75t_L g3322 ( 
.A(n_2506),
.B(n_2243),
.Y(n_3322)
);

OAI21xp5_ASAP7_75t_L g3323 ( 
.A1(n_2733),
.A2(n_2188),
.B(n_1946),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_SL g3324 ( 
.A(n_2677),
.B(n_2377),
.Y(n_3324)
);

AND2x2_ASAP7_75t_L g3325 ( 
.A(n_2815),
.B(n_1821),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_2621),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_2626),
.Y(n_3327)
);

CKINVDCx20_ASAP7_75t_R g3328 ( 
.A(n_2812),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_2626),
.Y(n_3329)
);

BUFx3_ASAP7_75t_L g3330 ( 
.A(n_2929),
.Y(n_3330)
);

NOR2xp33_ASAP7_75t_L g3331 ( 
.A(n_2556),
.B(n_2269),
.Y(n_3331)
);

HB1xp67_ASAP7_75t_L g3332 ( 
.A(n_2698),
.Y(n_3332)
);

INVx1_ASAP7_75t_L g3333 ( 
.A(n_2628),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_2628),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_2630),
.Y(n_3335)
);

AOI21xp5_ASAP7_75t_L g3336 ( 
.A1(n_2733),
.A2(n_1954),
.B(n_1933),
.Y(n_3336)
);

BUFx6f_ASAP7_75t_L g3337 ( 
.A(n_2547),
.Y(n_3337)
);

XOR2xp5_ASAP7_75t_L g3338 ( 
.A(n_2569),
.B(n_2318),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_2630),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_2632),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_2632),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_2633),
.Y(n_3342)
);

NOR2xp33_ASAP7_75t_L g3343 ( 
.A(n_2532),
.B(n_2269),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_2633),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_2634),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_2634),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_2637),
.Y(n_3347)
);

INVx1_ASAP7_75t_L g3348 ( 
.A(n_2637),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_2715),
.B(n_2274),
.Y(n_3349)
);

INVx4_ASAP7_75t_L g3350 ( 
.A(n_2557),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_2653),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_2653),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_2671),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_2671),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_2673),
.Y(n_3355)
);

BUFx6f_ASAP7_75t_SL g3356 ( 
.A(n_2856),
.Y(n_3356)
);

BUFx3_ASAP7_75t_L g3357 ( 
.A(n_2929),
.Y(n_3357)
);

XOR2xp5_ASAP7_75t_L g3358 ( 
.A(n_2672),
.B(n_2318),
.Y(n_3358)
);

AND2x2_ASAP7_75t_L g3359 ( 
.A(n_2726),
.B(n_1479),
.Y(n_3359)
);

AND2x2_ASAP7_75t_L g3360 ( 
.A(n_2784),
.B(n_1480),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_2673),
.Y(n_3361)
);

CKINVDCx20_ASAP7_75t_R g3362 ( 
.A(n_2674),
.Y(n_3362)
);

XNOR2xp5_ASAP7_75t_L g3363 ( 
.A(n_2541),
.B(n_1792),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_2681),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_2681),
.Y(n_3365)
);

INVx1_ASAP7_75t_L g3366 ( 
.A(n_2685),
.Y(n_3366)
);

XOR2x2_ASAP7_75t_L g3367 ( 
.A(n_2919),
.B(n_1797),
.Y(n_3367)
);

AND2x2_ASAP7_75t_L g3368 ( 
.A(n_2688),
.B(n_1481),
.Y(n_3368)
);

NOR2xp33_ASAP7_75t_L g3369 ( 
.A(n_2532),
.B(n_2274),
.Y(n_3369)
);

INVxp33_ASAP7_75t_L g3370 ( 
.A(n_2724),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_2685),
.Y(n_3371)
);

CKINVDCx5p33_ASAP7_75t_R g3372 ( 
.A(n_2677),
.Y(n_3372)
);

NOR2xp33_ASAP7_75t_SL g3373 ( 
.A(n_2557),
.B(n_2488),
.Y(n_3373)
);

INVxp67_ASAP7_75t_L g3374 ( 
.A(n_2856),
.Y(n_3374)
);

XOR2xp5_ASAP7_75t_L g3375 ( 
.A(n_2670),
.B(n_1797),
.Y(n_3375)
);

INVx2_ASAP7_75t_L g3376 ( 
.A(n_2687),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_2687),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_2690),
.Y(n_3378)
);

NOR2xp33_ASAP7_75t_L g3379 ( 
.A(n_2743),
.B(n_2331),
.Y(n_3379)
);

BUFx6f_ASAP7_75t_L g3380 ( 
.A(n_2547),
.Y(n_3380)
);

CKINVDCx20_ASAP7_75t_R g3381 ( 
.A(n_2743),
.Y(n_3381)
);

OR2x2_ASAP7_75t_SL g3382 ( 
.A(n_2772),
.B(n_1804),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_2690),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_2692),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_SL g3385 ( 
.A(n_3114),
.B(n_2769),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_L g3386 ( 
.A(n_3012),
.B(n_2715),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_3012),
.B(n_2715),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_L g3388 ( 
.A(n_2964),
.B(n_2856),
.Y(n_3388)
);

AND2x6_ASAP7_75t_SL g3389 ( 
.A(n_3182),
.B(n_1804),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_2964),
.B(n_2856),
.Y(n_3390)
);

AND2x4_ASAP7_75t_L g3391 ( 
.A(n_3216),
.B(n_2769),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_2941),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_SL g3393 ( 
.A(n_3232),
.B(n_2841),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_2944),
.Y(n_3394)
);

NOR2xp33_ASAP7_75t_L g3395 ( 
.A(n_3089),
.B(n_1918),
.Y(n_3395)
);

NOR2xp33_ASAP7_75t_L g3396 ( 
.A(n_2945),
.B(n_1918),
.Y(n_3396)
);

INVx2_ASAP7_75t_L g3397 ( 
.A(n_2949),
.Y(n_3397)
);

INVx3_ASAP7_75t_L g3398 ( 
.A(n_3350),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_3028),
.B(n_2856),
.Y(n_3399)
);

OAI22x1_ASAP7_75t_SL g3400 ( 
.A1(n_3059),
.A2(n_1098),
.B1(n_1126),
.B2(n_1092),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_3028),
.B(n_2773),
.Y(n_3401)
);

AND2x6_ASAP7_75t_L g3402 ( 
.A(n_3159),
.B(n_3216),
.Y(n_3402)
);

AND2x2_ASAP7_75t_L g3403 ( 
.A(n_2940),
.B(n_1482),
.Y(n_3403)
);

INVx2_ASAP7_75t_L g3404 ( 
.A(n_2953),
.Y(n_3404)
);

O2A1O1Ixp33_ASAP7_75t_L g3405 ( 
.A1(n_2945),
.A2(n_2631),
.B(n_2656),
.C(n_2652),
.Y(n_3405)
);

NOR2x1p5_ASAP7_75t_L g3406 ( 
.A(n_3072),
.B(n_2488),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_3049),
.B(n_2773),
.Y(n_3407)
);

INVx4_ASAP7_75t_L g3408 ( 
.A(n_3287),
.Y(n_3408)
);

AND2x2_ASAP7_75t_L g3409 ( 
.A(n_2951),
.B(n_1484),
.Y(n_3409)
);

O2A1O1Ixp5_ASAP7_75t_L g3410 ( 
.A1(n_2976),
.A2(n_2824),
.B(n_2659),
.C(n_2852),
.Y(n_3410)
);

AOI22xp33_ASAP7_75t_L g3411 ( 
.A1(n_3027),
.A2(n_2996),
.B1(n_2969),
.B2(n_3067),
.Y(n_3411)
);

INVxp67_ASAP7_75t_L g3412 ( 
.A(n_2955),
.Y(n_3412)
);

INVxp67_ASAP7_75t_L g3413 ( 
.A(n_2971),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_L g3414 ( 
.A(n_3049),
.B(n_2777),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3202),
.B(n_2777),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_L g3416 ( 
.A(n_2969),
.B(n_2778),
.Y(n_3416)
);

AOI22xp5_ASAP7_75t_L g3417 ( 
.A1(n_2981),
.A2(n_2599),
.B1(n_2712),
.B2(n_2709),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_L g3418 ( 
.A(n_3058),
.B(n_2778),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_3058),
.B(n_2781),
.Y(n_3419)
);

INVx2_ASAP7_75t_L g3420 ( 
.A(n_2974),
.Y(n_3420)
);

NOR2xp33_ASAP7_75t_SL g3421 ( 
.A(n_3015),
.B(n_2488),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_2950),
.Y(n_3422)
);

AND2x2_ASAP7_75t_L g3423 ( 
.A(n_2973),
.B(n_1486),
.Y(n_3423)
);

INVx2_ASAP7_75t_SL g3424 ( 
.A(n_2965),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_2947),
.B(n_2781),
.Y(n_3425)
);

INVx2_ASAP7_75t_L g3426 ( 
.A(n_2989),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_SL g3427 ( 
.A(n_2971),
.B(n_2841),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_L g3428 ( 
.A(n_2947),
.B(n_2782),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_2954),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_2957),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_L g3431 ( 
.A(n_2956),
.B(n_2782),
.Y(n_3431)
);

NOR2xp33_ASAP7_75t_L g3432 ( 
.A(n_3179),
.B(n_1978),
.Y(n_3432)
);

OAI22xp5_ASAP7_75t_L g3433 ( 
.A1(n_2976),
.A2(n_2544),
.B1(n_2907),
.B2(n_2867),
.Y(n_3433)
);

NAND2xp5_ASAP7_75t_L g3434 ( 
.A(n_2956),
.B(n_2785),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_2959),
.Y(n_3435)
);

AO221x1_ASAP7_75t_L g3436 ( 
.A1(n_2939),
.A2(n_1226),
.B1(n_2623),
.B2(n_2646),
.C(n_2547),
.Y(n_3436)
);

BUFx8_ASAP7_75t_L g3437 ( 
.A(n_3287),
.Y(n_3437)
);

NOR2xp33_ASAP7_75t_L g3438 ( 
.A(n_3003),
.B(n_3009),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_SL g3439 ( 
.A(n_3007),
.B(n_3040),
.Y(n_3439)
);

BUFx3_ASAP7_75t_L g3440 ( 
.A(n_3252),
.Y(n_3440)
);

NOR2xp33_ASAP7_75t_L g3441 ( 
.A(n_3007),
.B(n_3040),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_2960),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_L g3443 ( 
.A(n_2992),
.B(n_3134),
.Y(n_3443)
);

INVx8_ASAP7_75t_L g3444 ( 
.A(n_3356),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_L g3445 ( 
.A(n_2992),
.B(n_2867),
.Y(n_3445)
);

AND2x2_ASAP7_75t_L g3446 ( 
.A(n_3057),
.B(n_1488),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_SL g3447 ( 
.A(n_3060),
.B(n_2907),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_L g3448 ( 
.A(n_3093),
.B(n_2599),
.Y(n_3448)
);

INVx2_ASAP7_75t_L g3449 ( 
.A(n_2995),
.Y(n_3449)
);

NAND3xp33_ASAP7_75t_L g3450 ( 
.A(n_3093),
.B(n_3019),
.C(n_3021),
.Y(n_3450)
);

NOR2xp33_ASAP7_75t_L g3451 ( 
.A(n_3060),
.B(n_1978),
.Y(n_3451)
);

BUFx8_ASAP7_75t_L g3452 ( 
.A(n_3084),
.Y(n_3452)
);

BUFx6f_ASAP7_75t_SL g3453 ( 
.A(n_3199),
.Y(n_3453)
);

NOR3xp33_ASAP7_75t_L g3454 ( 
.A(n_3325),
.B(n_1228),
.C(n_1227),
.Y(n_3454)
);

INVx2_ASAP7_75t_SL g3455 ( 
.A(n_3223),
.Y(n_3455)
);

BUFx3_ASAP7_75t_L g3456 ( 
.A(n_3063),
.Y(n_3456)
);

AND2x2_ASAP7_75t_L g3457 ( 
.A(n_3032),
.B(n_1489),
.Y(n_3457)
);

NOR2xp33_ASAP7_75t_L g3458 ( 
.A(n_3075),
.B(n_2904),
.Y(n_3458)
);

INVxp67_ASAP7_75t_SL g3459 ( 
.A(n_3099),
.Y(n_3459)
);

INVxp67_ASAP7_75t_L g3460 ( 
.A(n_3055),
.Y(n_3460)
);

NOR2xp33_ASAP7_75t_L g3461 ( 
.A(n_3025),
.B(n_2745),
.Y(n_3461)
);

AOI21xp5_ASAP7_75t_L g3462 ( 
.A1(n_3024),
.A2(n_2684),
.B(n_2622),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_2961),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_L g3464 ( 
.A(n_3054),
.B(n_2800),
.Y(n_3464)
);

AOI21xp5_ASAP7_75t_L g3465 ( 
.A1(n_3024),
.A2(n_2684),
.B(n_2622),
.Y(n_3465)
);

INVxp67_ASAP7_75t_L g3466 ( 
.A(n_3001),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_L g3467 ( 
.A(n_3054),
.B(n_2785),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_2963),
.Y(n_3468)
);

INVx2_ASAP7_75t_L g3469 ( 
.A(n_3018),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_L g3470 ( 
.A(n_3164),
.B(n_2790),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_L g3471 ( 
.A(n_3164),
.B(n_2790),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_L g3472 ( 
.A(n_3139),
.B(n_2791),
.Y(n_3472)
);

INVx2_ASAP7_75t_L g3473 ( 
.A(n_3041),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_SL g3474 ( 
.A(n_3002),
.B(n_2623),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_SL g3475 ( 
.A(n_2946),
.B(n_2623),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_3231),
.B(n_2791),
.Y(n_3476)
);

BUFx4_ASAP7_75t_L g3477 ( 
.A(n_3015),
.Y(n_3477)
);

O2A1O1Ixp33_ASAP7_75t_L g3478 ( 
.A1(n_3019),
.A2(n_2934),
.B(n_2839),
.C(n_2854),
.Y(n_3478)
);

NAND2xp5_ASAP7_75t_SL g3479 ( 
.A(n_3160),
.B(n_2623),
.Y(n_3479)
);

AOI22xp5_ASAP7_75t_L g3480 ( 
.A1(n_2990),
.A2(n_1196),
.B1(n_1221),
.B2(n_1150),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_SL g3481 ( 
.A(n_3160),
.B(n_2948),
.Y(n_3481)
);

INVx2_ASAP7_75t_L g3482 ( 
.A(n_3070),
.Y(n_3482)
);

NOR2xp33_ASAP7_75t_L g3483 ( 
.A(n_3029),
.B(n_2748),
.Y(n_3483)
);

INVx8_ASAP7_75t_L g3484 ( 
.A(n_3356),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_2966),
.Y(n_3485)
);

NOR2xp33_ASAP7_75t_L g3486 ( 
.A(n_2978),
.B(n_2819),
.Y(n_3486)
);

NAND3xp33_ASAP7_75t_L g3487 ( 
.A(n_3021),
.B(n_2495),
.C(n_2437),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_2967),
.Y(n_3488)
);

AOI22xp33_ASAP7_75t_L g3489 ( 
.A1(n_3116),
.A2(n_1248),
.B1(n_1250),
.B2(n_2936),
.Y(n_3489)
);

AOI22xp33_ASAP7_75t_L g3490 ( 
.A1(n_3101),
.A2(n_2936),
.B1(n_2557),
.B2(n_2587),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_SL g3491 ( 
.A(n_2991),
.B(n_2623),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_SL g3492 ( 
.A(n_2991),
.B(n_2646),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_SL g3493 ( 
.A(n_3091),
.B(n_2646),
.Y(n_3493)
);

O2A1O1Ixp5_ASAP7_75t_L g3494 ( 
.A1(n_3120),
.A2(n_2738),
.B(n_2744),
.C(n_2735),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_L g3495 ( 
.A(n_3231),
.B(n_2793),
.Y(n_3495)
);

NOR2xp33_ASAP7_75t_L g3496 ( 
.A(n_3165),
.B(n_1885),
.Y(n_3496)
);

INVx2_ASAP7_75t_L g3497 ( 
.A(n_3104),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_2970),
.Y(n_3498)
);

AND2x2_ASAP7_75t_L g3499 ( 
.A(n_3165),
.B(n_1490),
.Y(n_3499)
);

NAND3xp33_ASAP7_75t_L g3500 ( 
.A(n_3004),
.B(n_2495),
.C(n_2437),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_L g3501 ( 
.A(n_3222),
.B(n_2800),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_2972),
.Y(n_3502)
);

BUFx8_ASAP7_75t_L g3503 ( 
.A(n_3109),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_L g3504 ( 
.A(n_3254),
.B(n_2793),
.Y(n_3504)
);

INVx3_ASAP7_75t_L g3505 ( 
.A(n_3350),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_L g3506 ( 
.A(n_3255),
.B(n_2788),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_SL g3507 ( 
.A(n_3372),
.B(n_2646),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_2977),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_SL g3509 ( 
.A(n_2952),
.B(n_2646),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_L g3510 ( 
.A(n_3258),
.B(n_2810),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_3260),
.B(n_2789),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_L g3512 ( 
.A(n_3272),
.B(n_2528),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_2980),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_3280),
.B(n_2528),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_SL g3515 ( 
.A(n_2952),
.B(n_2655),
.Y(n_3515)
);

NAND2xp5_ASAP7_75t_L g3516 ( 
.A(n_3283),
.B(n_2528),
.Y(n_3516)
);

BUFx3_ASAP7_75t_L g3517 ( 
.A(n_3381),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_SL g3518 ( 
.A(n_3136),
.B(n_2655),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_SL g3519 ( 
.A(n_3239),
.B(n_3143),
.Y(n_3519)
);

INVx2_ASAP7_75t_L g3520 ( 
.A(n_3113),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_3269),
.B(n_2826),
.Y(n_3521)
);

HB1xp67_ASAP7_75t_L g3522 ( 
.A(n_3269),
.Y(n_3522)
);

NOR2xp33_ASAP7_75t_L g3523 ( 
.A(n_3071),
.B(n_1885),
.Y(n_3523)
);

INVx2_ASAP7_75t_SL g3524 ( 
.A(n_2958),
.Y(n_3524)
);

NOR2xp33_ASAP7_75t_L g3525 ( 
.A(n_2984),
.B(n_2855),
.Y(n_3525)
);

NAND2xp5_ASAP7_75t_L g3526 ( 
.A(n_3293),
.B(n_2863),
.Y(n_3526)
);

OAI22xp33_ASAP7_75t_L g3527 ( 
.A1(n_3186),
.A2(n_2936),
.B1(n_2563),
.B2(n_2607),
.Y(n_3527)
);

AOI22xp33_ASAP7_75t_L g3528 ( 
.A1(n_3305),
.A2(n_2936),
.B1(n_2587),
.B2(n_2607),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_3133),
.B(n_2898),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_L g3530 ( 
.A(n_3151),
.B(n_2887),
.Y(n_3530)
);

AOI22xp5_ASAP7_75t_L g3531 ( 
.A1(n_3288),
.A2(n_2896),
.B1(n_2675),
.B2(n_2680),
.Y(n_3531)
);

INVx2_ASAP7_75t_SL g3532 ( 
.A(n_3094),
.Y(n_3532)
);

INVx2_ASAP7_75t_L g3533 ( 
.A(n_3118),
.Y(n_3533)
);

BUFx12f_ASAP7_75t_L g3534 ( 
.A(n_2962),
.Y(n_3534)
);

HB1xp67_ASAP7_75t_L g3535 ( 
.A(n_3271),
.Y(n_3535)
);

AND2x6_ASAP7_75t_SL g3536 ( 
.A(n_3034),
.B(n_1227),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_2982),
.Y(n_3537)
);

NAND2xp5_ASAP7_75t_SL g3538 ( 
.A(n_3051),
.B(n_2731),
.Y(n_3538)
);

NOR2xp33_ASAP7_75t_SL g3539 ( 
.A(n_3373),
.B(n_2563),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_2988),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3099),
.B(n_2692),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_3264),
.B(n_2694),
.Y(n_3542)
);

INVx1_ASAP7_75t_L g3543 ( 
.A(n_2997),
.Y(n_3543)
);

NAND2xp33_ASAP7_75t_L g3544 ( 
.A(n_3033),
.B(n_2563),
.Y(n_3544)
);

AND2x2_ASAP7_75t_L g3545 ( 
.A(n_3177),
.B(n_1491),
.Y(n_3545)
);

A2O1A1Ixp33_ASAP7_75t_L g3546 ( 
.A1(n_2993),
.A2(n_2895),
.B(n_2836),
.C(n_2876),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_SL g3547 ( 
.A(n_3085),
.B(n_2655),
.Y(n_3547)
);

INVx2_ASAP7_75t_SL g3548 ( 
.A(n_3149),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_3264),
.B(n_3079),
.Y(n_3549)
);

AOI22xp5_ASAP7_75t_L g3550 ( 
.A1(n_3328),
.A2(n_2423),
.B1(n_2607),
.B2(n_2587),
.Y(n_3550)
);

INVx2_ASAP7_75t_SL g3551 ( 
.A(n_3168),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_L g3552 ( 
.A(n_3079),
.B(n_2694),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_2998),
.Y(n_3553)
);

BUFx6f_ASAP7_75t_SL g3554 ( 
.A(n_3199),
.Y(n_3554)
);

NOR2xp33_ASAP7_75t_L g3555 ( 
.A(n_3187),
.B(n_2804),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_SL g3556 ( 
.A(n_3107),
.B(n_2655),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_L g3557 ( 
.A(n_3016),
.B(n_2695),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3000),
.Y(n_3558)
);

HB1xp67_ASAP7_75t_L g3559 ( 
.A(n_2975),
.Y(n_3559)
);

NOR2xp33_ASAP7_75t_L g3560 ( 
.A(n_3218),
.B(n_2804),
.Y(n_3560)
);

NOR2xp67_ASAP7_75t_L g3561 ( 
.A(n_3147),
.B(n_2845),
.Y(n_3561)
);

INVxp67_ASAP7_75t_L g3562 ( 
.A(n_3052),
.Y(n_3562)
);

NAND3xp33_ASAP7_75t_L g3563 ( 
.A(n_3004),
.B(n_2895),
.C(n_2188),
.Y(n_3563)
);

INVx2_ASAP7_75t_L g3564 ( 
.A(n_3125),
.Y(n_3564)
);

BUFx8_ASAP7_75t_L g3565 ( 
.A(n_3100),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_L g3566 ( 
.A(n_3016),
.B(n_2695),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_L g3567 ( 
.A(n_2993),
.B(n_2696),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_L g3568 ( 
.A(n_3097),
.B(n_2696),
.Y(n_3568)
);

NAND2xp5_ASAP7_75t_L g3569 ( 
.A(n_3098),
.B(n_2697),
.Y(n_3569)
);

OAI22xp33_ASAP7_75t_L g3570 ( 
.A1(n_3373),
.A2(n_2587),
.B1(n_2833),
.B2(n_2607),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_SL g3571 ( 
.A(n_3100),
.B(n_2655),
.Y(n_3571)
);

NAND2x1p5_ASAP7_75t_L g3572 ( 
.A(n_3279),
.B(n_2932),
.Y(n_3572)
);

NOR2xp33_ASAP7_75t_L g3573 ( 
.A(n_3227),
.B(n_2804),
.Y(n_3573)
);

INVx2_ASAP7_75t_L g3574 ( 
.A(n_3127),
.Y(n_3574)
);

INVx2_ASAP7_75t_L g3575 ( 
.A(n_3148),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3103),
.B(n_3105),
.Y(n_3576)
);

AOI21xp5_ASAP7_75t_L g3577 ( 
.A1(n_3155),
.A2(n_2779),
.B(n_2738),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_L g3578 ( 
.A(n_3110),
.B(n_2697),
.Y(n_3578)
);

OAI22xp5_ASAP7_75t_L g3579 ( 
.A1(n_3138),
.A2(n_2833),
.B1(n_2377),
.B2(n_2485),
.Y(n_3579)
);

AOI21x1_ASAP7_75t_L g3580 ( 
.A1(n_3154),
.A2(n_3191),
.B(n_3336),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_L g3581 ( 
.A(n_3111),
.B(n_2700),
.Y(n_3581)
);

INVx2_ASAP7_75t_SL g3582 ( 
.A(n_3285),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_3112),
.B(n_3119),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_L g3584 ( 
.A(n_3121),
.B(n_2700),
.Y(n_3584)
);

NAND3xp33_ASAP7_75t_L g3585 ( 
.A(n_3011),
.B(n_2073),
.C(n_2183),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3122),
.B(n_2701),
.Y(n_3586)
);

NOR2xp67_ASAP7_75t_L g3587 ( 
.A(n_3201),
.B(n_2845),
.Y(n_3587)
);

NOR2xp33_ASAP7_75t_L g3588 ( 
.A(n_3227),
.B(n_2813),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_3005),
.Y(n_3589)
);

NOR2xp33_ASAP7_75t_L g3590 ( 
.A(n_2942),
.B(n_2813),
.Y(n_3590)
);

INVx1_ASAP7_75t_L g3591 ( 
.A(n_3006),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_L g3592 ( 
.A(n_3123),
.B(n_3128),
.Y(n_3592)
);

NOR2xp33_ASAP7_75t_L g3593 ( 
.A(n_2943),
.B(n_2813),
.Y(n_3593)
);

NOR2xp33_ASAP7_75t_L g3594 ( 
.A(n_2979),
.B(n_2828),
.Y(n_3594)
);

AND2x6_ASAP7_75t_L g3595 ( 
.A(n_3159),
.B(n_3216),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_3130),
.B(n_2701),
.Y(n_3596)
);

OAI22xp5_ASAP7_75t_SL g3597 ( 
.A1(n_3124),
.A2(n_1244),
.B1(n_818),
.B2(n_819),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3008),
.Y(n_3598)
);

OAI22xp5_ASAP7_75t_L g3599 ( 
.A1(n_3141),
.A2(n_3144),
.B1(n_3145),
.B2(n_3142),
.Y(n_3599)
);

AOI22xp33_ASAP7_75t_L g3600 ( 
.A1(n_3014),
.A2(n_2833),
.B1(n_2423),
.B2(n_2787),
.Y(n_3600)
);

INVxp67_ASAP7_75t_SL g3601 ( 
.A(n_2938),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3010),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_3017),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_SL g3604 ( 
.A(n_3036),
.B(n_2731),
.Y(n_3604)
);

INVx1_ASAP7_75t_L g3605 ( 
.A(n_3023),
.Y(n_3605)
);

CKINVDCx5p33_ASAP7_75t_R g3606 ( 
.A(n_3013),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3135),
.B(n_2703),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_3146),
.B(n_2703),
.Y(n_3608)
);

NOR2xp33_ASAP7_75t_L g3609 ( 
.A(n_2999),
.B(n_2828),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_SL g3610 ( 
.A(n_3036),
.B(n_2770),
.Y(n_3610)
);

AOI22xp33_ASAP7_75t_L g3611 ( 
.A1(n_3014),
.A2(n_2833),
.B1(n_2423),
.B2(n_2787),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3026),
.Y(n_3612)
);

INVx2_ASAP7_75t_L g3613 ( 
.A(n_3166),
.Y(n_3613)
);

INVx2_ASAP7_75t_L g3614 ( 
.A(n_3172),
.Y(n_3614)
);

NOR2xp33_ASAP7_75t_L g3615 ( 
.A(n_3370),
.B(n_2828),
.Y(n_3615)
);

BUFx6f_ASAP7_75t_L g3616 ( 
.A(n_2938),
.Y(n_3616)
);

INVx2_ASAP7_75t_L g3617 ( 
.A(n_3176),
.Y(n_3617)
);

INVx2_ASAP7_75t_L g3618 ( 
.A(n_3180),
.Y(n_3618)
);

INVx2_ASAP7_75t_L g3619 ( 
.A(n_3213),
.Y(n_3619)
);

NAND2xp33_ASAP7_75t_L g3620 ( 
.A(n_3033),
.B(n_2568),
.Y(n_3620)
);

NOR2xp33_ASAP7_75t_L g3621 ( 
.A(n_3056),
.B(n_2830),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_L g3622 ( 
.A(n_3192),
.B(n_2707),
.Y(n_3622)
);

AO22x1_ASAP7_75t_L g3623 ( 
.A1(n_3178),
.A2(n_2423),
.B1(n_2055),
.B2(n_2045),
.Y(n_3623)
);

INVx2_ASAP7_75t_L g3624 ( 
.A(n_3278),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_SL g3625 ( 
.A(n_3037),
.B(n_2770),
.Y(n_3625)
);

INVx2_ASAP7_75t_L g3626 ( 
.A(n_3289),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_L g3627 ( 
.A(n_3360),
.B(n_2707),
.Y(n_3627)
);

INVxp67_ASAP7_75t_L g3628 ( 
.A(n_3158),
.Y(n_3628)
);

INVx1_ASAP7_75t_SL g3629 ( 
.A(n_3245),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_L g3630 ( 
.A(n_3292),
.B(n_2710),
.Y(n_3630)
);

INVx2_ASAP7_75t_L g3631 ( 
.A(n_3306),
.Y(n_3631)
);

NOR2xp33_ASAP7_75t_L g3632 ( 
.A(n_3056),
.B(n_3037),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_3011),
.B(n_2710),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_3030),
.Y(n_3634)
);

INVx2_ASAP7_75t_L g3635 ( 
.A(n_3309),
.Y(n_3635)
);

NAND3xp33_ASAP7_75t_L g3636 ( 
.A(n_3129),
.B(n_2073),
.C(n_2184),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_L g3637 ( 
.A(n_3035),
.B(n_2714),
.Y(n_3637)
);

INVx1_ASAP7_75t_L g3638 ( 
.A(n_3038),
.Y(n_3638)
);

NAND2xp5_ASAP7_75t_L g3639 ( 
.A(n_3035),
.B(n_2714),
.Y(n_3639)
);

NOR2xp67_ASAP7_75t_L g3640 ( 
.A(n_3235),
.B(n_2845),
.Y(n_3640)
);

INVxp67_ASAP7_75t_L g3641 ( 
.A(n_3158),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_L g3642 ( 
.A(n_3132),
.B(n_2716),
.Y(n_3642)
);

AND2x2_ASAP7_75t_L g3643 ( 
.A(n_3190),
.B(n_1492),
.Y(n_3643)
);

INVx8_ASAP7_75t_L g3644 ( 
.A(n_3046),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_SL g3645 ( 
.A(n_3279),
.B(n_2731),
.Y(n_3645)
);

INVx2_ASAP7_75t_L g3646 ( 
.A(n_3315),
.Y(n_3646)
);

INVx1_ASAP7_75t_L g3647 ( 
.A(n_3042),
.Y(n_3647)
);

NAND2xp5_ASAP7_75t_L g3648 ( 
.A(n_3132),
.B(n_2716),
.Y(n_3648)
);

INVx1_ASAP7_75t_L g3649 ( 
.A(n_3044),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_SL g3650 ( 
.A(n_3310),
.B(n_2731),
.Y(n_3650)
);

INVx2_ASAP7_75t_L g3651 ( 
.A(n_3318),
.Y(n_3651)
);

INVx6_ASAP7_75t_L g3652 ( 
.A(n_3211),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_L g3653 ( 
.A(n_3129),
.B(n_2719),
.Y(n_3653)
);

INVx2_ASAP7_75t_L g3654 ( 
.A(n_3371),
.Y(n_3654)
);

OAI22xp5_ASAP7_75t_L g3655 ( 
.A1(n_3152),
.A2(n_2472),
.B1(n_2485),
.B2(n_2851),
.Y(n_3655)
);

OAI22xp5_ASAP7_75t_L g3656 ( 
.A1(n_3153),
.A2(n_2472),
.B1(n_2869),
.B2(n_2851),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_SL g3657 ( 
.A(n_3310),
.B(n_2770),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_L g3658 ( 
.A(n_3096),
.B(n_2719),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_3045),
.Y(n_3659)
);

INVx2_ASAP7_75t_L g3660 ( 
.A(n_3376),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_L g3661 ( 
.A(n_3096),
.B(n_2730),
.Y(n_3661)
);

CKINVDCx5p33_ASAP7_75t_R g3662 ( 
.A(n_3039),
.Y(n_3662)
);

INVx1_ASAP7_75t_L g3663 ( 
.A(n_3047),
.Y(n_3663)
);

AOI22xp5_ASAP7_75t_L g3664 ( 
.A1(n_3362),
.A2(n_2423),
.B1(n_2913),
.B2(n_2897),
.Y(n_3664)
);

INVx2_ASAP7_75t_SL g3665 ( 
.A(n_3248),
.Y(n_3665)
);

OAI22xp33_ASAP7_75t_L g3666 ( 
.A1(n_3088),
.A2(n_821),
.B1(n_827),
.B2(n_815),
.Y(n_3666)
);

NAND2xp5_ASAP7_75t_L g3667 ( 
.A(n_3156),
.B(n_2730),
.Y(n_3667)
);

A2O1A1Ixp33_ASAP7_75t_L g3668 ( 
.A1(n_3282),
.A2(n_2830),
.B(n_2331),
.C(n_2185),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_L g3669 ( 
.A(n_3157),
.B(n_2580),
.Y(n_3669)
);

INVx3_ASAP7_75t_L g3670 ( 
.A(n_2938),
.Y(n_3670)
);

NOR2xp33_ASAP7_75t_L g3671 ( 
.A(n_3300),
.B(n_2830),
.Y(n_3671)
);

INVxp67_ASAP7_75t_L g3672 ( 
.A(n_3263),
.Y(n_3672)
);

INVx2_ASAP7_75t_SL g3673 ( 
.A(n_3209),
.Y(n_3673)
);

NOR2xp33_ASAP7_75t_L g3674 ( 
.A(n_3234),
.B(n_2922),
.Y(n_3674)
);

HB1xp67_ASAP7_75t_L g3675 ( 
.A(n_3117),
.Y(n_3675)
);

INVx1_ASAP7_75t_L g3676 ( 
.A(n_3050),
.Y(n_3676)
);

INVx1_ASAP7_75t_L g3677 ( 
.A(n_3053),
.Y(n_3677)
);

NAND2xp5_ASAP7_75t_L g3678 ( 
.A(n_3161),
.B(n_2584),
.Y(n_3678)
);

NAND2xp5_ASAP7_75t_L g3679 ( 
.A(n_3162),
.B(n_2584),
.Y(n_3679)
);

INVxp67_ASAP7_75t_SL g3680 ( 
.A(n_2968),
.Y(n_3680)
);

AND2x2_ASAP7_75t_L g3681 ( 
.A(n_3359),
.B(n_1496),
.Y(n_3681)
);

AND2x2_ASAP7_75t_L g3682 ( 
.A(n_3368),
.B(n_1498),
.Y(n_3682)
);

OAI221xp5_ASAP7_75t_L g3683 ( 
.A1(n_3126),
.A2(n_1237),
.B1(n_1242),
.B2(n_1235),
.C(n_1228),
.Y(n_3683)
);

NAND2xp5_ASAP7_75t_SL g3684 ( 
.A(n_3374),
.B(n_2731),
.Y(n_3684)
);

NAND3xp33_ASAP7_75t_L g3685 ( 
.A(n_3343),
.B(n_2073),
.C(n_2191),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_SL g3686 ( 
.A(n_3374),
.B(n_2770),
.Y(n_3686)
);

NOR2xp33_ASAP7_75t_L g3687 ( 
.A(n_3313),
.B(n_2925),
.Y(n_3687)
);

INVx2_ASAP7_75t_SL g3688 ( 
.A(n_3090),
.Y(n_3688)
);

NAND2xp5_ASAP7_75t_L g3689 ( 
.A(n_3163),
.B(n_3167),
.Y(n_3689)
);

AOI22xp5_ASAP7_75t_L g3690 ( 
.A1(n_3140),
.A2(n_3115),
.B1(n_3106),
.B2(n_3206),
.Y(n_3690)
);

NAND2xp5_ASAP7_75t_L g3691 ( 
.A(n_3169),
.B(n_2508),
.Y(n_3691)
);

OR2x6_ASAP7_75t_L g3692 ( 
.A(n_3311),
.B(n_2506),
.Y(n_3692)
);

AOI22xp33_ASAP7_75t_L g3693 ( 
.A1(n_3299),
.A2(n_2774),
.B1(n_2795),
.B2(n_2794),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_SL g3694 ( 
.A(n_3343),
.B(n_2770),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_L g3695 ( 
.A(n_3170),
.B(n_2508),
.Y(n_3695)
);

BUFx2_ASAP7_75t_L g3696 ( 
.A(n_3074),
.Y(n_3696)
);

NOR2xp33_ASAP7_75t_L g3697 ( 
.A(n_3313),
.B(n_2935),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_L g3698 ( 
.A(n_3171),
.B(n_2509),
.Y(n_3698)
);

NAND2xp5_ASAP7_75t_L g3699 ( 
.A(n_3173),
.B(n_3175),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3061),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_L g3701 ( 
.A(n_3181),
.B(n_2509),
.Y(n_3701)
);

INVx1_ASAP7_75t_L g3702 ( 
.A(n_3062),
.Y(n_3702)
);

OR2x2_ASAP7_75t_L g3703 ( 
.A(n_3064),
.B(n_2192),
.Y(n_3703)
);

AND2x2_ASAP7_75t_L g3704 ( 
.A(n_3117),
.B(n_1502),
.Y(n_3704)
);

NAND2xp5_ASAP7_75t_L g3705 ( 
.A(n_3183),
.B(n_2519),
.Y(n_3705)
);

NAND2xp5_ASAP7_75t_SL g3706 ( 
.A(n_3369),
.B(n_2877),
.Y(n_3706)
);

AND2x2_ASAP7_75t_SL g3707 ( 
.A(n_3198),
.B(n_2717),
.Y(n_3707)
);

NOR2xp33_ASAP7_75t_R g3708 ( 
.A(n_3043),
.B(n_2928),
.Y(n_3708)
);

INVx2_ASAP7_75t_L g3709 ( 
.A(n_2983),
.Y(n_3709)
);

INVx2_ASAP7_75t_SL g3710 ( 
.A(n_3330),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_L g3711 ( 
.A(n_3185),
.B(n_3188),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_L g3712 ( 
.A(n_3189),
.B(n_2519),
.Y(n_3712)
);

OAI221xp5_ASAP7_75t_L g3713 ( 
.A1(n_3363),
.A2(n_1242),
.B1(n_1249),
.B2(n_1237),
.C(n_1235),
.Y(n_3713)
);

NOR3xp33_ASAP7_75t_L g3714 ( 
.A(n_3066),
.B(n_1249),
.C(n_1234),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_3193),
.B(n_3194),
.Y(n_3715)
);

AND2x6_ASAP7_75t_L g3716 ( 
.A(n_2968),
.B(n_2774),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_SL g3717 ( 
.A(n_3369),
.B(n_3211),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3065),
.Y(n_3718)
);

INVx2_ASAP7_75t_L g3719 ( 
.A(n_2985),
.Y(n_3719)
);

AOI21xp5_ASAP7_75t_L g3720 ( 
.A1(n_3155),
.A2(n_2779),
.B(n_2744),
.Y(n_3720)
);

INVx2_ASAP7_75t_L g3721 ( 
.A(n_2986),
.Y(n_3721)
);

AND2x2_ASAP7_75t_L g3722 ( 
.A(n_3367),
.B(n_1503),
.Y(n_3722)
);

OR2x2_ASAP7_75t_L g3723 ( 
.A(n_3068),
.B(n_2199),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3195),
.Y(n_3724)
);

NOR2xp33_ASAP7_75t_L g3725 ( 
.A(n_3066),
.B(n_2832),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3196),
.Y(n_3726)
);

O2A1O1Ixp5_ASAP7_75t_L g3727 ( 
.A1(n_3154),
.A2(n_2746),
.B(n_2735),
.C(n_2851),
.Y(n_3727)
);

INVx2_ASAP7_75t_SL g3728 ( 
.A(n_3357),
.Y(n_3728)
);

NOR2xp33_ASAP7_75t_L g3729 ( 
.A(n_3230),
.B(n_2832),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_SL g3730 ( 
.A(n_3274),
.B(n_2877),
.Y(n_3730)
);

INVx2_ASAP7_75t_L g3731 ( 
.A(n_2987),
.Y(n_3731)
);

NAND2xp5_ASAP7_75t_L g3732 ( 
.A(n_3197),
.B(n_2801),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_L g3733 ( 
.A(n_3200),
.B(n_2801),
.Y(n_3733)
);

NOR2xp33_ASAP7_75t_L g3734 ( 
.A(n_3230),
.B(n_2842),
.Y(n_3734)
);

NAND2xp5_ASAP7_75t_L g3735 ( 
.A(n_3069),
.B(n_2802),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3073),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_L g3737 ( 
.A(n_3076),
.B(n_2802),
.Y(n_3737)
);

NAND2xp5_ASAP7_75t_SL g3738 ( 
.A(n_3274),
.B(n_2877),
.Y(n_3738)
);

NAND2xp5_ASAP7_75t_L g3739 ( 
.A(n_3332),
.B(n_2806),
.Y(n_3739)
);

INVx8_ASAP7_75t_L g3740 ( 
.A(n_3046),
.Y(n_3740)
);

BUFx3_ASAP7_75t_L g3741 ( 
.A(n_3174),
.Y(n_3741)
);

NAND2xp5_ASAP7_75t_L g3742 ( 
.A(n_3332),
.B(n_2806),
.Y(n_3742)
);

INVxp67_ASAP7_75t_L g3743 ( 
.A(n_3250),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3077),
.Y(n_3744)
);

NAND2xp5_ASAP7_75t_L g3745 ( 
.A(n_3031),
.B(n_2807),
.Y(n_3745)
);

NAND2xp5_ASAP7_75t_L g3746 ( 
.A(n_3031),
.B(n_2807),
.Y(n_3746)
);

NOR2xp33_ASAP7_75t_L g3747 ( 
.A(n_3250),
.B(n_2842),
.Y(n_3747)
);

OAI21xp33_ASAP7_75t_L g3748 ( 
.A1(n_3102),
.A2(n_832),
.B(n_831),
.Y(n_3748)
);

BUFx3_ASAP7_75t_L g3749 ( 
.A(n_3208),
.Y(n_3749)
);

NAND2xp5_ASAP7_75t_L g3750 ( 
.A(n_3020),
.B(n_2817),
.Y(n_3750)
);

OR2x2_ASAP7_75t_L g3751 ( 
.A(n_3078),
.B(n_2211),
.Y(n_3751)
);

AOI22xp33_ASAP7_75t_L g3752 ( 
.A1(n_3020),
.A2(n_2795),
.B1(n_2860),
.B2(n_2794),
.Y(n_3752)
);

NAND2xp5_ASAP7_75t_L g3753 ( 
.A(n_3020),
.B(n_3240),
.Y(n_3753)
);

NOR3xp33_ASAP7_75t_L g3754 ( 
.A(n_3312),
.B(n_1234),
.C(n_1188),
.Y(n_3754)
);

INVx2_ASAP7_75t_L g3755 ( 
.A(n_3241),
.Y(n_3755)
);

O2A1O1Ixp33_ASAP7_75t_L g3756 ( 
.A1(n_3102),
.A2(n_1506),
.B(n_1508),
.C(n_1505),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3080),
.Y(n_3757)
);

NOR2xp33_ASAP7_75t_L g3758 ( 
.A(n_3317),
.B(n_2843),
.Y(n_3758)
);

NAND2xp5_ASAP7_75t_SL g3759 ( 
.A(n_3311),
.B(n_2877),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_3020),
.B(n_2817),
.Y(n_3760)
);

INVx2_ASAP7_75t_L g3761 ( 
.A(n_3242),
.Y(n_3761)
);

A2O1A1Ixp33_ASAP7_75t_L g3762 ( 
.A1(n_3282),
.A2(n_2218),
.B(n_2222),
.C(n_2219),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_L g3763 ( 
.A(n_3020),
.B(n_2818),
.Y(n_3763)
);

AND2x2_ASAP7_75t_L g3764 ( 
.A(n_3259),
.B(n_1509),
.Y(n_3764)
);

NAND2xp5_ASAP7_75t_L g3765 ( 
.A(n_3243),
.B(n_2818),
.Y(n_3765)
);

INVx2_ASAP7_75t_SL g3766 ( 
.A(n_3338),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_3081),
.Y(n_3767)
);

INVx2_ASAP7_75t_SL g3768 ( 
.A(n_3358),
.Y(n_3768)
);

AND2x2_ASAP7_75t_L g3769 ( 
.A(n_3082),
.B(n_1510),
.Y(n_3769)
);

INVx2_ASAP7_75t_L g3770 ( 
.A(n_3244),
.Y(n_3770)
);

INVx3_ASAP7_75t_L g3771 ( 
.A(n_2968),
.Y(n_3771)
);

NOR2xp33_ASAP7_75t_L g3772 ( 
.A(n_3083),
.B(n_2843),
.Y(n_3772)
);

NAND2xp5_ASAP7_75t_L g3773 ( 
.A(n_3246),
.B(n_2821),
.Y(n_3773)
);

NOR2xp67_ASAP7_75t_L g3774 ( 
.A(n_3086),
.B(n_2869),
.Y(n_3774)
);

BUFx3_ASAP7_75t_L g3775 ( 
.A(n_3382),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_SL g3776 ( 
.A(n_2994),
.B(n_2877),
.Y(n_3776)
);

NAND2xp5_ASAP7_75t_L g3777 ( 
.A(n_3247),
.B(n_2821),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3087),
.Y(n_3778)
);

NAND2xp5_ASAP7_75t_L g3779 ( 
.A(n_3249),
.B(n_2822),
.Y(n_3779)
);

NOR2xp33_ASAP7_75t_L g3780 ( 
.A(n_3092),
.B(n_2846),
.Y(n_3780)
);

NAND2xp33_ASAP7_75t_L g3781 ( 
.A(n_3033),
.B(n_2994),
.Y(n_3781)
);

INVxp67_ASAP7_75t_L g3782 ( 
.A(n_3095),
.Y(n_3782)
);

NAND2xp5_ASAP7_75t_SL g3783 ( 
.A(n_2994),
.B(n_2869),
.Y(n_3783)
);

NOR2xp33_ASAP7_75t_L g3784 ( 
.A(n_3375),
.B(n_2846),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_L g3785 ( 
.A(n_3253),
.B(n_2822),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_3203),
.Y(n_3786)
);

INVx2_ASAP7_75t_L g3787 ( 
.A(n_3256),
.Y(n_3787)
);

BUFx6f_ASAP7_75t_L g3788 ( 
.A(n_3022),
.Y(n_3788)
);

AOI22xp5_ASAP7_75t_L g3789 ( 
.A1(n_3296),
.A2(n_2848),
.B1(n_2861),
.B2(n_2858),
.Y(n_3789)
);

AND2x4_ASAP7_75t_SL g3790 ( 
.A(n_3022),
.B(n_2901),
.Y(n_3790)
);

NAND2x1p5_ASAP7_75t_L g3791 ( 
.A(n_3022),
.B(n_2568),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_L g3792 ( 
.A(n_3261),
.B(n_2827),
.Y(n_3792)
);

NAND2xp5_ASAP7_75t_L g3793 ( 
.A(n_3262),
.B(n_2827),
.Y(n_3793)
);

NAND2xp5_ASAP7_75t_L g3794 ( 
.A(n_3265),
.B(n_2829),
.Y(n_3794)
);

NOR2xp67_ASAP7_75t_L g3795 ( 
.A(n_3379),
.B(n_2901),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_L g3796 ( 
.A(n_3266),
.B(n_2829),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_L g3797 ( 
.A(n_3267),
.B(n_2860),
.Y(n_3797)
);

AO221x1_ASAP7_75t_L g3798 ( 
.A1(n_3048),
.A2(n_2930),
.B1(n_2928),
.B2(n_2901),
.C(n_2238),
.Y(n_3798)
);

BUFx2_ASAP7_75t_L g3799 ( 
.A(n_3440),
.Y(n_3799)
);

AOI21xp5_ASAP7_75t_L g3800 ( 
.A1(n_3620),
.A2(n_3323),
.B(n_3336),
.Y(n_3800)
);

INVx2_ASAP7_75t_L g3801 ( 
.A(n_3709),
.Y(n_3801)
);

NOR2xp33_ASAP7_75t_SL g3802 ( 
.A(n_3644),
.B(n_3046),
.Y(n_3802)
);

AO21x1_ASAP7_75t_L g3803 ( 
.A1(n_3448),
.A2(n_3296),
.B(n_3319),
.Y(n_3803)
);

HB1xp67_ASAP7_75t_L g3804 ( 
.A(n_3441),
.Y(n_3804)
);

NAND2xp5_ASAP7_75t_L g3805 ( 
.A(n_3443),
.B(n_3131),
.Y(n_3805)
);

NAND2xp5_ASAP7_75t_L g3806 ( 
.A(n_3628),
.B(n_3205),
.Y(n_3806)
);

AND2x2_ASAP7_75t_L g3807 ( 
.A(n_3411),
.B(n_1511),
.Y(n_3807)
);

NOR2xp33_ASAP7_75t_R g3808 ( 
.A(n_3606),
.B(n_3048),
.Y(n_3808)
);

CKINVDCx10_ASAP7_75t_R g3809 ( 
.A(n_3453),
.Y(n_3809)
);

OAI21x1_ASAP7_75t_L g3810 ( 
.A1(n_3580),
.A2(n_2746),
.B(n_3323),
.Y(n_3810)
);

AOI21xp5_ASAP7_75t_L g3811 ( 
.A1(n_3544),
.A2(n_3184),
.B(n_3204),
.Y(n_3811)
);

INVx1_ASAP7_75t_L g3812 ( 
.A(n_3392),
.Y(n_3812)
);

AOI21xp5_ASAP7_75t_L g3813 ( 
.A1(n_3450),
.A2(n_3184),
.B(n_3204),
.Y(n_3813)
);

OAI22xp5_ASAP7_75t_L g3814 ( 
.A1(n_3445),
.A2(n_3150),
.B1(n_3331),
.B2(n_3319),
.Y(n_3814)
);

AOI21xp5_ASAP7_75t_L g3815 ( 
.A1(n_3462),
.A2(n_3225),
.B(n_3214),
.Y(n_3815)
);

NAND2x1p5_ASAP7_75t_L g3816 ( 
.A(n_3391),
.B(n_3048),
.Y(n_3816)
);

BUFx6f_ASAP7_75t_L g3817 ( 
.A(n_3444),
.Y(n_3817)
);

INVx2_ASAP7_75t_L g3818 ( 
.A(n_3719),
.Y(n_3818)
);

OAI21xp33_ASAP7_75t_L g3819 ( 
.A1(n_3396),
.A2(n_3331),
.B(n_874),
.Y(n_3819)
);

AOI21xp5_ASAP7_75t_L g3820 ( 
.A1(n_3465),
.A2(n_3225),
.B(n_3214),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_L g3821 ( 
.A(n_3641),
.B(n_3207),
.Y(n_3821)
);

AOI21xp5_ASAP7_75t_L g3822 ( 
.A1(n_3781),
.A2(n_3251),
.B(n_3236),
.Y(n_3822)
);

OAI21xp33_ASAP7_75t_L g3823 ( 
.A1(n_3714),
.A2(n_875),
.B(n_854),
.Y(n_3823)
);

BUFx2_ASAP7_75t_L g3824 ( 
.A(n_3452),
.Y(n_3824)
);

AOI21x1_ASAP7_75t_L g3825 ( 
.A1(n_3577),
.A2(n_3286),
.B(n_3229),
.Y(n_3825)
);

NAND2xp5_ASAP7_75t_L g3826 ( 
.A(n_3743),
.B(n_3210),
.Y(n_3826)
);

OAI21xp5_ASAP7_75t_L g3827 ( 
.A1(n_3563),
.A2(n_3150),
.B(n_3236),
.Y(n_3827)
);

NAND2xp5_ASAP7_75t_L g3828 ( 
.A(n_3446),
.B(n_3212),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_3499),
.B(n_3215),
.Y(n_3829)
);

OAI21xp33_ASAP7_75t_L g3830 ( 
.A1(n_3416),
.A2(n_877),
.B(n_856),
.Y(n_3830)
);

INVx1_ASAP7_75t_SL g3831 ( 
.A(n_3652),
.Y(n_3831)
);

A2O1A1Ixp33_ASAP7_75t_L g3832 ( 
.A1(n_3417),
.A2(n_3379),
.B(n_3281),
.C(n_3324),
.Y(n_3832)
);

OAI21xp5_ASAP7_75t_L g3833 ( 
.A1(n_3388),
.A2(n_3297),
.B(n_3251),
.Y(n_3833)
);

OAI21xp33_ASAP7_75t_L g3834 ( 
.A1(n_3416),
.A2(n_882),
.B(n_861),
.Y(n_3834)
);

AOI21xp5_ASAP7_75t_L g3835 ( 
.A1(n_3459),
.A2(n_3349),
.B(n_3297),
.Y(n_3835)
);

AO21x1_ASAP7_75t_L g3836 ( 
.A1(n_3388),
.A2(n_3349),
.B(n_3219),
.Y(n_3836)
);

OAI21xp33_ASAP7_75t_L g3837 ( 
.A1(n_3748),
.A2(n_889),
.B(n_862),
.Y(n_3837)
);

AOI21xp5_ASAP7_75t_L g3838 ( 
.A1(n_3390),
.A2(n_2679),
.B(n_2524),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_L g3839 ( 
.A(n_3457),
.B(n_3217),
.Y(n_3839)
);

AOI21xp5_ASAP7_75t_L g3840 ( 
.A1(n_3390),
.A2(n_2679),
.B(n_2524),
.Y(n_3840)
);

INVx1_ASAP7_75t_SL g3841 ( 
.A(n_3652),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_L g3842 ( 
.A(n_3403),
.B(n_3220),
.Y(n_3842)
);

AOI21x1_ASAP7_75t_L g3843 ( 
.A1(n_3720),
.A2(n_2227),
.B(n_2224),
.Y(n_3843)
);

OAI22xp5_ASAP7_75t_L g3844 ( 
.A1(n_3573),
.A2(n_3295),
.B1(n_3337),
.B2(n_3137),
.Y(n_3844)
);

OAI21xp5_ASAP7_75t_L g3845 ( 
.A1(n_3725),
.A2(n_3621),
.B(n_3549),
.Y(n_3845)
);

INVx2_ASAP7_75t_SL g3846 ( 
.A(n_3437),
.Y(n_3846)
);

AOI21xp5_ASAP7_75t_L g3847 ( 
.A1(n_3549),
.A2(n_2679),
.B(n_2524),
.Y(n_3847)
);

AOI21xp5_ASAP7_75t_L g3848 ( 
.A1(n_3478),
.A2(n_2779),
.B(n_3137),
.Y(n_3848)
);

AOI21xp5_ASAP7_75t_L g3849 ( 
.A1(n_3425),
.A2(n_3295),
.B(n_3137),
.Y(n_3849)
);

NAND2xp5_ASAP7_75t_L g3850 ( 
.A(n_3409),
.B(n_3221),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_SL g3851 ( 
.A(n_3588),
.B(n_3399),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_L g3852 ( 
.A(n_3423),
.B(n_3224),
.Y(n_3852)
);

NAND2xp5_ASAP7_75t_SL g3853 ( 
.A(n_3399),
.B(n_3295),
.Y(n_3853)
);

AO21x1_ASAP7_75t_L g3854 ( 
.A1(n_3433),
.A2(n_3734),
.B(n_3729),
.Y(n_3854)
);

INVx1_ASAP7_75t_L g3855 ( 
.A(n_3394),
.Y(n_3855)
);

NAND2xp5_ASAP7_75t_SL g3856 ( 
.A(n_3632),
.B(n_3337),
.Y(n_3856)
);

AOI21xp5_ASAP7_75t_L g3857 ( 
.A1(n_3425),
.A2(n_3380),
.B(n_3337),
.Y(n_3857)
);

AOI21xp5_ASAP7_75t_L g3858 ( 
.A1(n_3428),
.A2(n_3434),
.B(n_3431),
.Y(n_3858)
);

BUFx10_ASAP7_75t_L g3859 ( 
.A(n_3662),
.Y(n_3859)
);

A2O1A1Ixp33_ASAP7_75t_L g3860 ( 
.A1(n_3405),
.A2(n_2239),
.B(n_2250),
.C(n_2249),
.Y(n_3860)
);

A2O1A1Ixp33_ASAP7_75t_L g3861 ( 
.A1(n_3687),
.A2(n_3697),
.B(n_3747),
.C(n_3454),
.Y(n_3861)
);

AOI21xp5_ASAP7_75t_L g3862 ( 
.A1(n_3428),
.A2(n_3434),
.B(n_3431),
.Y(n_3862)
);

HB1xp67_ASAP7_75t_L g3863 ( 
.A(n_3522),
.Y(n_3863)
);

AOI21xp5_ASAP7_75t_L g3864 ( 
.A1(n_3386),
.A2(n_3380),
.B(n_2577),
.Y(n_3864)
);

AND2x2_ASAP7_75t_L g3865 ( 
.A(n_3764),
.B(n_1513),
.Y(n_3865)
);

NAND2x1p5_ASAP7_75t_L g3866 ( 
.A(n_3391),
.B(n_3380),
.Y(n_3866)
);

NOR3xp33_ASAP7_75t_L g3867 ( 
.A(n_3713),
.B(n_1517),
.C(n_1516),
.Y(n_3867)
);

NAND2xp5_ASAP7_75t_L g3868 ( 
.A(n_3545),
.B(n_3226),
.Y(n_3868)
);

AOI21xp5_ASAP7_75t_L g3869 ( 
.A1(n_3386),
.A2(n_2577),
.B(n_3033),
.Y(n_3869)
);

OAI22xp5_ASAP7_75t_L g3870 ( 
.A1(n_3412),
.A2(n_2930),
.B1(n_2928),
.B2(n_846),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_3422),
.Y(n_3871)
);

NAND2xp5_ASAP7_75t_L g3872 ( 
.A(n_3704),
.B(n_3228),
.Y(n_3872)
);

AO21x1_ASAP7_75t_L g3873 ( 
.A1(n_3753),
.A2(n_3237),
.B(n_3233),
.Y(n_3873)
);

NAND2xp5_ASAP7_75t_SL g3874 ( 
.A(n_3594),
.B(n_3033),
.Y(n_3874)
);

AOI21xp5_ASAP7_75t_L g3875 ( 
.A1(n_3387),
.A2(n_2577),
.B(n_3033),
.Y(n_3875)
);

NAND2xp5_ASAP7_75t_L g3876 ( 
.A(n_3681),
.B(n_3682),
.Y(n_3876)
);

NOR2xp33_ASAP7_75t_L g3877 ( 
.A(n_3562),
.B(n_836),
.Y(n_3877)
);

NAND2xp5_ASAP7_75t_L g3878 ( 
.A(n_3413),
.B(n_3238),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_3429),
.Y(n_3879)
);

NOR2xp33_ASAP7_75t_L g3880 ( 
.A(n_3590),
.B(n_850),
.Y(n_3880)
);

AOI21xp5_ASAP7_75t_L g3881 ( 
.A1(n_3387),
.A2(n_2930),
.B(n_2857),
.Y(n_3881)
);

AOI21xp5_ASAP7_75t_L g3882 ( 
.A1(n_3401),
.A2(n_2857),
.B(n_2848),
.Y(n_3882)
);

AND2x2_ASAP7_75t_L g3883 ( 
.A(n_3643),
.B(n_1520),
.Y(n_3883)
);

AOI21xp5_ASAP7_75t_L g3884 ( 
.A1(n_3401),
.A2(n_2861),
.B(n_2858),
.Y(n_3884)
);

AOI21xp5_ASAP7_75t_L g3885 ( 
.A1(n_3541),
.A2(n_2872),
.B(n_2870),
.Y(n_3885)
);

OAI21xp5_ASAP7_75t_L g3886 ( 
.A1(n_3410),
.A2(n_3108),
.B(n_3046),
.Y(n_3886)
);

NAND2xp5_ASAP7_75t_L g3887 ( 
.A(n_3675),
.B(n_3268),
.Y(n_3887)
);

BUFx8_ASAP7_75t_L g3888 ( 
.A(n_3534),
.Y(n_3888)
);

AOI21xp5_ASAP7_75t_L g3889 ( 
.A1(n_3541),
.A2(n_2872),
.B(n_2870),
.Y(n_3889)
);

NAND2xp5_ASAP7_75t_L g3890 ( 
.A(n_3472),
.B(n_3270),
.Y(n_3890)
);

O2A1O1Ixp33_ASAP7_75t_L g3891 ( 
.A1(n_3666),
.A2(n_1523),
.B(n_1524),
.C(n_1521),
.Y(n_3891)
);

BUFx6f_ASAP7_75t_L g3892 ( 
.A(n_3444),
.Y(n_3892)
);

NOR2xp33_ASAP7_75t_L g3893 ( 
.A(n_3593),
.B(n_851),
.Y(n_3893)
);

INVx1_ASAP7_75t_L g3894 ( 
.A(n_3430),
.Y(n_3894)
);

NAND2xp5_ASAP7_75t_L g3895 ( 
.A(n_3769),
.B(n_3273),
.Y(n_3895)
);

NAND2xp5_ASAP7_75t_SL g3896 ( 
.A(n_3424),
.B(n_2879),
.Y(n_3896)
);

NAND2xp5_ASAP7_75t_L g3897 ( 
.A(n_3438),
.B(n_3275),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_L g3898 ( 
.A(n_3627),
.B(n_3276),
.Y(n_3898)
);

AOI21xp5_ASAP7_75t_L g3899 ( 
.A1(n_3542),
.A2(n_2881),
.B(n_2879),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_L g3900 ( 
.A(n_3689),
.B(n_3277),
.Y(n_3900)
);

AOI21xp5_ASAP7_75t_L g3901 ( 
.A1(n_3542),
.A2(n_2883),
.B(n_2881),
.Y(n_3901)
);

AOI21xp5_ASAP7_75t_L g3902 ( 
.A1(n_3546),
.A2(n_2884),
.B(n_2883),
.Y(n_3902)
);

CKINVDCx5p33_ASAP7_75t_R g3903 ( 
.A(n_3437),
.Y(n_3903)
);

AND2x2_ASAP7_75t_L g3904 ( 
.A(n_3722),
.B(n_1528),
.Y(n_3904)
);

AOI21xp5_ASAP7_75t_L g3905 ( 
.A1(n_3494),
.A2(n_2889),
.B(n_2884),
.Y(n_3905)
);

AOI21xp5_ASAP7_75t_L g3906 ( 
.A1(n_3727),
.A2(n_3579),
.B(n_3552),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_L g3907 ( 
.A(n_3699),
.B(n_3284),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_L g3908 ( 
.A(n_3711),
.B(n_3290),
.Y(n_3908)
);

BUFx6f_ASAP7_75t_L g3909 ( 
.A(n_3444),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3435),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_L g3911 ( 
.A(n_3715),
.B(n_3291),
.Y(n_3911)
);

NAND2xp5_ASAP7_75t_L g3912 ( 
.A(n_3466),
.B(n_3294),
.Y(n_3912)
);

INVx2_ASAP7_75t_SL g3913 ( 
.A(n_3406),
.Y(n_3913)
);

INVx2_ASAP7_75t_L g3914 ( 
.A(n_3721),
.Y(n_3914)
);

OR2x2_ASAP7_75t_L g3915 ( 
.A(n_3559),
.B(n_3298),
.Y(n_3915)
);

NAND2xp5_ASAP7_75t_L g3916 ( 
.A(n_3460),
.B(n_3301),
.Y(n_3916)
);

AOI21xp5_ASAP7_75t_L g3917 ( 
.A1(n_3552),
.A2(n_2892),
.B(n_2889),
.Y(n_3917)
);

NOR2xp33_ASAP7_75t_L g3918 ( 
.A(n_3451),
.B(n_852),
.Y(n_3918)
);

O2A1O1Ixp33_ASAP7_75t_SL g3919 ( 
.A1(n_3547),
.A2(n_1985),
.B(n_1993),
.C(n_1963),
.Y(n_3919)
);

NAND2xp5_ASAP7_75t_L g3920 ( 
.A(n_3489),
.B(n_3302),
.Y(n_3920)
);

OAI21xp5_ASAP7_75t_L g3921 ( 
.A1(n_3512),
.A2(n_3108),
.B(n_3046),
.Y(n_3921)
);

NOR2xp33_ASAP7_75t_L g3922 ( 
.A(n_3481),
.B(n_868),
.Y(n_3922)
);

INVx3_ASAP7_75t_L g3923 ( 
.A(n_3644),
.Y(n_3923)
);

NOR2xp33_ASAP7_75t_L g3924 ( 
.A(n_3480),
.B(n_870),
.Y(n_3924)
);

NAND2xp5_ASAP7_75t_L g3925 ( 
.A(n_3782),
.B(n_3303),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_L g3926 ( 
.A(n_3439),
.B(n_3304),
.Y(n_3926)
);

AOI21xp5_ASAP7_75t_L g3927 ( 
.A1(n_3487),
.A2(n_2900),
.B(n_2892),
.Y(n_3927)
);

AOI21xp5_ASAP7_75t_L g3928 ( 
.A1(n_3642),
.A2(n_2902),
.B(n_2900),
.Y(n_3928)
);

BUFx4f_ASAP7_75t_L g3929 ( 
.A(n_3484),
.Y(n_3929)
);

AOI21xp5_ASAP7_75t_L g3930 ( 
.A1(n_3648),
.A2(n_2906),
.B(n_2902),
.Y(n_3930)
);

AOI21xp5_ASAP7_75t_L g3931 ( 
.A1(n_3653),
.A2(n_2912),
.B(n_2906),
.Y(n_3931)
);

CKINVDCx5p33_ASAP7_75t_R g3932 ( 
.A(n_3708),
.Y(n_3932)
);

OAI22xp5_ASAP7_75t_L g3933 ( 
.A1(n_3511),
.A2(n_873),
.B1(n_876),
.B2(n_871),
.Y(n_3933)
);

OAI21xp5_ASAP7_75t_L g3934 ( 
.A1(n_3514),
.A2(n_3108),
.B(n_2262),
.Y(n_3934)
);

NAND2xp5_ASAP7_75t_SL g3935 ( 
.A(n_3531),
.B(n_2912),
.Y(n_3935)
);

INVx2_ASAP7_75t_L g3936 ( 
.A(n_3731),
.Y(n_3936)
);

INVx2_ASAP7_75t_L g3937 ( 
.A(n_3755),
.Y(n_3937)
);

NOR2xp33_ASAP7_75t_L g3938 ( 
.A(n_3458),
.B(n_881),
.Y(n_3938)
);

NAND2xp5_ASAP7_75t_L g3939 ( 
.A(n_3724),
.B(n_3307),
.Y(n_3939)
);

O2A1O1Ixp33_ASAP7_75t_L g3940 ( 
.A1(n_3385),
.A2(n_1542),
.B(n_1544),
.C(n_1529),
.Y(n_3940)
);

AO21x1_ASAP7_75t_L g3941 ( 
.A1(n_3753),
.A2(n_3314),
.B(n_3308),
.Y(n_3941)
);

BUFx12f_ASAP7_75t_L g3942 ( 
.A(n_3452),
.Y(n_3942)
);

O2A1O1Ixp33_ASAP7_75t_L g3943 ( 
.A1(n_3683),
.A2(n_3530),
.B(n_3529),
.C(n_3395),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3442),
.Y(n_3944)
);

NOR2xp33_ASAP7_75t_L g3945 ( 
.A(n_3525),
.B(n_883),
.Y(n_3945)
);

A2O1A1Ixp33_ASAP7_75t_L g3946 ( 
.A1(n_3500),
.A2(n_2254),
.B(n_2265),
.C(n_2263),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_3463),
.Y(n_3947)
);

OAI21xp5_ASAP7_75t_L g3948 ( 
.A1(n_3516),
.A2(n_3108),
.B(n_2270),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_3726),
.B(n_3316),
.Y(n_3949)
);

AOI21xp5_ASAP7_75t_L g3950 ( 
.A1(n_3798),
.A2(n_2923),
.B(n_2914),
.Y(n_3950)
);

INVx3_ASAP7_75t_L g3951 ( 
.A(n_3644),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_L g3952 ( 
.A(n_3576),
.B(n_3320),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_L g3953 ( 
.A(n_3576),
.B(n_3321),
.Y(n_3953)
);

NAND2xp5_ASAP7_75t_SL g3954 ( 
.A(n_3506),
.B(n_2914),
.Y(n_3954)
);

AND2x2_ASAP7_75t_L g3955 ( 
.A(n_3784),
.B(n_1547),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3583),
.B(n_3326),
.Y(n_3956)
);

O2A1O1Ixp5_ASAP7_75t_L g3957 ( 
.A1(n_3507),
.A2(n_2933),
.B(n_2937),
.C(n_2923),
.Y(n_3957)
);

NAND2xp5_ASAP7_75t_L g3958 ( 
.A(n_3583),
.B(n_3592),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_L g3959 ( 
.A(n_3592),
.B(n_3327),
.Y(n_3959)
);

NOR2xp33_ASAP7_75t_L g3960 ( 
.A(n_3432),
.B(n_890),
.Y(n_3960)
);

NAND2xp5_ASAP7_75t_L g3961 ( 
.A(n_3496),
.B(n_3329),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_L g3962 ( 
.A(n_3468),
.B(n_3333),
.Y(n_3962)
);

OAI21xp5_ASAP7_75t_L g3963 ( 
.A1(n_3418),
.A2(n_3108),
.B(n_2271),
.Y(n_3963)
);

NOR2xp33_ASAP7_75t_L g3964 ( 
.A(n_3629),
.B(n_895),
.Y(n_3964)
);

AOI21xp5_ASAP7_75t_L g3965 ( 
.A1(n_3464),
.A2(n_2937),
.B(n_2933),
.Y(n_3965)
);

INVx3_ASAP7_75t_L g3966 ( 
.A(n_3740),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_3485),
.Y(n_3967)
);

AOI21xp5_ASAP7_75t_L g3968 ( 
.A1(n_3467),
.A2(n_3678),
.B(n_3669),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_L g3969 ( 
.A(n_3488),
.B(n_3334),
.Y(n_3969)
);

AOI21xp5_ASAP7_75t_L g3970 ( 
.A1(n_3679),
.A2(n_3339),
.B(n_3335),
.Y(n_3970)
);

NAND2xp5_ASAP7_75t_SL g3971 ( 
.A(n_3510),
.B(n_3340),
.Y(n_3971)
);

INVx2_ASAP7_75t_L g3972 ( 
.A(n_3761),
.Y(n_3972)
);

AND2x2_ASAP7_75t_L g3973 ( 
.A(n_3671),
.B(n_1549),
.Y(n_3973)
);

BUFx2_ASAP7_75t_SL g3974 ( 
.A(n_3408),
.Y(n_3974)
);

BUFx6f_ASAP7_75t_L g3975 ( 
.A(n_3484),
.Y(n_3975)
);

NAND2xp5_ASAP7_75t_SL g3976 ( 
.A(n_3717),
.B(n_3341),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_L g3977 ( 
.A(n_3498),
.B(n_3342),
.Y(n_3977)
);

AOI21xp5_ASAP7_75t_L g3978 ( 
.A1(n_3740),
.A2(n_3345),
.B(n_3344),
.Y(n_3978)
);

INVx1_ASAP7_75t_L g3979 ( 
.A(n_3502),
.Y(n_3979)
);

AOI21x1_ASAP7_75t_L g3980 ( 
.A1(n_3694),
.A2(n_2275),
.B(n_2266),
.Y(n_3980)
);

O2A1O1Ixp33_ASAP7_75t_L g3981 ( 
.A1(n_3393),
.A2(n_1555),
.B(n_1556),
.C(n_1552),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3508),
.Y(n_3982)
);

AOI21xp5_ASAP7_75t_L g3983 ( 
.A1(n_3740),
.A2(n_3347),
.B(n_3346),
.Y(n_3983)
);

OAI21xp5_ASAP7_75t_L g3984 ( 
.A1(n_3418),
.A2(n_2288),
.B(n_2276),
.Y(n_3984)
);

INVx2_ASAP7_75t_L g3985 ( 
.A(n_3770),
.Y(n_3985)
);

HB1xp67_ASAP7_75t_L g3986 ( 
.A(n_3517),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3513),
.Y(n_3987)
);

INVx2_ASAP7_75t_L g3988 ( 
.A(n_3787),
.Y(n_3988)
);

OAI21xp5_ASAP7_75t_L g3989 ( 
.A1(n_3419),
.A2(n_2291),
.B(n_2290),
.Y(n_3989)
);

INVx3_ASAP7_75t_L g3990 ( 
.A(n_3572),
.Y(n_3990)
);

NAND2xp5_ASAP7_75t_L g3991 ( 
.A(n_3537),
.B(n_3348),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3540),
.Y(n_3992)
);

NOR2xp33_ASAP7_75t_L g3993 ( 
.A(n_3652),
.B(n_897),
.Y(n_3993)
);

INVx2_ASAP7_75t_L g3994 ( 
.A(n_3397),
.Y(n_3994)
);

AND2x2_ASAP7_75t_L g3995 ( 
.A(n_3674),
.B(n_1557),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_SL g3996 ( 
.A(n_3555),
.B(n_3351),
.Y(n_3996)
);

A2O1A1Ixp33_ASAP7_75t_L g3997 ( 
.A1(n_3772),
.A2(n_2295),
.B(n_2302),
.C(n_2298),
.Y(n_3997)
);

INVx1_ASAP7_75t_L g3998 ( 
.A(n_3543),
.Y(n_3998)
);

AND2x2_ASAP7_75t_L g3999 ( 
.A(n_3741),
.B(n_1559),
.Y(n_3999)
);

AOI21xp5_ASAP7_75t_L g4000 ( 
.A1(n_3407),
.A2(n_3353),
.B(n_3352),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_3553),
.Y(n_4001)
);

AO21x1_ASAP7_75t_L g4002 ( 
.A1(n_3650),
.A2(n_3355),
.B(n_3354),
.Y(n_4002)
);

NAND2x1p5_ASAP7_75t_L g4003 ( 
.A(n_3509),
.B(n_3361),
.Y(n_4003)
);

INVx2_ASAP7_75t_L g4004 ( 
.A(n_3404),
.Y(n_4004)
);

OAI22xp5_ASAP7_75t_L g4005 ( 
.A1(n_3486),
.A2(n_899),
.B1(n_906),
.B2(n_898),
.Y(n_4005)
);

NAND2xp5_ASAP7_75t_SL g4006 ( 
.A(n_3560),
.B(n_3364),
.Y(n_4006)
);

A2O1A1Ixp33_ASAP7_75t_L g4007 ( 
.A1(n_3780),
.A2(n_2307),
.B(n_2314),
.C(n_2311),
.Y(n_4007)
);

AND2x2_ASAP7_75t_L g4008 ( 
.A(n_3749),
.B(n_1561),
.Y(n_4008)
);

OAI21xp33_ASAP7_75t_L g4009 ( 
.A1(n_3419),
.A2(n_935),
.B(n_923),
.Y(n_4009)
);

O2A1O1Ixp33_ASAP7_75t_L g4010 ( 
.A1(n_3521),
.A2(n_1567),
.B(n_1569),
.C(n_1562),
.Y(n_4010)
);

AND2x4_ASAP7_75t_L g4011 ( 
.A(n_3587),
.B(n_3365),
.Y(n_4011)
);

NOR2x1_ASAP7_75t_L g4012 ( 
.A(n_3408),
.B(n_2315),
.Y(n_4012)
);

AOI22xp33_ASAP7_75t_L g4013 ( 
.A1(n_3597),
.A2(n_3377),
.B1(n_3378),
.B2(n_3366),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_L g4014 ( 
.A(n_3558),
.B(n_3383),
.Y(n_4014)
);

INVxp67_ASAP7_75t_L g4015 ( 
.A(n_3503),
.Y(n_4015)
);

AOI21xp5_ASAP7_75t_L g4016 ( 
.A1(n_3407),
.A2(n_3384),
.B(n_2862),
.Y(n_4016)
);

NAND2xp5_ASAP7_75t_L g4017 ( 
.A(n_3589),
.B(n_907),
.Y(n_4017)
);

AND2x2_ASAP7_75t_L g4018 ( 
.A(n_3535),
.B(n_1571),
.Y(n_4018)
);

OAI21xp5_ASAP7_75t_L g4019 ( 
.A1(n_3668),
.A2(n_2320),
.B(n_2319),
.Y(n_4019)
);

NAND2xp5_ASAP7_75t_L g4020 ( 
.A(n_3591),
.B(n_3598),
.Y(n_4020)
);

AOI22xp5_ASAP7_75t_L g4021 ( 
.A1(n_3523),
.A2(n_916),
.B1(n_917),
.B2(n_908),
.Y(n_4021)
);

AOI21xp5_ASAP7_75t_L g4022 ( 
.A1(n_3414),
.A2(n_2862),
.B(n_2721),
.Y(n_4022)
);

INVx5_ASAP7_75t_L g4023 ( 
.A(n_3402),
.Y(n_4023)
);

OAI22xp5_ASAP7_75t_L g4024 ( 
.A1(n_3599),
.A2(n_925),
.B1(n_926),
.B2(n_919),
.Y(n_4024)
);

AOI21xp5_ASAP7_75t_L g4025 ( 
.A1(n_3414),
.A2(n_2721),
.B(n_2568),
.Y(n_4025)
);

NAND2xp5_ASAP7_75t_SL g4026 ( 
.A(n_3615),
.B(n_2281),
.Y(n_4026)
);

INVx11_ASAP7_75t_L g4027 ( 
.A(n_3503),
.Y(n_4027)
);

BUFx8_ASAP7_75t_L g4028 ( 
.A(n_3696),
.Y(n_4028)
);

BUFx6f_ASAP7_75t_L g4029 ( 
.A(n_3484),
.Y(n_4029)
);

INVx2_ASAP7_75t_L g4030 ( 
.A(n_3420),
.Y(n_4030)
);

INVx2_ASAP7_75t_SL g4031 ( 
.A(n_3477),
.Y(n_4031)
);

BUFx3_ASAP7_75t_L g4032 ( 
.A(n_3456),
.Y(n_4032)
);

AOI21xp5_ASAP7_75t_L g4033 ( 
.A1(n_3570),
.A2(n_2721),
.B(n_2568),
.Y(n_4033)
);

NAND2xp5_ASAP7_75t_L g4034 ( 
.A(n_3602),
.B(n_927),
.Y(n_4034)
);

INVx1_ASAP7_75t_L g4035 ( 
.A(n_3603),
.Y(n_4035)
);

AOI21xp5_ASAP7_75t_L g4036 ( 
.A1(n_3655),
.A2(n_2721),
.B(n_2568),
.Y(n_4036)
);

INVx4_ASAP7_75t_L g4037 ( 
.A(n_3616),
.Y(n_4037)
);

AOI21xp5_ASAP7_75t_L g4038 ( 
.A1(n_3739),
.A2(n_2725),
.B(n_2721),
.Y(n_4038)
);

AND2x2_ASAP7_75t_L g4039 ( 
.A(n_3461),
.B(n_1577),
.Y(n_4039)
);

NAND2xp5_ASAP7_75t_L g4040 ( 
.A(n_3605),
.B(n_928),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_L g4041 ( 
.A(n_3612),
.B(n_929),
.Y(n_4041)
);

OAI22xp5_ASAP7_75t_L g4042 ( 
.A1(n_3470),
.A2(n_3471),
.B1(n_3504),
.B2(n_3501),
.Y(n_4042)
);

AND2x2_ASAP7_75t_L g4043 ( 
.A(n_3483),
.B(n_1580),
.Y(n_4043)
);

NAND2xp5_ASAP7_75t_SL g4044 ( 
.A(n_3630),
.B(n_2281),
.Y(n_4044)
);

A2O1A1Ixp33_ASAP7_75t_L g4045 ( 
.A1(n_3756),
.A2(n_2323),
.B(n_2326),
.C(n_2325),
.Y(n_4045)
);

AOI21xp5_ASAP7_75t_L g4046 ( 
.A1(n_3739),
.A2(n_2756),
.B(n_2725),
.Y(n_4046)
);

AOI21xp5_ASAP7_75t_L g4047 ( 
.A1(n_3742),
.A2(n_2756),
.B(n_2725),
.Y(n_4047)
);

AND2x2_ASAP7_75t_L g4048 ( 
.A(n_3609),
.B(n_1582),
.Y(n_4048)
);

INVx2_ASAP7_75t_L g4049 ( 
.A(n_3426),
.Y(n_4049)
);

INVx2_ASAP7_75t_L g4050 ( 
.A(n_3449),
.Y(n_4050)
);

A2O1A1Ixp33_ASAP7_75t_L g4051 ( 
.A1(n_3622),
.A2(n_2327),
.B(n_2335),
.C(n_2330),
.Y(n_4051)
);

INVx2_ASAP7_75t_L g4052 ( 
.A(n_3469),
.Y(n_4052)
);

NAND2xp5_ASAP7_75t_SL g4053 ( 
.A(n_3616),
.B(n_2281),
.Y(n_4053)
);

INVxp67_ASAP7_75t_SL g4054 ( 
.A(n_3691),
.Y(n_4054)
);

AOI21x1_ASAP7_75t_L g4055 ( 
.A1(n_3706),
.A2(n_3657),
.B(n_3475),
.Y(n_4055)
);

INVx4_ASAP7_75t_L g4056 ( 
.A(n_3616),
.Y(n_4056)
);

AOI21xp5_ASAP7_75t_L g4057 ( 
.A1(n_3742),
.A2(n_2756),
.B(n_2725),
.Y(n_4057)
);

NAND2xp5_ASAP7_75t_SL g4058 ( 
.A(n_3788),
.B(n_2281),
.Y(n_4058)
);

INVxp67_ASAP7_75t_L g4059 ( 
.A(n_3582),
.Y(n_4059)
);

HB1xp67_ASAP7_75t_L g4060 ( 
.A(n_3634),
.Y(n_4060)
);

NAND2xp5_ASAP7_75t_L g4061 ( 
.A(n_3638),
.B(n_932),
.Y(n_4061)
);

OAI21xp5_ASAP7_75t_L g4062 ( 
.A1(n_3762),
.A2(n_2011),
.B(n_2003),
.Y(n_4062)
);

AOI33xp33_ASAP7_75t_L g4063 ( 
.A1(n_3647),
.A2(n_1588),
.A3(n_1585),
.B1(n_1591),
.B2(n_1586),
.B3(n_1583),
.Y(n_4063)
);

A2O1A1Ixp33_ASAP7_75t_L g4064 ( 
.A1(n_3774),
.A2(n_2339),
.B(n_2343),
.C(n_2340),
.Y(n_4064)
);

BUFx2_ASAP7_75t_L g4065 ( 
.A(n_3565),
.Y(n_4065)
);

OAI21x1_ASAP7_75t_L g4066 ( 
.A1(n_3567),
.A2(n_3322),
.B(n_2348),
.Y(n_4066)
);

INVx3_ASAP7_75t_L g4067 ( 
.A(n_3572),
.Y(n_4067)
);

NAND2xp5_ASAP7_75t_L g4068 ( 
.A(n_3649),
.B(n_933),
.Y(n_4068)
);

NAND2xp5_ASAP7_75t_L g4069 ( 
.A(n_3659),
.B(n_936),
.Y(n_4069)
);

NAND2xp5_ASAP7_75t_L g4070 ( 
.A(n_3663),
.B(n_939),
.Y(n_4070)
);

AOI21xp5_ASAP7_75t_L g4071 ( 
.A1(n_3567),
.A2(n_2756),
.B(n_2725),
.Y(n_4071)
);

A2O1A1Ixp33_ASAP7_75t_L g4072 ( 
.A1(n_3664),
.A2(n_2344),
.B(n_2351),
.C(n_2502),
.Y(n_4072)
);

A2O1A1Ixp33_ASAP7_75t_L g4073 ( 
.A1(n_3758),
.A2(n_3636),
.B(n_3526),
.C(n_3658),
.Y(n_4073)
);

AOI21xp5_ASAP7_75t_L g4074 ( 
.A1(n_3695),
.A2(n_2849),
.B(n_2756),
.Y(n_4074)
);

NAND2xp5_ASAP7_75t_L g4075 ( 
.A(n_3676),
.B(n_3677),
.Y(n_4075)
);

NAND2xp5_ASAP7_75t_L g4076 ( 
.A(n_3700),
.B(n_941),
.Y(n_4076)
);

AOI21x1_ASAP7_75t_L g4077 ( 
.A1(n_3685),
.A2(n_2418),
.B(n_2413),
.Y(n_4077)
);

BUFx6f_ASAP7_75t_L g4078 ( 
.A(n_3788),
.Y(n_4078)
);

INVx2_ASAP7_75t_L g4079 ( 
.A(n_3473),
.Y(n_4079)
);

NOR2xp33_ASAP7_75t_L g4080 ( 
.A(n_3688),
.B(n_3447),
.Y(n_4080)
);

NAND2xp5_ASAP7_75t_L g4081 ( 
.A(n_3702),
.B(n_944),
.Y(n_4081)
);

INVx2_ASAP7_75t_L g4082 ( 
.A(n_3482),
.Y(n_4082)
);

NAND2xp5_ASAP7_75t_SL g4083 ( 
.A(n_3788),
.B(n_2297),
.Y(n_4083)
);

NAND2xp5_ASAP7_75t_L g4084 ( 
.A(n_3718),
.B(n_945),
.Y(n_4084)
);

NAND2xp5_ASAP7_75t_SL g4085 ( 
.A(n_3661),
.B(n_3707),
.Y(n_4085)
);

AOI22xp5_ASAP7_75t_L g4086 ( 
.A1(n_3474),
.A2(n_3421),
.B1(n_3515),
.B2(n_3754),
.Y(n_4086)
);

AND2x2_ASAP7_75t_L g4087 ( 
.A(n_3736),
.B(n_1593),
.Y(n_4087)
);

OAI21xp5_ASAP7_75t_L g4088 ( 
.A1(n_3656),
.A2(n_1990),
.B(n_2151),
.Y(n_4088)
);

NAND2xp5_ASAP7_75t_SL g4089 ( 
.A(n_3550),
.B(n_3561),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_L g4090 ( 
.A(n_3744),
.B(n_951),
.Y(n_4090)
);

INVxp67_ASAP7_75t_L g4091 ( 
.A(n_3710),
.Y(n_4091)
);

NAND2xp5_ASAP7_75t_L g4092 ( 
.A(n_3757),
.B(n_953),
.Y(n_4092)
);

NAND2xp5_ASAP7_75t_L g4093 ( 
.A(n_3767),
.B(n_955),
.Y(n_4093)
);

NOR2xp33_ASAP7_75t_L g4094 ( 
.A(n_3427),
.B(n_958),
.Y(n_4094)
);

AOI21xp5_ASAP7_75t_L g4095 ( 
.A1(n_3698),
.A2(n_2932),
.B(n_2849),
.Y(n_4095)
);

NAND2xp5_ASAP7_75t_L g4096 ( 
.A(n_3778),
.B(n_962),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_3876),
.B(n_3565),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_SL g4098 ( 
.A(n_3845),
.B(n_3633),
.Y(n_4098)
);

AOI21xp5_ASAP7_75t_L g4099 ( 
.A1(n_3858),
.A2(n_3436),
.B(n_3776),
.Y(n_4099)
);

O2A1O1Ixp33_ASAP7_75t_L g4100 ( 
.A1(n_3861),
.A2(n_3519),
.B(n_3524),
.C(n_3491),
.Y(n_4100)
);

AOI21xp5_ASAP7_75t_L g4101 ( 
.A1(n_3862),
.A2(n_3705),
.B(n_3701),
.Y(n_4101)
);

NAND2xp5_ASAP7_75t_SL g4102 ( 
.A(n_3958),
.B(n_3795),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_4060),
.Y(n_4103)
);

NOR2xp33_ASAP7_75t_L g4104 ( 
.A(n_3938),
.B(n_3690),
.Y(n_4104)
);

AOI21xp5_ASAP7_75t_L g4105 ( 
.A1(n_3800),
.A2(n_3712),
.B(n_3750),
.Y(n_4105)
);

AOI21xp5_ASAP7_75t_L g4106 ( 
.A1(n_3886),
.A2(n_3968),
.B(n_3848),
.Y(n_4106)
);

O2A1O1Ixp33_ASAP7_75t_L g4107 ( 
.A1(n_3819),
.A2(n_3492),
.B(n_3518),
.C(n_3493),
.Y(n_4107)
);

NOR2xp33_ASAP7_75t_SL g4108 ( 
.A(n_3942),
.B(n_3453),
.Y(n_4108)
);

AND2x2_ASAP7_75t_L g4109 ( 
.A(n_3995),
.B(n_3728),
.Y(n_4109)
);

CKINVDCx8_ASAP7_75t_R g4110 ( 
.A(n_3809),
.Y(n_4110)
);

INVx2_ASAP7_75t_L g4111 ( 
.A(n_3801),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_L g4112 ( 
.A(n_3804),
.B(n_3786),
.Y(n_4112)
);

INVx3_ASAP7_75t_L g4113 ( 
.A(n_3929),
.Y(n_4113)
);

INVx1_ASAP7_75t_L g4114 ( 
.A(n_4020),
.Y(n_4114)
);

OAI22xp5_ASAP7_75t_L g4115 ( 
.A1(n_3945),
.A2(n_3495),
.B1(n_3476),
.B2(n_3490),
.Y(n_4115)
);

O2A1O1Ixp5_ASAP7_75t_L g4116 ( 
.A1(n_3854),
.A2(n_3556),
.B(n_3645),
.C(n_3730),
.Y(n_4116)
);

BUFx12f_ASAP7_75t_L g4117 ( 
.A(n_3888),
.Y(n_4117)
);

AOI21xp5_ASAP7_75t_L g4118 ( 
.A1(n_3886),
.A2(n_3760),
.B(n_3750),
.Y(n_4118)
);

AND2x4_ASAP7_75t_L g4119 ( 
.A(n_4023),
.B(n_3571),
.Y(n_4119)
);

AOI22x1_ASAP7_75t_L g4120 ( 
.A1(n_3813),
.A2(n_3932),
.B1(n_3799),
.B2(n_3875),
.Y(n_4120)
);

NOR2xp33_ASAP7_75t_L g4121 ( 
.A(n_3918),
.B(n_3389),
.Y(n_4121)
);

AOI22xp5_ASAP7_75t_L g4122 ( 
.A1(n_3880),
.A2(n_3400),
.B1(n_3766),
.B2(n_3768),
.Y(n_4122)
);

NAND2xp5_ASAP7_75t_L g4123 ( 
.A(n_3883),
.B(n_3637),
.Y(n_4123)
);

OAI22xp5_ASAP7_75t_L g4124 ( 
.A1(n_3960),
.A2(n_3532),
.B1(n_3551),
.B2(n_3548),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_4075),
.Y(n_4125)
);

NAND2xp5_ASAP7_75t_L g4126 ( 
.A(n_3807),
.B(n_3639),
.Y(n_4126)
);

AOI21xp5_ASAP7_75t_L g4127 ( 
.A1(n_3869),
.A2(n_3811),
.B(n_3906),
.Y(n_4127)
);

OAI22xp5_ASAP7_75t_L g4128 ( 
.A1(n_3893),
.A2(n_3528),
.B1(n_3665),
.B2(n_3640),
.Y(n_4128)
);

NOR2xp33_ASAP7_75t_L g4129 ( 
.A(n_3805),
.B(n_3672),
.Y(n_4129)
);

NAND2xp5_ASAP7_75t_L g4130 ( 
.A(n_3865),
.B(n_3673),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_3812),
.Y(n_4131)
);

OAI22xp5_ASAP7_75t_L g4132 ( 
.A1(n_3943),
.A2(n_3611),
.B1(n_3600),
.B2(n_3415),
.Y(n_4132)
);

NAND2xp5_ASAP7_75t_L g4133 ( 
.A(n_3973),
.B(n_3415),
.Y(n_4133)
);

BUFx10_ASAP7_75t_L g4134 ( 
.A(n_3903),
.Y(n_4134)
);

INVx8_ASAP7_75t_L g4135 ( 
.A(n_3817),
.Y(n_4135)
);

A2O1A1Ixp33_ASAP7_75t_L g4136 ( 
.A1(n_3830),
.A2(n_3834),
.B(n_3837),
.C(n_4009),
.Y(n_4136)
);

OAI22x1_ASAP7_75t_L g4137 ( 
.A1(n_4031),
.A2(n_3538),
.B1(n_3455),
.B2(n_3536),
.Y(n_4137)
);

OAI22x1_ASAP7_75t_L g4138 ( 
.A1(n_4086),
.A2(n_3479),
.B1(n_3738),
.B2(n_3789),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_L g4139 ( 
.A(n_4039),
.B(n_3608),
.Y(n_4139)
);

INVx2_ASAP7_75t_L g4140 ( 
.A(n_3818),
.Y(n_4140)
);

AOI21xp5_ASAP7_75t_L g4141 ( 
.A1(n_3847),
.A2(n_3763),
.B(n_3760),
.Y(n_4141)
);

AOI21xp33_ASAP7_75t_L g4142 ( 
.A1(n_4042),
.A2(n_3585),
.B(n_3763),
.Y(n_4142)
);

AOI21xp5_ASAP7_75t_L g4143 ( 
.A1(n_3921),
.A2(n_3608),
.B(n_3566),
.Y(n_4143)
);

NOR2xp33_ASAP7_75t_L g4144 ( 
.A(n_3986),
.B(n_3775),
.Y(n_4144)
);

INVx2_ASAP7_75t_L g4145 ( 
.A(n_3914),
.Y(n_4145)
);

BUFx2_ASAP7_75t_L g4146 ( 
.A(n_3808),
.Y(n_4146)
);

NAND2xp5_ASAP7_75t_L g4147 ( 
.A(n_4043),
.B(n_3703),
.Y(n_4147)
);

AOI21x1_ASAP7_75t_L g4148 ( 
.A1(n_3843),
.A2(n_3840),
.B(n_3838),
.Y(n_4148)
);

NAND2xp5_ASAP7_75t_L g4149 ( 
.A(n_3828),
.B(n_3497),
.Y(n_4149)
);

AOI21xp5_ASAP7_75t_L g4150 ( 
.A1(n_3921),
.A2(n_3566),
.B(n_3557),
.Y(n_4150)
);

AOI21xp5_ASAP7_75t_L g4151 ( 
.A1(n_3822),
.A2(n_3864),
.B(n_4036),
.Y(n_4151)
);

OR2x2_ASAP7_75t_L g4152 ( 
.A(n_3863),
.B(n_3797),
.Y(n_4152)
);

AOI21xp5_ASAP7_75t_L g4153 ( 
.A1(n_3835),
.A2(n_3557),
.B(n_3527),
.Y(n_4153)
);

A2O1A1Ixp33_ASAP7_75t_L g4154 ( 
.A1(n_3823),
.A2(n_3604),
.B(n_3625),
.C(n_3610),
.Y(n_4154)
);

AO32x1_ASAP7_75t_L g4155 ( 
.A1(n_3814),
.A2(n_3844),
.A3(n_3855),
.B1(n_3879),
.B2(n_3871),
.Y(n_4155)
);

O2A1O1Ixp33_ASAP7_75t_L g4156 ( 
.A1(n_4005),
.A2(n_1602),
.B(n_1603),
.C(n_1599),
.Y(n_4156)
);

NOR2xp33_ASAP7_75t_L g4157 ( 
.A(n_3877),
.B(n_3554),
.Y(n_4157)
);

AOI21xp5_ASAP7_75t_L g4158 ( 
.A1(n_3963),
.A2(n_3797),
.B(n_3569),
.Y(n_4158)
);

NAND2xp5_ASAP7_75t_L g4159 ( 
.A(n_3955),
.B(n_3829),
.Y(n_4159)
);

CKINVDCx6p67_ASAP7_75t_R g4160 ( 
.A(n_3859),
.Y(n_4160)
);

OR2x6_ASAP7_75t_L g4161 ( 
.A(n_3913),
.B(n_3692),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_3894),
.Y(n_4162)
);

AOI21xp5_ASAP7_75t_L g4163 ( 
.A1(n_3963),
.A2(n_3569),
.B(n_3568),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_L g4164 ( 
.A(n_4048),
.B(n_3520),
.Y(n_4164)
);

NOR2xp33_ASAP7_75t_L g4165 ( 
.A(n_4032),
.B(n_3554),
.Y(n_4165)
);

NAND2xp5_ASAP7_75t_L g4166 ( 
.A(n_3839),
.B(n_3533),
.Y(n_4166)
);

OAI22xp5_ASAP7_75t_L g4167 ( 
.A1(n_3922),
.A2(n_4021),
.B1(n_3924),
.B2(n_4024),
.Y(n_4167)
);

AOI21xp5_ASAP7_75t_L g4168 ( 
.A1(n_3802),
.A2(n_3578),
.B(n_3568),
.Y(n_4168)
);

INVx1_ASAP7_75t_L g4169 ( 
.A(n_3910),
.Y(n_4169)
);

BUFx6f_ASAP7_75t_L g4170 ( 
.A(n_3929),
.Y(n_4170)
);

A2O1A1Ixp33_ASAP7_75t_L g4171 ( 
.A1(n_4094),
.A2(n_3752),
.B(n_3723),
.C(n_3751),
.Y(n_4171)
);

AOI21xp5_ASAP7_75t_L g4172 ( 
.A1(n_3802),
.A2(n_3581),
.B(n_3578),
.Y(n_4172)
);

O2A1O1Ixp33_ASAP7_75t_L g4173 ( 
.A1(n_3933),
.A2(n_1607),
.B(n_1609),
.C(n_1606),
.Y(n_4173)
);

BUFx2_ASAP7_75t_SL g4174 ( 
.A(n_3859),
.Y(n_4174)
);

OAI22xp5_ASAP7_75t_L g4175 ( 
.A1(n_3961),
.A2(n_3692),
.B1(n_3505),
.B2(n_3398),
.Y(n_4175)
);

INVx3_ASAP7_75t_L g4176 ( 
.A(n_4078),
.Y(n_4176)
);

BUFx6f_ASAP7_75t_L g4177 ( 
.A(n_3817),
.Y(n_4177)
);

AOI21xp5_ASAP7_75t_L g4178 ( 
.A1(n_4071),
.A2(n_3584),
.B(n_3581),
.Y(n_4178)
);

AOI21xp5_ASAP7_75t_L g4179 ( 
.A1(n_4033),
.A2(n_3586),
.B(n_3584),
.Y(n_4179)
);

NAND2xp5_ASAP7_75t_L g4180 ( 
.A(n_3842),
.B(n_3564),
.Y(n_4180)
);

INVx4_ASAP7_75t_L g4181 ( 
.A(n_4027),
.Y(n_4181)
);

NAND2x1_ASAP7_75t_L g4182 ( 
.A(n_3923),
.B(n_3716),
.Y(n_4182)
);

INVx6_ASAP7_75t_L g4183 ( 
.A(n_4028),
.Y(n_4183)
);

AOI21xp5_ASAP7_75t_L g4184 ( 
.A1(n_4025),
.A2(n_4046),
.B(n_4038),
.Y(n_4184)
);

AOI22xp33_ASAP7_75t_L g4185 ( 
.A1(n_3904),
.A2(n_3574),
.B1(n_3613),
.B2(n_3575),
.Y(n_4185)
);

OAI21x1_ASAP7_75t_L g4186 ( 
.A1(n_3815),
.A2(n_3746),
.B(n_3745),
.Y(n_4186)
);

AOI21xp5_ASAP7_75t_L g4187 ( 
.A1(n_4047),
.A2(n_3596),
.B(n_3586),
.Y(n_4187)
);

AND2x2_ASAP7_75t_L g4188 ( 
.A(n_3999),
.B(n_1610),
.Y(n_4188)
);

AND2x2_ASAP7_75t_L g4189 ( 
.A(n_4008),
.B(n_1611),
.Y(n_4189)
);

AOI21xp5_ASAP7_75t_L g4190 ( 
.A1(n_4057),
.A2(n_3607),
.B(n_3596),
.Y(n_4190)
);

NAND2xp5_ASAP7_75t_L g4191 ( 
.A(n_3850),
.B(n_3614),
.Y(n_4191)
);

OAI22xp5_ASAP7_75t_L g4192 ( 
.A1(n_4080),
.A2(n_3692),
.B1(n_3505),
.B2(n_3398),
.Y(n_4192)
);

A2O1A1Ixp33_ASAP7_75t_L g4193 ( 
.A1(n_4085),
.A2(n_3539),
.B(n_3759),
.C(n_3733),
.Y(n_4193)
);

AND2x2_ASAP7_75t_L g4194 ( 
.A(n_4018),
.B(n_1613),
.Y(n_4194)
);

AND2x2_ASAP7_75t_L g4195 ( 
.A(n_4087),
.B(n_3915),
.Y(n_4195)
);

OAI22xp5_ASAP7_75t_L g4196 ( 
.A1(n_4013),
.A2(n_3732),
.B1(n_3667),
.B2(n_3670),
.Y(n_4196)
);

NOR2xp33_ASAP7_75t_L g4197 ( 
.A(n_4059),
.B(n_963),
.Y(n_4197)
);

O2A1O1Ixp5_ASAP7_75t_L g4198 ( 
.A1(n_3803),
.A2(n_3686),
.B(n_3684),
.C(n_3783),
.Y(n_4198)
);

INVx1_ASAP7_75t_L g4199 ( 
.A(n_3944),
.Y(n_4199)
);

INVx3_ASAP7_75t_L g4200 ( 
.A(n_4078),
.Y(n_4200)
);

NAND2xp5_ASAP7_75t_L g4201 ( 
.A(n_3852),
.B(n_3617),
.Y(n_4201)
);

INVx4_ASAP7_75t_L g4202 ( 
.A(n_4078),
.Y(n_4202)
);

OAI21xp5_ASAP7_75t_L g4203 ( 
.A1(n_3832),
.A2(n_4073),
.B(n_3827),
.Y(n_4203)
);

AND2x2_ASAP7_75t_L g4204 ( 
.A(n_4065),
.B(n_1615),
.Y(n_4204)
);

AND2x2_ASAP7_75t_SL g4205 ( 
.A(n_3824),
.B(n_3693),
.Y(n_4205)
);

BUFx6f_ASAP7_75t_L g4206 ( 
.A(n_3817),
.Y(n_4206)
);

BUFx8_ASAP7_75t_L g4207 ( 
.A(n_3846),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_SL g4208 ( 
.A(n_4011),
.B(n_3670),
.Y(n_4208)
);

NAND3xp33_ASAP7_75t_SL g4209 ( 
.A(n_3867),
.B(n_966),
.C(n_964),
.Y(n_4209)
);

INVx1_ASAP7_75t_L g4210 ( 
.A(n_3947),
.Y(n_4210)
);

AOI22xp33_ASAP7_75t_L g4211 ( 
.A1(n_3920),
.A2(n_3619),
.B1(n_3624),
.B2(n_3618),
.Y(n_4211)
);

NAND2xp5_ASAP7_75t_L g4212 ( 
.A(n_3872),
.B(n_3626),
.Y(n_4212)
);

AOI21xp5_ASAP7_75t_L g4213 ( 
.A1(n_3820),
.A2(n_3607),
.B(n_3746),
.Y(n_4213)
);

O2A1O1Ixp33_ASAP7_75t_L g4214 ( 
.A1(n_3964),
.A2(n_3891),
.B(n_4010),
.C(n_3870),
.Y(n_4214)
);

AND2x4_ASAP7_75t_L g4215 ( 
.A(n_4023),
.B(n_3771),
.Y(n_4215)
);

NOR2xp33_ASAP7_75t_L g4216 ( 
.A(n_4091),
.B(n_969),
.Y(n_4216)
);

OAI22xp5_ASAP7_75t_L g4217 ( 
.A1(n_4023),
.A2(n_3771),
.B1(n_3737),
.B2(n_3735),
.Y(n_4217)
);

NAND2xp5_ASAP7_75t_SL g4218 ( 
.A(n_4011),
.B(n_3785),
.Y(n_4218)
);

NAND2xp5_ASAP7_75t_L g4219 ( 
.A(n_3868),
.B(n_3631),
.Y(n_4219)
);

OAI21xp33_ASAP7_75t_L g4220 ( 
.A1(n_4063),
.A2(n_975),
.B(n_972),
.Y(n_4220)
);

AOI21xp5_ASAP7_75t_L g4221 ( 
.A1(n_3934),
.A2(n_3745),
.B(n_3792),
.Y(n_4221)
);

INVxp33_ASAP7_75t_SL g4222 ( 
.A(n_3974),
.Y(n_4222)
);

INVx1_ASAP7_75t_L g4223 ( 
.A(n_3967),
.Y(n_4223)
);

NAND2xp5_ASAP7_75t_L g4224 ( 
.A(n_3826),
.B(n_3635),
.Y(n_4224)
);

CKINVDCx16_ASAP7_75t_R g4225 ( 
.A(n_3892),
.Y(n_4225)
);

NAND2xp5_ASAP7_75t_L g4226 ( 
.A(n_3806),
.B(n_3646),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_L g4227 ( 
.A(n_3821),
.B(n_3651),
.Y(n_4227)
);

NAND2xp5_ASAP7_75t_SL g4228 ( 
.A(n_3851),
.B(n_3765),
.Y(n_4228)
);

NAND2xp5_ASAP7_75t_L g4229 ( 
.A(n_3897),
.B(n_3895),
.Y(n_4229)
);

NOR2xp33_ASAP7_75t_L g4230 ( 
.A(n_4015),
.B(n_976),
.Y(n_4230)
);

INVxp67_ASAP7_75t_SL g4231 ( 
.A(n_4054),
.Y(n_4231)
);

AOI21xp5_ASAP7_75t_L g4232 ( 
.A1(n_3934),
.A2(n_3773),
.B(n_3765),
.Y(n_4232)
);

INVx1_ASAP7_75t_L g4233 ( 
.A(n_3979),
.Y(n_4233)
);

OAI22x1_ASAP7_75t_L g4234 ( 
.A1(n_3982),
.A2(n_978),
.B1(n_982),
.B2(n_977),
.Y(n_4234)
);

AND2x2_ASAP7_75t_L g4235 ( 
.A(n_3993),
.B(n_1618),
.Y(n_4235)
);

AOI21xp5_ASAP7_75t_L g4236 ( 
.A1(n_3948),
.A2(n_3777),
.B(n_3773),
.Y(n_4236)
);

AOI21xp5_ASAP7_75t_L g4237 ( 
.A1(n_3948),
.A2(n_3779),
.B(n_3777),
.Y(n_4237)
);

OAI21xp5_ASAP7_75t_L g4238 ( 
.A1(n_3827),
.A2(n_1990),
.B(n_3791),
.Y(n_4238)
);

NOR2xp33_ASAP7_75t_L g4239 ( 
.A(n_4028),
.B(n_985),
.Y(n_4239)
);

AOI21xp5_ASAP7_75t_L g4240 ( 
.A1(n_4074),
.A2(n_3793),
.B(n_3792),
.Y(n_4240)
);

AOI22xp5_ASAP7_75t_L g4241 ( 
.A1(n_3856),
.A2(n_3716),
.B1(n_3595),
.B2(n_3402),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_3987),
.Y(n_4242)
);

INVx2_ASAP7_75t_SL g4243 ( 
.A(n_3892),
.Y(n_4243)
);

BUFx6f_ASAP7_75t_L g4244 ( 
.A(n_3892),
.Y(n_4244)
);

OAI22xp5_ASAP7_75t_L g4245 ( 
.A1(n_4017),
.A2(n_3791),
.B1(n_993),
.B2(n_994),
.Y(n_4245)
);

NAND2xp5_ASAP7_75t_L g4246 ( 
.A(n_3936),
.B(n_3654),
.Y(n_4246)
);

NAND2xp5_ASAP7_75t_L g4247 ( 
.A(n_3831),
.B(n_3660),
.Y(n_4247)
);

O2A1O1Ixp33_ASAP7_75t_L g4248 ( 
.A1(n_3940),
.A2(n_1622),
.B(n_1623),
.C(n_1619),
.Y(n_4248)
);

BUFx6f_ASAP7_75t_L g4249 ( 
.A(n_3909),
.Y(n_4249)
);

NAND2xp5_ASAP7_75t_SL g4250 ( 
.A(n_3831),
.B(n_3779),
.Y(n_4250)
);

OAI22xp5_ASAP7_75t_L g4251 ( 
.A1(n_4034),
.A2(n_995),
.B1(n_997),
.B2(n_987),
.Y(n_4251)
);

BUFx3_ASAP7_75t_L g4252 ( 
.A(n_3888),
.Y(n_4252)
);

NAND2xp5_ASAP7_75t_L g4253 ( 
.A(n_3841),
.B(n_3601),
.Y(n_4253)
);

NOR2xp33_ASAP7_75t_L g4254 ( 
.A(n_3841),
.B(n_999),
.Y(n_4254)
);

O2A1O1Ixp33_ASAP7_75t_L g4255 ( 
.A1(n_3981),
.A2(n_1626),
.B(n_1628),
.C(n_1625),
.Y(n_4255)
);

AND2x4_ASAP7_75t_L g4256 ( 
.A(n_3990),
.B(n_3680),
.Y(n_4256)
);

BUFx6f_ASAP7_75t_L g4257 ( 
.A(n_3909),
.Y(n_4257)
);

AOI21xp5_ASAP7_75t_L g4258 ( 
.A1(n_4095),
.A2(n_3794),
.B(n_3793),
.Y(n_4258)
);

NAND2xp5_ASAP7_75t_SL g4259 ( 
.A(n_4089),
.B(n_3794),
.Y(n_4259)
);

NAND2xp5_ASAP7_75t_SL g4260 ( 
.A(n_3978),
.B(n_3796),
.Y(n_4260)
);

NOR2xp33_ASAP7_75t_L g4261 ( 
.A(n_3916),
.B(n_1000),
.Y(n_4261)
);

INVx2_ASAP7_75t_L g4262 ( 
.A(n_3937),
.Y(n_4262)
);

AND2x2_ASAP7_75t_SL g4263 ( 
.A(n_3909),
.B(n_3790),
.Y(n_4263)
);

NAND2xp5_ASAP7_75t_SL g4264 ( 
.A(n_3983),
.B(n_3785),
.Y(n_4264)
);

NAND2xp5_ASAP7_75t_L g4265 ( 
.A(n_3992),
.B(n_3796),
.Y(n_4265)
);

NAND3xp33_ASAP7_75t_L g4266 ( 
.A(n_3935),
.B(n_3874),
.C(n_3996),
.Y(n_4266)
);

AOI22x1_ASAP7_75t_L g4267 ( 
.A1(n_4037),
.A2(n_1004),
.B1(n_1006),
.B2(n_1001),
.Y(n_4267)
);

BUFx6f_ASAP7_75t_L g4268 ( 
.A(n_3975),
.Y(n_4268)
);

NAND2xp5_ASAP7_75t_L g4269 ( 
.A(n_3998),
.B(n_3716),
.Y(n_4269)
);

AOI22xp33_ASAP7_75t_L g4270 ( 
.A1(n_3994),
.A2(n_3595),
.B1(n_3402),
.B2(n_2055),
.Y(n_4270)
);

O2A1O1Ixp33_ASAP7_75t_L g4271 ( 
.A1(n_3860),
.A2(n_4041),
.B(n_4061),
.C(n_4040),
.Y(n_4271)
);

OAI21xp5_ASAP7_75t_L g4272 ( 
.A1(n_3950),
.A2(n_4072),
.B(n_3833),
.Y(n_4272)
);

O2A1O1Ixp33_ASAP7_75t_L g4273 ( 
.A1(n_4068),
.A2(n_1630),
.B(n_1631),
.C(n_1629),
.Y(n_4273)
);

AND2x2_ASAP7_75t_L g4274 ( 
.A(n_4001),
.B(n_1632),
.Y(n_4274)
);

OAI22xp5_ASAP7_75t_L g4275 ( 
.A1(n_4069),
.A2(n_1009),
.B1(n_1010),
.B2(n_1008),
.Y(n_4275)
);

NAND3xp33_ASAP7_75t_L g4276 ( 
.A(n_4006),
.B(n_1013),
.C(n_1011),
.Y(n_4276)
);

AOI21xp5_ASAP7_75t_L g4277 ( 
.A1(n_3919),
.A2(n_3716),
.B(n_2932),
.Y(n_4277)
);

AOI22xp5_ASAP7_75t_L g4278 ( 
.A1(n_3971),
.A2(n_3976),
.B1(n_3925),
.B2(n_3716),
.Y(n_4278)
);

NOR2xp33_ASAP7_75t_L g4279 ( 
.A(n_3975),
.B(n_1015),
.Y(n_4279)
);

NAND2xp5_ASAP7_75t_SL g4280 ( 
.A(n_3990),
.B(n_2297),
.Y(n_4280)
);

AND2x4_ASAP7_75t_L g4281 ( 
.A(n_4067),
.B(n_3402),
.Y(n_4281)
);

INVxp67_ASAP7_75t_L g4282 ( 
.A(n_3912),
.Y(n_4282)
);

INVxp67_ASAP7_75t_SL g4283 ( 
.A(n_3952),
.Y(n_4283)
);

NAND2xp5_ASAP7_75t_L g4284 ( 
.A(n_4035),
.B(n_1633),
.Y(n_4284)
);

NAND2xp5_ASAP7_75t_SL g4285 ( 
.A(n_4067),
.B(n_2297),
.Y(n_4285)
);

AOI22x1_ASAP7_75t_L g4286 ( 
.A1(n_4037),
.A2(n_1019),
.B1(n_1020),
.B2(n_1017),
.Y(n_4286)
);

AOI21x1_ASAP7_75t_L g4287 ( 
.A1(n_4077),
.A2(n_3623),
.B(n_2418),
.Y(n_4287)
);

NAND2xp5_ASAP7_75t_L g4288 ( 
.A(n_3878),
.B(n_1634),
.Y(n_4288)
);

A2O1A1Ixp33_ASAP7_75t_L g4289 ( 
.A1(n_3953),
.A2(n_3959),
.B(n_3956),
.C(n_3984),
.Y(n_4289)
);

NOR2xp33_ASAP7_75t_L g4290 ( 
.A(n_3975),
.B(n_1023),
.Y(n_4290)
);

OR2x2_ASAP7_75t_L g4291 ( 
.A(n_3887),
.B(n_1639),
.Y(n_4291)
);

NAND2xp5_ASAP7_75t_L g4292 ( 
.A(n_3900),
.B(n_1640),
.Y(n_4292)
);

NAND2xp5_ASAP7_75t_L g4293 ( 
.A(n_3907),
.B(n_1641),
.Y(n_4293)
);

AOI21xp5_ASAP7_75t_L g4294 ( 
.A1(n_4022),
.A2(n_3857),
.B(n_3849),
.Y(n_4294)
);

NOR2x1_ASAP7_75t_R g4295 ( 
.A(n_4029),
.B(n_1024),
.Y(n_4295)
);

INVx2_ASAP7_75t_L g4296 ( 
.A(n_3972),
.Y(n_4296)
);

AOI21xp5_ASAP7_75t_L g4297 ( 
.A1(n_3881),
.A2(n_2932),
.B(n_2849),
.Y(n_4297)
);

AOI21xp5_ASAP7_75t_L g4298 ( 
.A1(n_3902),
.A2(n_2932),
.B(n_2849),
.Y(n_4298)
);

O2A1O1Ixp33_ASAP7_75t_L g4299 ( 
.A1(n_4070),
.A2(n_1646),
.B(n_1647),
.C(n_1642),
.Y(n_4299)
);

AOI21xp33_ASAP7_75t_L g4300 ( 
.A1(n_3898),
.A2(n_2301),
.B(n_2297),
.Y(n_4300)
);

AO32x1_ASAP7_75t_L g4301 ( 
.A1(n_3985),
.A2(n_3988),
.A3(n_4056),
.B1(n_3873),
.B2(n_3941),
.Y(n_4301)
);

HB1xp67_ASAP7_75t_L g4302 ( 
.A(n_3926),
.Y(n_4302)
);

AOI21xp5_ASAP7_75t_L g4303 ( 
.A1(n_3836),
.A2(n_4062),
.B(n_3889),
.Y(n_4303)
);

NOR2xp33_ASAP7_75t_L g4304 ( 
.A(n_4029),
.B(n_1026),
.Y(n_4304)
);

NAND2xp5_ASAP7_75t_L g4305 ( 
.A(n_3908),
.B(n_1650),
.Y(n_4305)
);

CKINVDCx5p33_ASAP7_75t_R g4306 ( 
.A(n_4029),
.Y(n_4306)
);

AOI21xp5_ASAP7_75t_L g4307 ( 
.A1(n_3885),
.A2(n_2849),
.B(n_3402),
.Y(n_4307)
);

BUFx6f_ASAP7_75t_L g4308 ( 
.A(n_3923),
.Y(n_4308)
);

NAND2xp5_ASAP7_75t_L g4309 ( 
.A(n_3911),
.B(n_1651),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_4004),
.Y(n_4310)
);

INVx1_ASAP7_75t_L g4311 ( 
.A(n_4030),
.Y(n_4311)
);

NAND2xp5_ASAP7_75t_L g4312 ( 
.A(n_3890),
.B(n_1653),
.Y(n_4312)
);

NAND2xp5_ASAP7_75t_SL g4313 ( 
.A(n_4056),
.B(n_2301),
.Y(n_4313)
);

AOI21xp5_ASAP7_75t_L g4314 ( 
.A1(n_3899),
.A2(n_3595),
.B(n_3322),
.Y(n_4314)
);

AOI21xp5_ASAP7_75t_L g4315 ( 
.A1(n_3901),
.A2(n_3595),
.B(n_2303),
.Y(n_4315)
);

OR2x2_ASAP7_75t_L g4316 ( 
.A(n_3962),
.B(n_1654),
.Y(n_4316)
);

NOR2xp33_ASAP7_75t_L g4317 ( 
.A(n_4096),
.B(n_1027),
.Y(n_4317)
);

AOI21xp5_ASAP7_75t_L g4318 ( 
.A1(n_3905),
.A2(n_3595),
.B(n_2303),
.Y(n_4318)
);

O2A1O1Ixp5_ASAP7_75t_L g4319 ( 
.A1(n_3853),
.A2(n_2420),
.B(n_2421),
.C(n_2413),
.Y(n_4319)
);

AOI22x1_ASAP7_75t_L g4320 ( 
.A1(n_3816),
.A2(n_1029),
.B1(n_1034),
.B2(n_1028),
.Y(n_4320)
);

NAND2xp5_ASAP7_75t_L g4321 ( 
.A(n_3969),
.B(n_1656),
.Y(n_4321)
);

NOR2xp33_ASAP7_75t_L g4322 ( 
.A(n_4093),
.B(n_1035),
.Y(n_4322)
);

OR2x6_ASAP7_75t_SL g4323 ( 
.A(n_4076),
.B(n_1037),
.Y(n_4323)
);

OAI22x1_ASAP7_75t_L g4324 ( 
.A1(n_4003),
.A2(n_4055),
.B1(n_4012),
.B2(n_3896),
.Y(n_4324)
);

NAND2xp5_ASAP7_75t_L g4325 ( 
.A(n_3977),
.B(n_1659),
.Y(n_4325)
);

A2O1A1Ixp33_ASAP7_75t_L g4326 ( 
.A1(n_3984),
.A2(n_1673),
.B(n_1674),
.C(n_1672),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_4049),
.Y(n_4327)
);

NAND2xp5_ASAP7_75t_L g4328 ( 
.A(n_3991),
.B(n_1677),
.Y(n_4328)
);

BUFx6f_ASAP7_75t_L g4329 ( 
.A(n_3951),
.Y(n_4329)
);

BUFx2_ASAP7_75t_SL g4330 ( 
.A(n_3951),
.Y(n_4330)
);

NAND2xp5_ASAP7_75t_SL g4331 ( 
.A(n_3966),
.B(n_2301),
.Y(n_4331)
);

NAND2xp5_ASAP7_75t_L g4332 ( 
.A(n_4014),
.B(n_1678),
.Y(n_4332)
);

AOI22xp5_ASAP7_75t_L g4333 ( 
.A1(n_4081),
.A2(n_1040),
.B1(n_1041),
.B2(n_1038),
.Y(n_4333)
);

AOI21xp5_ASAP7_75t_L g4334 ( 
.A1(n_3927),
.A2(n_2303),
.B(n_2301),
.Y(n_4334)
);

AO21x1_ASAP7_75t_L g4335 ( 
.A1(n_4026),
.A2(n_1701),
.B(n_1684),
.Y(n_4335)
);

INVx2_ASAP7_75t_L g4336 ( 
.A(n_4050),
.Y(n_4336)
);

NAND2xp5_ASAP7_75t_SL g4337 ( 
.A(n_3966),
.B(n_2303),
.Y(n_4337)
);

NOR2xp33_ASAP7_75t_L g4338 ( 
.A(n_4092),
.B(n_1042),
.Y(n_4338)
);

AOI21xp5_ASAP7_75t_L g4339 ( 
.A1(n_3970),
.A2(n_2333),
.B(n_2304),
.Y(n_4339)
);

AOI21xp5_ASAP7_75t_L g4340 ( 
.A1(n_4088),
.A2(n_2333),
.B(n_2304),
.Y(n_4340)
);

AOI21xp5_ASAP7_75t_L g4341 ( 
.A1(n_3882),
.A2(n_2333),
.B(n_2304),
.Y(n_4341)
);

NAND2xp5_ASAP7_75t_L g4342 ( 
.A(n_3939),
.B(n_2045),
.Y(n_4342)
);

NAND2xp5_ASAP7_75t_L g4343 ( 
.A(n_3949),
.B(n_2045),
.Y(n_4343)
);

CKINVDCx5p33_ASAP7_75t_R g4344 ( 
.A(n_4052),
.Y(n_4344)
);

AOI21xp5_ASAP7_75t_L g4345 ( 
.A1(n_3884),
.A2(n_2333),
.B(n_2304),
.Y(n_4345)
);

AOI21xp5_ASAP7_75t_L g4346 ( 
.A1(n_3917),
.A2(n_2352),
.B(n_2346),
.Y(n_4346)
);

NOR2xp67_ASAP7_75t_L g4347 ( 
.A(n_4084),
.B(n_2420),
.Y(n_4347)
);

NAND2xp5_ASAP7_75t_L g4348 ( 
.A(n_4079),
.B(n_2055),
.Y(n_4348)
);

NAND2xp5_ASAP7_75t_L g4349 ( 
.A(n_4082),
.B(n_2055),
.Y(n_4349)
);

OAI22xp5_ASAP7_75t_L g4350 ( 
.A1(n_4090),
.A2(n_1045),
.B1(n_1046),
.B2(n_1044),
.Y(n_4350)
);

INVx2_ASAP7_75t_L g4351 ( 
.A(n_4003),
.Y(n_4351)
);

AOI21x1_ASAP7_75t_L g4352 ( 
.A1(n_3825),
.A2(n_2424),
.B(n_2421),
.Y(n_4352)
);

AOI21xp5_ASAP7_75t_L g4353 ( 
.A1(n_4016),
.A2(n_2352),
.B(n_2346),
.Y(n_4353)
);

OAI22xp5_ASAP7_75t_L g4354 ( 
.A1(n_4045),
.A2(n_4007),
.B1(n_3997),
.B2(n_4051),
.Y(n_4354)
);

A2O1A1Ixp33_ASAP7_75t_L g4355 ( 
.A1(n_3989),
.A2(n_1048),
.B(n_1049),
.C(n_1047),
.Y(n_4355)
);

OAI21xp5_ASAP7_75t_L g4356 ( 
.A1(n_3989),
.A2(n_2438),
.B(n_2424),
.Y(n_4356)
);

AND2x2_ASAP7_75t_SL g4357 ( 
.A(n_3816),
.B(n_2438),
.Y(n_4357)
);

NAND2xp5_ASAP7_75t_L g4358 ( 
.A(n_4000),
.B(n_2055),
.Y(n_4358)
);

NAND2xp5_ASAP7_75t_L g4359 ( 
.A(n_3954),
.B(n_1050),
.Y(n_4359)
);

INVx3_ASAP7_75t_SL g4360 ( 
.A(n_4053),
.Y(n_4360)
);

INVx4_ASAP7_75t_L g4361 ( 
.A(n_3866),
.Y(n_4361)
);

INVx2_ASAP7_75t_L g4362 ( 
.A(n_3980),
.Y(n_4362)
);

NOR2xp33_ASAP7_75t_L g4363 ( 
.A(n_3866),
.B(n_1052),
.Y(n_4363)
);

NOR3xp33_ASAP7_75t_L g4364 ( 
.A(n_3957),
.B(n_1055),
.C(n_1053),
.Y(n_4364)
);

INVx6_ASAP7_75t_L g4365 ( 
.A(n_4058),
.Y(n_4365)
);

NAND2xp5_ASAP7_75t_SL g4366 ( 
.A(n_4002),
.B(n_2346),
.Y(n_4366)
);

NOR2xp67_ASAP7_75t_L g4367 ( 
.A(n_4083),
.B(n_2443),
.Y(n_4367)
);

AO31x2_ASAP7_75t_L g4368 ( 
.A1(n_4303),
.A2(n_3931),
.A3(n_3930),
.B(n_3928),
.Y(n_4368)
);

INVx2_ASAP7_75t_L g4369 ( 
.A(n_4111),
.Y(n_4369)
);

NAND2xp5_ASAP7_75t_L g4370 ( 
.A(n_4195),
.B(n_3965),
.Y(n_4370)
);

NAND2xp5_ASAP7_75t_L g4371 ( 
.A(n_4229),
.B(n_1056),
.Y(n_4371)
);

NAND2xp5_ASAP7_75t_L g4372 ( 
.A(n_4114),
.B(n_1057),
.Y(n_4372)
);

BUFx6f_ASAP7_75t_L g4373 ( 
.A(n_4170),
.Y(n_4373)
);

AO31x2_ASAP7_75t_L g4374 ( 
.A1(n_4362),
.A2(n_3946),
.A3(n_4064),
.B(n_2445),
.Y(n_4374)
);

AOI21xp5_ASAP7_75t_L g4375 ( 
.A1(n_4106),
.A2(n_4044),
.B(n_4019),
.Y(n_4375)
);

BUFx3_ASAP7_75t_L g4376 ( 
.A(n_4146),
.Y(n_4376)
);

AOI21xp33_ASAP7_75t_L g4377 ( 
.A1(n_4271),
.A2(n_4019),
.B(n_4066),
.Y(n_4377)
);

BUFx6f_ASAP7_75t_L g4378 ( 
.A(n_4170),
.Y(n_4378)
);

AO31x2_ASAP7_75t_L g4379 ( 
.A1(n_4099),
.A2(n_2445),
.A3(n_2452),
.B(n_2443),
.Y(n_4379)
);

NAND2xp5_ASAP7_75t_L g4380 ( 
.A(n_4125),
.B(n_1061),
.Y(n_4380)
);

AOI21xp5_ASAP7_75t_L g4381 ( 
.A1(n_4127),
.A2(n_3810),
.B(n_3257),
.Y(n_4381)
);

INVx1_ASAP7_75t_L g4382 ( 
.A(n_4131),
.Y(n_4382)
);

AND2x2_ASAP7_75t_L g4383 ( 
.A(n_4109),
.B(n_7),
.Y(n_4383)
);

AOI21x1_ASAP7_75t_SL g4384 ( 
.A1(n_4204),
.A2(n_7),
.B(n_8),
.Y(n_4384)
);

OAI21x1_ASAP7_75t_L g4385 ( 
.A1(n_4352),
.A2(n_3257),
.B(n_2459),
.Y(n_4385)
);

INVx2_ASAP7_75t_L g4386 ( 
.A(n_4140),
.Y(n_4386)
);

BUFx6f_ASAP7_75t_L g4387 ( 
.A(n_4170),
.Y(n_4387)
);

OA21x2_ASAP7_75t_L g4388 ( 
.A1(n_4151),
.A2(n_4294),
.B(n_4272),
.Y(n_4388)
);

BUFx2_ASAP7_75t_L g4389 ( 
.A(n_4103),
.Y(n_4389)
);

OAI22xp5_ASAP7_75t_L g4390 ( 
.A1(n_4167),
.A2(n_1094),
.B1(n_1110),
.B2(n_1073),
.Y(n_4390)
);

BUFx12f_ASAP7_75t_L g4391 ( 
.A(n_4117),
.Y(n_4391)
);

OAI21x1_ASAP7_75t_L g4392 ( 
.A1(n_4184),
.A2(n_2459),
.B(n_2452),
.Y(n_4392)
);

AND2x2_ASAP7_75t_L g4393 ( 
.A(n_4112),
.B(n_8),
.Y(n_4393)
);

AOI21xp5_ASAP7_75t_L g4394 ( 
.A1(n_4213),
.A2(n_2352),
.B(n_2346),
.Y(n_4394)
);

OAI21xp5_ASAP7_75t_L g4395 ( 
.A1(n_4214),
.A2(n_1101),
.B(n_1078),
.Y(n_4395)
);

AOI21xp5_ASAP7_75t_L g4396 ( 
.A1(n_4153),
.A2(n_2355),
.B(n_2352),
.Y(n_4396)
);

OR2x2_ASAP7_75t_L g4397 ( 
.A(n_4152),
.B(n_9),
.Y(n_4397)
);

NAND3xp33_ASAP7_75t_SL g4398 ( 
.A(n_4104),
.B(n_1085),
.C(n_1063),
.Y(n_4398)
);

INVx3_ASAP7_75t_L g4399 ( 
.A(n_4202),
.Y(n_4399)
);

INVx1_ASAP7_75t_L g4400 ( 
.A(n_4162),
.Y(n_4400)
);

OAI21xp5_ASAP7_75t_L g4401 ( 
.A1(n_4136),
.A2(n_1088),
.B(n_1066),
.Y(n_4401)
);

NAND2xp5_ASAP7_75t_L g4402 ( 
.A(n_4282),
.B(n_1068),
.Y(n_4402)
);

O2A1O1Ixp5_ASAP7_75t_L g4403 ( 
.A1(n_4203),
.A2(n_2466),
.B(n_2479),
.C(n_2463),
.Y(n_4403)
);

OAI21xp5_ASAP7_75t_L g4404 ( 
.A1(n_4116),
.A2(n_1097),
.B(n_1069),
.Y(n_4404)
);

NAND2xp5_ASAP7_75t_SL g4405 ( 
.A(n_4175),
.B(n_2463),
.Y(n_4405)
);

INVx2_ASAP7_75t_L g4406 ( 
.A(n_4145),
.Y(n_4406)
);

OAI21x1_ASAP7_75t_L g4407 ( 
.A1(n_4148),
.A2(n_2479),
.B(n_2466),
.Y(n_4407)
);

OAI22xp5_ASAP7_75t_L g4408 ( 
.A1(n_4355),
.A2(n_1103),
.B1(n_1123),
.B2(n_1070),
.Y(n_4408)
);

OAI21x1_ASAP7_75t_L g4409 ( 
.A1(n_4287),
.A2(n_2496),
.B(n_2484),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4169),
.Y(n_4410)
);

AOI21xp5_ASAP7_75t_L g4411 ( 
.A1(n_4158),
.A2(n_2376),
.B(n_2355),
.Y(n_4411)
);

OAI21xp5_ASAP7_75t_L g4412 ( 
.A1(n_4209),
.A2(n_1108),
.B(n_1072),
.Y(n_4412)
);

AOI221x1_ASAP7_75t_L g4413 ( 
.A1(n_4138),
.A2(n_1775),
.B1(n_1788),
.B2(n_1771),
.C(n_1770),
.Y(n_4413)
);

OAI21x1_ASAP7_75t_L g4414 ( 
.A1(n_4340),
.A2(n_4277),
.B(n_4353),
.Y(n_4414)
);

BUFx6f_ASAP7_75t_L g4415 ( 
.A(n_4263),
.Y(n_4415)
);

AOI21xp5_ASAP7_75t_L g4416 ( 
.A1(n_4179),
.A2(n_4101),
.B(n_4187),
.Y(n_4416)
);

OAI21x1_ASAP7_75t_L g4417 ( 
.A1(n_4341),
.A2(n_2496),
.B(n_2484),
.Y(n_4417)
);

OAI21x1_ASAP7_75t_L g4418 ( 
.A1(n_4345),
.A2(n_2376),
.B(n_2355),
.Y(n_4418)
);

NAND2xp5_ASAP7_75t_L g4419 ( 
.A(n_4139),
.B(n_1076),
.Y(n_4419)
);

INVx2_ASAP7_75t_L g4420 ( 
.A(n_4262),
.Y(n_4420)
);

INVx2_ASAP7_75t_L g4421 ( 
.A(n_4296),
.Y(n_4421)
);

OAI21xp5_ASAP7_75t_L g4422 ( 
.A1(n_4317),
.A2(n_1120),
.B(n_1079),
.Y(n_4422)
);

BUFx4_ASAP7_75t_SL g4423 ( 
.A(n_4252),
.Y(n_4423)
);

AND2x2_ASAP7_75t_L g4424 ( 
.A(n_4097),
.B(n_11),
.Y(n_4424)
);

AO31x2_ASAP7_75t_L g4425 ( 
.A1(n_4141),
.A2(n_4240),
.A3(n_4258),
.B(n_4178),
.Y(n_4425)
);

NOR2xp33_ASAP7_75t_L g4426 ( 
.A(n_4323),
.B(n_1086),
.Y(n_4426)
);

NAND2xp5_ASAP7_75t_L g4427 ( 
.A(n_4133),
.B(n_1091),
.Y(n_4427)
);

OA21x2_ASAP7_75t_L g4428 ( 
.A1(n_4366),
.A2(n_1102),
.B(n_1095),
.Y(n_4428)
);

AOI21x1_ASAP7_75t_L g4429 ( 
.A1(n_4324),
.A2(n_1798),
.B(n_1756),
.Y(n_4429)
);

NOR2xp33_ASAP7_75t_L g4430 ( 
.A(n_4121),
.B(n_1104),
.Y(n_4430)
);

OAI221xp5_ASAP7_75t_L g4431 ( 
.A1(n_4322),
.A2(n_1121),
.B1(n_1122),
.B2(n_1117),
.C(n_1112),
.Y(n_4431)
);

INVx1_ASAP7_75t_L g4432 ( 
.A(n_4199),
.Y(n_4432)
);

INVxp67_ASAP7_75t_L g4433 ( 
.A(n_4130),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_L g4434 ( 
.A(n_4283),
.B(n_1129),
.Y(n_4434)
);

BUFx3_ASAP7_75t_L g4435 ( 
.A(n_4183),
.Y(n_4435)
);

NAND2xp5_ASAP7_75t_L g4436 ( 
.A(n_4147),
.B(n_1130),
.Y(n_4436)
);

NAND2xp5_ASAP7_75t_L g4437 ( 
.A(n_4159),
.B(n_1135),
.Y(n_4437)
);

INVx1_ASAP7_75t_L g4438 ( 
.A(n_4210),
.Y(n_4438)
);

NAND2xp5_ASAP7_75t_L g4439 ( 
.A(n_4098),
.B(n_1136),
.Y(n_4439)
);

NAND2xp5_ASAP7_75t_L g4440 ( 
.A(n_4302),
.B(n_1143),
.Y(n_4440)
);

AND2x2_ASAP7_75t_L g4441 ( 
.A(n_4205),
.B(n_11),
.Y(n_4441)
);

NAND2xp5_ASAP7_75t_L g4442 ( 
.A(n_4224),
.B(n_4226),
.Y(n_4442)
);

OAI21xp5_ASAP7_75t_L g4443 ( 
.A1(n_4338),
.A2(n_4354),
.B(n_4198),
.Y(n_4443)
);

NAND2xp5_ASAP7_75t_L g4444 ( 
.A(n_4227),
.B(n_4265),
.Y(n_4444)
);

NOR2xp33_ASAP7_75t_L g4445 ( 
.A(n_4222),
.B(n_1146),
.Y(n_4445)
);

OAI22xp5_ASAP7_75t_L g4446 ( 
.A1(n_4276),
.A2(n_1151),
.B1(n_1194),
.B2(n_1171),
.Y(n_4446)
);

AO31x2_ASAP7_75t_L g4447 ( 
.A1(n_4217),
.A2(n_2853),
.A3(n_2865),
.B(n_2506),
.Y(n_4447)
);

OAI21x1_ASAP7_75t_L g4448 ( 
.A1(n_4346),
.A2(n_2376),
.B(n_2355),
.Y(n_4448)
);

AOI21xp5_ASAP7_75t_L g4449 ( 
.A1(n_4190),
.A2(n_2379),
.B(n_2376),
.Y(n_4449)
);

INVx1_ASAP7_75t_L g4450 ( 
.A(n_4223),
.Y(n_4450)
);

OAI21x1_ASAP7_75t_L g4451 ( 
.A1(n_4334),
.A2(n_4314),
.B(n_4339),
.Y(n_4451)
);

OAI21x1_ASAP7_75t_L g4452 ( 
.A1(n_4318),
.A2(n_2384),
.B(n_2379),
.Y(n_4452)
);

NAND2xp5_ASAP7_75t_L g4453 ( 
.A(n_4231),
.B(n_1147),
.Y(n_4453)
);

INVx2_ASAP7_75t_L g4454 ( 
.A(n_4336),
.Y(n_4454)
);

OAI21x1_ASAP7_75t_L g4455 ( 
.A1(n_4315),
.A2(n_4307),
.B(n_4105),
.Y(n_4455)
);

OAI21xp5_ASAP7_75t_L g4456 ( 
.A1(n_4115),
.A2(n_1179),
.B(n_1158),
.Y(n_4456)
);

INVxp67_ASAP7_75t_L g4457 ( 
.A(n_4188),
.Y(n_4457)
);

BUFx6f_ASAP7_75t_L g4458 ( 
.A(n_4177),
.Y(n_4458)
);

BUFx6f_ASAP7_75t_L g4459 ( 
.A(n_4177),
.Y(n_4459)
);

OAI21x1_ASAP7_75t_L g4460 ( 
.A1(n_4186),
.A2(n_2384),
.B(n_2379),
.Y(n_4460)
);

OAI21x1_ASAP7_75t_L g4461 ( 
.A1(n_4120),
.A2(n_2384),
.B(n_2379),
.Y(n_4461)
);

NAND2xp5_ASAP7_75t_L g4462 ( 
.A(n_4233),
.B(n_4242),
.Y(n_4462)
);

AOI221x1_ASAP7_75t_L g4463 ( 
.A1(n_4137),
.A2(n_1788),
.B1(n_1795),
.B2(n_1775),
.C(n_1771),
.Y(n_4463)
);

OR2x2_ASAP7_75t_L g4464 ( 
.A(n_4123),
.B(n_12),
.Y(n_4464)
);

NAND2xp5_ASAP7_75t_L g4465 ( 
.A(n_4189),
.B(n_1156),
.Y(n_4465)
);

CKINVDCx16_ASAP7_75t_R g4466 ( 
.A(n_4108),
.Y(n_4466)
);

OAI21x1_ASAP7_75t_L g4467 ( 
.A1(n_4168),
.A2(n_2394),
.B(n_2384),
.Y(n_4467)
);

NAND2xp5_ASAP7_75t_L g4468 ( 
.A(n_4194),
.B(n_1162),
.Y(n_4468)
);

OAI21x1_ASAP7_75t_L g4469 ( 
.A1(n_4172),
.A2(n_2409),
.B(n_2394),
.Y(n_4469)
);

INVx1_ASAP7_75t_L g4470 ( 
.A(n_4269),
.Y(n_4470)
);

AOI211x1_ASAP7_75t_L g4471 ( 
.A1(n_4124),
.A2(n_14),
.B(n_12),
.C(n_13),
.Y(n_4471)
);

AOI21xp5_ASAP7_75t_L g4472 ( 
.A1(n_4163),
.A2(n_2409),
.B(n_2394),
.Y(n_4472)
);

A2O1A1Ixp33_ASAP7_75t_L g4473 ( 
.A1(n_4261),
.A2(n_1168),
.B(n_1169),
.C(n_1166),
.Y(n_4473)
);

OAI21x1_ASAP7_75t_L g4474 ( 
.A1(n_4298),
.A2(n_2409),
.B(n_2394),
.Y(n_4474)
);

OAI21x1_ASAP7_75t_L g4475 ( 
.A1(n_4297),
.A2(n_2410),
.B(n_2409),
.Y(n_4475)
);

NAND2xp5_ASAP7_75t_L g4476 ( 
.A(n_4289),
.B(n_1170),
.Y(n_4476)
);

O2A1O1Ixp33_ASAP7_75t_L g4477 ( 
.A1(n_4100),
.A2(n_1177),
.B(n_1182),
.C(n_1175),
.Y(n_4477)
);

AO22x2_ASAP7_75t_L g4478 ( 
.A1(n_4218),
.A2(n_1822),
.B1(n_1826),
.B2(n_1756),
.Y(n_4478)
);

INVx1_ASAP7_75t_L g4479 ( 
.A(n_4301),
.Y(n_4479)
);

AO31x2_ASAP7_75t_L g4480 ( 
.A1(n_4232),
.A2(n_2853),
.A3(n_2865),
.B(n_1826),
.Y(n_4480)
);

NAND2xp5_ASAP7_75t_L g4481 ( 
.A(n_4149),
.B(n_1184),
.Y(n_4481)
);

OAI21x1_ASAP7_75t_L g4482 ( 
.A1(n_4260),
.A2(n_2410),
.B(n_1890),
.Y(n_4482)
);

NOR2xp33_ASAP7_75t_L g4483 ( 
.A(n_4239),
.B(n_1190),
.Y(n_4483)
);

OA21x2_ASAP7_75t_L g4484 ( 
.A1(n_4142),
.A2(n_4118),
.B(n_4264),
.Y(n_4484)
);

AO31x2_ASAP7_75t_L g4485 ( 
.A1(n_4236),
.A2(n_2865),
.A3(n_2853),
.B(n_2336),
.Y(n_4485)
);

OAI21x1_ASAP7_75t_L g4486 ( 
.A1(n_4237),
.A2(n_2410),
.B(n_1890),
.Y(n_4486)
);

OAI22xp5_ASAP7_75t_L g4487 ( 
.A1(n_4171),
.A2(n_1222),
.B1(n_1243),
.B2(n_1203),
.Y(n_4487)
);

OA22x2_ASAP7_75t_L g4488 ( 
.A1(n_4122),
.A2(n_4278),
.B1(n_4208),
.B2(n_4128),
.Y(n_4488)
);

INVx1_ASAP7_75t_L g4489 ( 
.A(n_4301),
.Y(n_4489)
);

AND2x2_ASAP7_75t_L g4490 ( 
.A(n_4225),
.B(n_14),
.Y(n_4490)
);

NAND2xp5_ASAP7_75t_L g4491 ( 
.A(n_4166),
.B(n_1191),
.Y(n_4491)
);

OR2x6_ASAP7_75t_L g4492 ( 
.A(n_4183),
.B(n_2410),
.Y(n_4492)
);

INVx2_ASAP7_75t_L g4493 ( 
.A(n_4310),
.Y(n_4493)
);

CKINVDCx11_ASAP7_75t_R g4494 ( 
.A(n_4110),
.Y(n_4494)
);

INVx3_ASAP7_75t_L g4495 ( 
.A(n_4202),
.Y(n_4495)
);

OAI21xp5_ASAP7_75t_L g4496 ( 
.A1(n_4193),
.A2(n_1232),
.B(n_1210),
.Y(n_4496)
);

AND2x2_ASAP7_75t_L g4497 ( 
.A(n_4274),
.B(n_15),
.Y(n_4497)
);

OAI21x1_ASAP7_75t_L g4498 ( 
.A1(n_4358),
.A2(n_1890),
.B(n_2431),
.Y(n_4498)
);

NAND3xp33_ASAP7_75t_SL g4499 ( 
.A(n_4333),
.B(n_1241),
.C(n_1213),
.Y(n_4499)
);

OAI21xp5_ASAP7_75t_L g4500 ( 
.A1(n_4364),
.A2(n_1247),
.B(n_1218),
.Y(n_4500)
);

AO22x1_ASAP7_75t_L g4501 ( 
.A1(n_4157),
.A2(n_1202),
.B1(n_1207),
.B2(n_1195),
.Y(n_4501)
);

AND2x4_ASAP7_75t_L g4502 ( 
.A(n_4161),
.B(n_2431),
.Y(n_4502)
);

INVx1_ASAP7_75t_L g4503 ( 
.A(n_4301),
.Y(n_4503)
);

OAI21x1_ASAP7_75t_L g4504 ( 
.A1(n_4221),
.A2(n_2435),
.B(n_2431),
.Y(n_4504)
);

AOI21xp5_ASAP7_75t_L g4505 ( 
.A1(n_4143),
.A2(n_2435),
.B(n_2431),
.Y(n_4505)
);

BUFx8_ASAP7_75t_SL g4506 ( 
.A(n_4306),
.Y(n_4506)
);

AOI21xp33_ASAP7_75t_L g4507 ( 
.A1(n_4107),
.A2(n_2426),
.B(n_1211),
.Y(n_4507)
);

AOI21xp5_ASAP7_75t_L g4508 ( 
.A1(n_4150),
.A2(n_2450),
.B(n_2435),
.Y(n_4508)
);

OAI21x1_ASAP7_75t_L g4509 ( 
.A1(n_4319),
.A2(n_2450),
.B(n_2435),
.Y(n_4509)
);

NAND2xp5_ASAP7_75t_L g4510 ( 
.A(n_4180),
.B(n_1209),
.Y(n_4510)
);

OAI21x1_ASAP7_75t_L g4511 ( 
.A1(n_4238),
.A2(n_2457),
.B(n_2450),
.Y(n_4511)
);

AND2x2_ASAP7_75t_L g4512 ( 
.A(n_4235),
.B(n_4176),
.Y(n_4512)
);

INVx1_ASAP7_75t_L g4513 ( 
.A(n_4351),
.Y(n_4513)
);

OAI21x1_ASAP7_75t_L g4514 ( 
.A1(n_4182),
.A2(n_2457),
.B(n_2450),
.Y(n_4514)
);

INVx1_ASAP7_75t_L g4515 ( 
.A(n_4311),
.Y(n_4515)
);

A2O1A1Ixp33_ASAP7_75t_L g4516 ( 
.A1(n_4220),
.A2(n_1223),
.B(n_1225),
.C(n_1219),
.Y(n_4516)
);

OAI21x1_ASAP7_75t_L g4517 ( 
.A1(n_4356),
.A2(n_4102),
.B(n_4259),
.Y(n_4517)
);

AND2x2_ASAP7_75t_L g4518 ( 
.A(n_4176),
.B(n_16),
.Y(n_4518)
);

AND2x4_ASAP7_75t_SL g4519 ( 
.A(n_4181),
.B(n_2457),
.Y(n_4519)
);

OAI21xp33_ASAP7_75t_L g4520 ( 
.A1(n_4251),
.A2(n_1233),
.B(n_1229),
.Y(n_4520)
);

INVx2_ASAP7_75t_L g4521 ( 
.A(n_4327),
.Y(n_4521)
);

BUFx6f_ASAP7_75t_L g4522 ( 
.A(n_4177),
.Y(n_4522)
);

INVx1_ASAP7_75t_SL g4523 ( 
.A(n_4174),
.Y(n_4523)
);

OA22x2_ASAP7_75t_L g4524 ( 
.A1(n_4161),
.A2(n_1246),
.B1(n_1251),
.B2(n_1238),
.Y(n_4524)
);

A2O1A1Ixp33_ASAP7_75t_L g4525 ( 
.A1(n_4347),
.A2(n_1256),
.B(n_1257),
.C(n_1252),
.Y(n_4525)
);

OAI21x1_ASAP7_75t_L g4526 ( 
.A1(n_4228),
.A2(n_2471),
.B(n_2457),
.Y(n_4526)
);

OAI22xp5_ASAP7_75t_L g4527 ( 
.A1(n_4245),
.A2(n_1259),
.B1(n_1260),
.B2(n_1258),
.Y(n_4527)
);

OAI21x1_ASAP7_75t_L g4528 ( 
.A1(n_4132),
.A2(n_2475),
.B(n_2471),
.Y(n_4528)
);

OAI21x1_ASAP7_75t_L g4529 ( 
.A1(n_4348),
.A2(n_2475),
.B(n_2471),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_L g4530 ( 
.A(n_4191),
.B(n_17),
.Y(n_4530)
);

NOR2x1_ASAP7_75t_R g4531 ( 
.A(n_4181),
.B(n_2426),
.Y(n_4531)
);

AO21x2_ASAP7_75t_L g4532 ( 
.A1(n_4300),
.A2(n_2243),
.B(n_2426),
.Y(n_4532)
);

AOI21xp5_ASAP7_75t_L g4533 ( 
.A1(n_4155),
.A2(n_2475),
.B(n_2471),
.Y(n_4533)
);

AOI21xp5_ASAP7_75t_SL g4534 ( 
.A1(n_4154),
.A2(n_2481),
.B(n_2426),
.Y(n_4534)
);

BUFx6f_ASAP7_75t_L g4535 ( 
.A(n_4206),
.Y(n_4535)
);

OAI21x1_ASAP7_75t_L g4536 ( 
.A1(n_4349),
.A2(n_2476),
.B(n_2475),
.Y(n_4536)
);

AND3x2_ASAP7_75t_L g4537 ( 
.A(n_4165),
.B(n_21),
.C(n_19),
.Y(n_4537)
);

OAI21x1_ASAP7_75t_L g4538 ( 
.A1(n_4250),
.A2(n_2493),
.B(n_2476),
.Y(n_4538)
);

AOI21xp5_ASAP7_75t_L g4539 ( 
.A1(n_4155),
.A2(n_2493),
.B(n_2476),
.Y(n_4539)
);

OAI21x1_ASAP7_75t_L g4540 ( 
.A1(n_4196),
.A2(n_2493),
.B(n_2476),
.Y(n_4540)
);

AOI21xp5_ASAP7_75t_L g4541 ( 
.A1(n_4331),
.A2(n_2493),
.B(n_2243),
.Y(n_4541)
);

NAND2x1p5_ASAP7_75t_L g4542 ( 
.A(n_4113),
.B(n_2243),
.Y(n_4542)
);

HB1xp67_ASAP7_75t_L g4543 ( 
.A(n_4253),
.Y(n_4543)
);

INVx2_ASAP7_75t_L g4544 ( 
.A(n_4246),
.Y(n_4544)
);

AOI21xp5_ASAP7_75t_L g4545 ( 
.A1(n_4337),
.A2(n_2353),
.B(n_2336),
.Y(n_4545)
);

INVx1_ASAP7_75t_L g4546 ( 
.A(n_4201),
.Y(n_4546)
);

OAI21x1_ASAP7_75t_SL g4547 ( 
.A1(n_4192),
.A2(n_18),
.B(n_22),
.Y(n_4547)
);

NAND2xp5_ASAP7_75t_L g4548 ( 
.A(n_4219),
.B(n_22),
.Y(n_4548)
);

AND2x2_ASAP7_75t_L g4549 ( 
.A(n_4200),
.B(n_23),
.Y(n_4549)
);

AOI21x1_ASAP7_75t_SL g4550 ( 
.A1(n_4359),
.A2(n_23),
.B(n_25),
.Y(n_4550)
);

O2A1O1Ixp5_ASAP7_75t_L g4551 ( 
.A1(n_4335),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_4551)
);

INVx3_ASAP7_75t_L g4552 ( 
.A(n_4365),
.Y(n_4552)
);

NAND3xp33_ASAP7_75t_SL g4553 ( 
.A(n_4230),
.B(n_26),
.C(n_27),
.Y(n_4553)
);

A2O1A1Ixp33_ASAP7_75t_L g4554 ( 
.A1(n_4363),
.A2(n_2481),
.B(n_30),
.C(n_28),
.Y(n_4554)
);

NAND2xp5_ASAP7_75t_L g4555 ( 
.A(n_4164),
.B(n_29),
.Y(n_4555)
);

OAI21x1_ASAP7_75t_L g4556 ( 
.A1(n_4342),
.A2(n_1775),
.B(n_1771),
.Y(n_4556)
);

OAI21x1_ASAP7_75t_L g4557 ( 
.A1(n_4343),
.A2(n_1775),
.B(n_1771),
.Y(n_4557)
);

OAI21x1_ASAP7_75t_L g4558 ( 
.A1(n_4270),
.A2(n_1795),
.B(n_1788),
.Y(n_4558)
);

NAND2xp5_ASAP7_75t_SL g4559 ( 
.A(n_4308),
.B(n_1788),
.Y(n_4559)
);

NAND2xp5_ASAP7_75t_L g4560 ( 
.A(n_4212),
.B(n_30),
.Y(n_4560)
);

BUFx6f_ASAP7_75t_L g4561 ( 
.A(n_4206),
.Y(n_4561)
);

INVx1_ASAP7_75t_L g4562 ( 
.A(n_4247),
.Y(n_4562)
);

OAI21x1_ASAP7_75t_L g4563 ( 
.A1(n_4241),
.A2(n_1800),
.B(n_1795),
.Y(n_4563)
);

NAND2xp5_ASAP7_75t_SL g4564 ( 
.A(n_4308),
.B(n_1795),
.Y(n_4564)
);

AOI21xp5_ASAP7_75t_L g4565 ( 
.A1(n_4313),
.A2(n_2336),
.B(n_2353),
.Y(n_4565)
);

OAI21xp5_ASAP7_75t_L g4566 ( 
.A1(n_4254),
.A2(n_1724),
.B(n_1723),
.Y(n_4566)
);

NOR2x1_ASAP7_75t_L g4567 ( 
.A(n_4266),
.B(n_1800),
.Y(n_4567)
);

OAI21x1_ASAP7_75t_L g4568 ( 
.A1(n_4280),
.A2(n_1812),
.B(n_1800),
.Y(n_4568)
);

OAI21xp5_ASAP7_75t_L g4569 ( 
.A1(n_4197),
.A2(n_1724),
.B(n_1723),
.Y(n_4569)
);

BUFx10_ASAP7_75t_L g4570 ( 
.A(n_4279),
.Y(n_4570)
);

NOR2xp33_ASAP7_75t_L g4571 ( 
.A(n_4144),
.B(n_31),
.Y(n_4571)
);

AOI21xp5_ASAP7_75t_L g4572 ( 
.A1(n_4357),
.A2(n_4285),
.B(n_4215),
.Y(n_4572)
);

OAI21x1_ASAP7_75t_L g4573 ( 
.A1(n_4200),
.A2(n_4367),
.B(n_4211),
.Y(n_4573)
);

NOR2xp67_ASAP7_75t_SL g4574 ( 
.A(n_4113),
.B(n_4330),
.Y(n_4574)
);

NAND2xp5_ASAP7_75t_L g4575 ( 
.A(n_4291),
.B(n_32),
.Y(n_4575)
);

AO31x2_ASAP7_75t_L g4576 ( 
.A1(n_4126),
.A2(n_2353),
.A3(n_1871),
.B(n_1875),
.Y(n_4576)
);

OAI21x1_ASAP7_75t_L g4577 ( 
.A1(n_4284),
.A2(n_1812),
.B(n_1800),
.Y(n_4577)
);

AOI21xp5_ASAP7_75t_L g4578 ( 
.A1(n_4215),
.A2(n_2015),
.B(n_1813),
.Y(n_4578)
);

BUFx2_ASAP7_75t_L g4579 ( 
.A(n_4206),
.Y(n_4579)
);

AND2x2_ASAP7_75t_L g4580 ( 
.A(n_4129),
.B(n_33),
.Y(n_4580)
);

NAND2x1p5_ASAP7_75t_L g4581 ( 
.A(n_4244),
.B(n_1812),
.Y(n_4581)
);

OAI21x1_ASAP7_75t_SL g4582 ( 
.A1(n_4320),
.A2(n_33),
.B(n_34),
.Y(n_4582)
);

AOI21xp5_ASAP7_75t_L g4583 ( 
.A1(n_4281),
.A2(n_2015),
.B(n_1813),
.Y(n_4583)
);

OAI21x1_ASAP7_75t_SL g4584 ( 
.A1(n_4243),
.A2(n_35),
.B(n_36),
.Y(n_4584)
);

INVx2_ASAP7_75t_L g4585 ( 
.A(n_4344),
.Y(n_4585)
);

NAND2xp5_ASAP7_75t_L g4586 ( 
.A(n_4288),
.B(n_35),
.Y(n_4586)
);

OAI21xp5_ASAP7_75t_SL g4587 ( 
.A1(n_4290),
.A2(n_36),
.B(n_37),
.Y(n_4587)
);

OAI21x1_ASAP7_75t_L g4588 ( 
.A1(n_4292),
.A2(n_1813),
.B(n_1812),
.Y(n_4588)
);

NAND2xp5_ASAP7_75t_L g4589 ( 
.A(n_4316),
.B(n_37),
.Y(n_4589)
);

OA21x2_ASAP7_75t_L g4590 ( 
.A1(n_4326),
.A2(n_1843),
.B(n_1813),
.Y(n_4590)
);

INVx2_ASAP7_75t_L g4591 ( 
.A(n_4256),
.Y(n_4591)
);

HB1xp67_ASAP7_75t_L g4592 ( 
.A(n_4365),
.Y(n_4592)
);

AOI22xp5_ASAP7_75t_L g4593 ( 
.A1(n_4234),
.A2(n_1854),
.B1(n_1855),
.B2(n_1843),
.Y(n_4593)
);

OR2x6_ASAP7_75t_L g4594 ( 
.A(n_4135),
.B(n_1843),
.Y(n_4594)
);

INVx2_ASAP7_75t_SL g4595 ( 
.A(n_4135),
.Y(n_4595)
);

NAND2xp5_ASAP7_75t_L g4596 ( 
.A(n_4312),
.B(n_38),
.Y(n_4596)
);

OAI21x1_ASAP7_75t_L g4597 ( 
.A1(n_4293),
.A2(n_1854),
.B(n_1843),
.Y(n_4597)
);

OR2x2_ASAP7_75t_L g4598 ( 
.A(n_4321),
.B(n_38),
.Y(n_4598)
);

AO31x2_ASAP7_75t_L g4599 ( 
.A1(n_4361),
.A2(n_1871),
.A3(n_1875),
.B(n_1868),
.Y(n_4599)
);

OAI21xp5_ASAP7_75t_L g4600 ( 
.A1(n_4216),
.A2(n_1724),
.B(n_1723),
.Y(n_4600)
);

BUFx3_ASAP7_75t_L g4601 ( 
.A(n_4207),
.Y(n_4601)
);

AND2x2_ASAP7_75t_L g4602 ( 
.A(n_4244),
.B(n_39),
.Y(n_4602)
);

NAND2xp5_ASAP7_75t_L g4603 ( 
.A(n_4305),
.B(n_40),
.Y(n_4603)
);

AOI22xp33_ASAP7_75t_L g4604 ( 
.A1(n_4185),
.A2(n_1855),
.B1(n_1861),
.B2(n_1854),
.Y(n_4604)
);

AND2x2_ASAP7_75t_L g4605 ( 
.A(n_4244),
.B(n_4249),
.Y(n_4605)
);

A2O1A1Ixp33_ASAP7_75t_L g4606 ( 
.A1(n_4273),
.A2(n_42),
.B(n_40),
.C(n_41),
.Y(n_4606)
);

OAI21x1_ASAP7_75t_L g4607 ( 
.A1(n_4309),
.A2(n_1855),
.B(n_1854),
.Y(n_4607)
);

OAI21xp5_ASAP7_75t_L g4608 ( 
.A1(n_4275),
.A2(n_1724),
.B(n_1723),
.Y(n_4608)
);

NAND3xp33_ASAP7_75t_SL g4609 ( 
.A(n_4304),
.B(n_41),
.C(n_42),
.Y(n_4609)
);

OAI21x1_ASAP7_75t_L g4610 ( 
.A1(n_4325),
.A2(n_1861),
.B(n_1855),
.Y(n_4610)
);

AOI21x1_ASAP7_75t_SL g4611 ( 
.A1(n_4160),
.A2(n_45),
.B(n_46),
.Y(n_4611)
);

CKINVDCx5p33_ASAP7_75t_R g4612 ( 
.A(n_4207),
.Y(n_4612)
);

INVx1_ASAP7_75t_L g4613 ( 
.A(n_4328),
.Y(n_4613)
);

AOI21xp5_ASAP7_75t_L g4614 ( 
.A1(n_4281),
.A2(n_2015),
.B(n_1865),
.Y(n_4614)
);

OR2x2_ASAP7_75t_L g4615 ( 
.A(n_4332),
.B(n_47),
.Y(n_4615)
);

NAND2xp5_ASAP7_75t_L g4616 ( 
.A(n_4256),
.B(n_48),
.Y(n_4616)
);

BUFx6f_ASAP7_75t_L g4617 ( 
.A(n_4249),
.Y(n_4617)
);

AO21x1_ASAP7_75t_L g4618 ( 
.A1(n_4350),
.A2(n_50),
.B(n_51),
.Y(n_4618)
);

NAND2xp5_ASAP7_75t_SL g4619 ( 
.A(n_4308),
.B(n_1861),
.Y(n_4619)
);

NAND2xp5_ASAP7_75t_SL g4620 ( 
.A(n_4329),
.B(n_1861),
.Y(n_4620)
);

AOI21x1_ASAP7_75t_L g4621 ( 
.A1(n_4119),
.A2(n_1865),
.B(n_1753),
.Y(n_4621)
);

CKINVDCx5p33_ASAP7_75t_R g4622 ( 
.A(n_4134),
.Y(n_4622)
);

AOI21xp5_ASAP7_75t_L g4623 ( 
.A1(n_4119),
.A2(n_2015),
.B(n_1865),
.Y(n_4623)
);

BUFx2_ASAP7_75t_L g4624 ( 
.A(n_4249),
.Y(n_4624)
);

BUFx3_ASAP7_75t_L g4625 ( 
.A(n_4134),
.Y(n_4625)
);

OAI21x1_ASAP7_75t_L g4626 ( 
.A1(n_4248),
.A2(n_1865),
.B(n_1753),
.Y(n_4626)
);

NAND2xp5_ASAP7_75t_SL g4627 ( 
.A(n_4443),
.B(n_4257),
.Y(n_4627)
);

BUFx6f_ASAP7_75t_L g4628 ( 
.A(n_4415),
.Y(n_4628)
);

OR2x2_ASAP7_75t_L g4629 ( 
.A(n_4389),
.B(n_4360),
.Y(n_4629)
);

OR2x2_ASAP7_75t_L g4630 ( 
.A(n_4543),
.B(n_4257),
.Y(n_4630)
);

INVx2_ASAP7_75t_SL g4631 ( 
.A(n_4376),
.Y(n_4631)
);

INVx1_ASAP7_75t_L g4632 ( 
.A(n_4400),
.Y(n_4632)
);

AOI21xp5_ASAP7_75t_L g4633 ( 
.A1(n_4416),
.A2(n_4329),
.B(n_4361),
.Y(n_4633)
);

OAI22xp5_ASAP7_75t_L g4634 ( 
.A1(n_4587),
.A2(n_4329),
.B1(n_4257),
.B2(n_4268),
.Y(n_4634)
);

OR2x6_ASAP7_75t_L g4635 ( 
.A(n_4488),
.B(n_4268),
.Y(n_4635)
);

OAI22xp5_ASAP7_75t_L g4636 ( 
.A1(n_4390),
.A2(n_4268),
.B1(n_4267),
.B2(n_4286),
.Y(n_4636)
);

AND2x4_ASAP7_75t_L g4637 ( 
.A(n_4591),
.B(n_50),
.Y(n_4637)
);

NAND2xp5_ASAP7_75t_L g4638 ( 
.A(n_4444),
.B(n_4295),
.Y(n_4638)
);

AOI21xp5_ASAP7_75t_L g4639 ( 
.A1(n_4608),
.A2(n_4388),
.B(n_4375),
.Y(n_4639)
);

AND2x2_ASAP7_75t_L g4640 ( 
.A(n_4512),
.B(n_51),
.Y(n_4640)
);

OR2x6_ASAP7_75t_L g4641 ( 
.A(n_4534),
.B(n_4299),
.Y(n_4641)
);

INVx1_ASAP7_75t_L g4642 ( 
.A(n_4400),
.Y(n_4642)
);

HB1xp67_ASAP7_75t_L g4643 ( 
.A(n_4370),
.Y(n_4643)
);

NAND2xp5_ASAP7_75t_SL g4644 ( 
.A(n_4552),
.B(n_4156),
.Y(n_4644)
);

BUFx6f_ASAP7_75t_L g4645 ( 
.A(n_4415),
.Y(n_4645)
);

AOI21xp5_ASAP7_75t_L g4646 ( 
.A1(n_4388),
.A2(n_4255),
.B(n_4173),
.Y(n_4646)
);

O2A1O1Ixp33_ASAP7_75t_L g4647 ( 
.A1(n_4487),
.A2(n_54),
.B(n_52),
.C(n_53),
.Y(n_4647)
);

NAND2xp5_ASAP7_75t_L g4648 ( 
.A(n_4433),
.B(n_52),
.Y(n_4648)
);

INVx5_ASAP7_75t_L g4649 ( 
.A(n_4492),
.Y(n_4649)
);

BUFx2_ASAP7_75t_L g4650 ( 
.A(n_4470),
.Y(n_4650)
);

NOR2xp33_ASAP7_75t_L g4651 ( 
.A(n_4430),
.B(n_53),
.Y(n_4651)
);

INVx3_ASAP7_75t_L g4652 ( 
.A(n_4435),
.Y(n_4652)
);

BUFx3_ASAP7_75t_L g4653 ( 
.A(n_4391),
.Y(n_4653)
);

INVx1_ASAP7_75t_L g4654 ( 
.A(n_4410),
.Y(n_4654)
);

INVx1_ASAP7_75t_L g4655 ( 
.A(n_4410),
.Y(n_4655)
);

AOI21xp5_ASAP7_75t_SL g4656 ( 
.A1(n_4531),
.A2(n_55),
.B(n_56),
.Y(n_4656)
);

OAI22xp5_ASAP7_75t_L g4657 ( 
.A1(n_4554),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_4657)
);

AND2x4_ASAP7_75t_L g4658 ( 
.A(n_4470),
.B(n_58),
.Y(n_4658)
);

INVx1_ASAP7_75t_L g4659 ( 
.A(n_4438),
.Y(n_4659)
);

INVxp67_ASAP7_75t_SL g4660 ( 
.A(n_4484),
.Y(n_4660)
);

OAI22xp5_ASAP7_75t_L g4661 ( 
.A1(n_4606),
.A2(n_62),
.B1(n_59),
.B2(n_60),
.Y(n_4661)
);

INVx4_ASAP7_75t_L g4662 ( 
.A(n_4612),
.Y(n_4662)
);

NOR2xp33_ASAP7_75t_R g4663 ( 
.A(n_4494),
.B(n_63),
.Y(n_4663)
);

OR2x2_ASAP7_75t_L g4664 ( 
.A(n_4457),
.B(n_64),
.Y(n_4664)
);

BUFx3_ASAP7_75t_L g4665 ( 
.A(n_4601),
.Y(n_4665)
);

INVx1_ASAP7_75t_L g4666 ( 
.A(n_4438),
.Y(n_4666)
);

NAND2xp5_ASAP7_75t_L g4667 ( 
.A(n_4562),
.B(n_66),
.Y(n_4667)
);

INVx1_ASAP7_75t_SL g4668 ( 
.A(n_4523),
.Y(n_4668)
);

AND2x2_ASAP7_75t_L g4669 ( 
.A(n_4585),
.B(n_67),
.Y(n_4669)
);

BUFx3_ASAP7_75t_L g4670 ( 
.A(n_4506),
.Y(n_4670)
);

INVx1_ASAP7_75t_L g4671 ( 
.A(n_4450),
.Y(n_4671)
);

NAND2xp5_ASAP7_75t_L g4672 ( 
.A(n_4562),
.B(n_67),
.Y(n_4672)
);

A2O1A1Ixp33_ASAP7_75t_L g4673 ( 
.A1(n_4477),
.A2(n_4456),
.B(n_4401),
.C(n_4483),
.Y(n_4673)
);

INVx2_ASAP7_75t_L g4674 ( 
.A(n_4493),
.Y(n_4674)
);

INVx3_ASAP7_75t_L g4675 ( 
.A(n_4552),
.Y(n_4675)
);

INVx1_ASAP7_75t_L g4676 ( 
.A(n_4450),
.Y(n_4676)
);

INVx2_ASAP7_75t_SL g4677 ( 
.A(n_4423),
.Y(n_4677)
);

INVx3_ASAP7_75t_SL g4678 ( 
.A(n_4622),
.Y(n_4678)
);

AND2x4_ASAP7_75t_L g4679 ( 
.A(n_4382),
.B(n_69),
.Y(n_4679)
);

AOI21xp5_ASAP7_75t_L g4680 ( 
.A1(n_4396),
.A2(n_1753),
.B(n_1725),
.Y(n_4680)
);

A2O1A1Ixp33_ASAP7_75t_L g4681 ( 
.A1(n_4496),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_4681)
);

INVx1_ASAP7_75t_L g4682 ( 
.A(n_4515),
.Y(n_4682)
);

OA21x2_ASAP7_75t_L g4683 ( 
.A1(n_4479),
.A2(n_70),
.B(n_71),
.Y(n_4683)
);

AND2x2_ASAP7_75t_L g4684 ( 
.A(n_4592),
.B(n_4432),
.Y(n_4684)
);

NOR2xp67_ASAP7_75t_SL g4685 ( 
.A(n_4466),
.B(n_1783),
.Y(n_4685)
);

O2A1O1Ixp33_ASAP7_75t_L g4686 ( 
.A1(n_4553),
.A2(n_74),
.B(n_72),
.C(n_73),
.Y(n_4686)
);

INVx1_ASAP7_75t_L g4687 ( 
.A(n_4515),
.Y(n_4687)
);

INVx2_ASAP7_75t_L g4688 ( 
.A(n_4521),
.Y(n_4688)
);

INVx2_ASAP7_75t_SL g4689 ( 
.A(n_4625),
.Y(n_4689)
);

INVx4_ASAP7_75t_L g4690 ( 
.A(n_4373),
.Y(n_4690)
);

AOI22xp5_ASAP7_75t_L g4691 ( 
.A1(n_4441),
.A2(n_1753),
.B1(n_1765),
.B2(n_1725),
.Y(n_4691)
);

AOI22xp33_ASAP7_75t_L g4692 ( 
.A1(n_4618),
.A2(n_4609),
.B1(n_4524),
.B2(n_4613),
.Y(n_4692)
);

NOR2xp67_ASAP7_75t_L g4693 ( 
.A(n_4453),
.B(n_72),
.Y(n_4693)
);

AOI21xp5_ASAP7_75t_L g4694 ( 
.A1(n_4569),
.A2(n_1765),
.B(n_1725),
.Y(n_4694)
);

INVx3_ASAP7_75t_L g4695 ( 
.A(n_4415),
.Y(n_4695)
);

AOI21xp5_ASAP7_75t_L g4696 ( 
.A1(n_4600),
.A2(n_1765),
.B(n_1725),
.Y(n_4696)
);

NAND2xp5_ASAP7_75t_L g4697 ( 
.A(n_4442),
.B(n_4546),
.Y(n_4697)
);

BUFx2_ASAP7_75t_L g4698 ( 
.A(n_4484),
.Y(n_4698)
);

NAND2xp5_ASAP7_75t_L g4699 ( 
.A(n_4546),
.B(n_73),
.Y(n_4699)
);

INVx2_ASAP7_75t_SL g4700 ( 
.A(n_4605),
.Y(n_4700)
);

BUFx12f_ASAP7_75t_L g4701 ( 
.A(n_4570),
.Y(n_4701)
);

INVx2_ASAP7_75t_SL g4702 ( 
.A(n_4458),
.Y(n_4702)
);

BUFx2_ASAP7_75t_L g4703 ( 
.A(n_4425),
.Y(n_4703)
);

NAND2xp5_ASAP7_75t_L g4704 ( 
.A(n_4462),
.B(n_74),
.Y(n_4704)
);

OR2x2_ASAP7_75t_L g4705 ( 
.A(n_4397),
.B(n_75),
.Y(n_4705)
);

AOI21xp5_ASAP7_75t_L g4706 ( 
.A1(n_4566),
.A2(n_1767),
.B(n_1765),
.Y(n_4706)
);

AOI21xp5_ASAP7_75t_L g4707 ( 
.A1(n_4377),
.A2(n_1773),
.B(n_1767),
.Y(n_4707)
);

OR2x6_ASAP7_75t_L g4708 ( 
.A(n_4492),
.B(n_661),
.Y(n_4708)
);

AOI22xp33_ASAP7_75t_L g4709 ( 
.A1(n_4476),
.A2(n_1871),
.B1(n_1875),
.B2(n_1868),
.Y(n_4709)
);

HB1xp67_ASAP7_75t_L g4710 ( 
.A(n_4513),
.Y(n_4710)
);

AND2x2_ASAP7_75t_L g4711 ( 
.A(n_4393),
.B(n_75),
.Y(n_4711)
);

AOI22xp5_ASAP7_75t_L g4712 ( 
.A1(n_4398),
.A2(n_1773),
.B1(n_1783),
.B2(n_1767),
.Y(n_4712)
);

NAND2xp5_ASAP7_75t_L g4713 ( 
.A(n_4464),
.B(n_76),
.Y(n_4713)
);

INVx2_ASAP7_75t_SL g4714 ( 
.A(n_4458),
.Y(n_4714)
);

INVx1_ASAP7_75t_L g4715 ( 
.A(n_4513),
.Y(n_4715)
);

NAND2xp5_ASAP7_75t_L g4716 ( 
.A(n_4530),
.B(n_76),
.Y(n_4716)
);

BUFx6f_ASAP7_75t_L g4717 ( 
.A(n_4373),
.Y(n_4717)
);

CKINVDCx5p33_ASAP7_75t_R g4718 ( 
.A(n_4570),
.Y(n_4718)
);

INVx3_ASAP7_75t_L g4719 ( 
.A(n_4458),
.Y(n_4719)
);

INVx2_ASAP7_75t_L g4720 ( 
.A(n_4369),
.Y(n_4720)
);

AND2x2_ASAP7_75t_L g4721 ( 
.A(n_4383),
.B(n_4490),
.Y(n_4721)
);

A2O1A1Ixp33_ASAP7_75t_L g4722 ( 
.A1(n_4426),
.A2(n_80),
.B(n_77),
.C(n_79),
.Y(n_4722)
);

OAI22xp33_ASAP7_75t_L g4723 ( 
.A1(n_4593),
.A2(n_81),
.B1(n_77),
.B2(n_80),
.Y(n_4723)
);

INVx2_ASAP7_75t_L g4724 ( 
.A(n_4386),
.Y(n_4724)
);

NOR2xp33_ASAP7_75t_L g4725 ( 
.A(n_4571),
.B(n_82),
.Y(n_4725)
);

AND2x4_ASAP7_75t_L g4726 ( 
.A(n_4579),
.B(n_82),
.Y(n_4726)
);

NAND2xp5_ASAP7_75t_L g4727 ( 
.A(n_4548),
.B(n_83),
.Y(n_4727)
);

OR2x6_ASAP7_75t_L g4728 ( 
.A(n_4572),
.B(n_666),
.Y(n_4728)
);

CKINVDCx6p67_ASAP7_75t_R g4729 ( 
.A(n_4580),
.Y(n_4729)
);

NAND2xp5_ASAP7_75t_L g4730 ( 
.A(n_4560),
.B(n_4497),
.Y(n_4730)
);

AND2x2_ASAP7_75t_L g4731 ( 
.A(n_4624),
.B(n_83),
.Y(n_4731)
);

INVx3_ASAP7_75t_L g4732 ( 
.A(n_4459),
.Y(n_4732)
);

INVx2_ASAP7_75t_L g4733 ( 
.A(n_4406),
.Y(n_4733)
);

AND2x4_ASAP7_75t_L g4734 ( 
.A(n_4399),
.B(n_85),
.Y(n_4734)
);

AND2x2_ASAP7_75t_L g4735 ( 
.A(n_4424),
.B(n_85),
.Y(n_4735)
);

AND2x2_ASAP7_75t_L g4736 ( 
.A(n_4602),
.B(n_86),
.Y(n_4736)
);

AND2x4_ASAP7_75t_L g4737 ( 
.A(n_4399),
.B(n_86),
.Y(n_4737)
);

INVx1_ASAP7_75t_L g4738 ( 
.A(n_4544),
.Y(n_4738)
);

BUFx6f_ASAP7_75t_L g4739 ( 
.A(n_4373),
.Y(n_4739)
);

NAND2x1p5_ASAP7_75t_L g4740 ( 
.A(n_4574),
.B(n_1767),
.Y(n_4740)
);

NAND2xp5_ASAP7_75t_L g4741 ( 
.A(n_4555),
.B(n_87),
.Y(n_4741)
);

O2A1O1Ixp33_ASAP7_75t_L g4742 ( 
.A1(n_4473),
.A2(n_90),
.B(n_88),
.C(n_89),
.Y(n_4742)
);

AND2x2_ASAP7_75t_L g4743 ( 
.A(n_4459),
.B(n_88),
.Y(n_4743)
);

INVx1_ASAP7_75t_L g4744 ( 
.A(n_4420),
.Y(n_4744)
);

INVx2_ASAP7_75t_L g4745 ( 
.A(n_4421),
.Y(n_4745)
);

INVx2_ASAP7_75t_L g4746 ( 
.A(n_4454),
.Y(n_4746)
);

AOI21xp5_ASAP7_75t_L g4747 ( 
.A1(n_4381),
.A2(n_1783),
.B(n_1773),
.Y(n_4747)
);

INVx4_ASAP7_75t_SL g4748 ( 
.A(n_4378),
.Y(n_4748)
);

NAND2xp5_ASAP7_75t_L g4749 ( 
.A(n_4434),
.B(n_91),
.Y(n_4749)
);

BUFx2_ASAP7_75t_R g4750 ( 
.A(n_4465),
.Y(n_4750)
);

AND2x4_ASAP7_75t_L g4751 ( 
.A(n_4495),
.B(n_91),
.Y(n_4751)
);

AND2x2_ASAP7_75t_L g4752 ( 
.A(n_4459),
.B(n_92),
.Y(n_4752)
);

NAND2xp5_ASAP7_75t_L g4753 ( 
.A(n_4575),
.B(n_92),
.Y(n_4753)
);

AND2x2_ASAP7_75t_L g4754 ( 
.A(n_4522),
.B(n_93),
.Y(n_4754)
);

AND2x4_ASAP7_75t_L g4755 ( 
.A(n_4495),
.B(n_93),
.Y(n_4755)
);

BUFx2_ASAP7_75t_L g4756 ( 
.A(n_4425),
.Y(n_4756)
);

NAND2xp5_ASAP7_75t_L g4757 ( 
.A(n_4598),
.B(n_94),
.Y(n_4757)
);

AOI21xp5_ASAP7_75t_L g4758 ( 
.A1(n_4449),
.A2(n_1783),
.B(n_1773),
.Y(n_4758)
);

NAND2xp5_ASAP7_75t_L g4759 ( 
.A(n_4615),
.B(n_95),
.Y(n_4759)
);

AND2x2_ASAP7_75t_L g4760 ( 
.A(n_4522),
.B(n_97),
.Y(n_4760)
);

NAND2xp5_ASAP7_75t_L g4761 ( 
.A(n_4589),
.B(n_97),
.Y(n_4761)
);

OR2x2_ASAP7_75t_L g4762 ( 
.A(n_4440),
.B(n_98),
.Y(n_4762)
);

CKINVDCx5p33_ASAP7_75t_R g4763 ( 
.A(n_4595),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_4616),
.Y(n_4764)
);

INVx1_ASAP7_75t_L g4765 ( 
.A(n_4573),
.Y(n_4765)
);

NAND2xp5_ASAP7_75t_L g4766 ( 
.A(n_4596),
.B(n_99),
.Y(n_4766)
);

OR2x2_ASAP7_75t_L g4767 ( 
.A(n_4603),
.B(n_4586),
.Y(n_4767)
);

AOI22xp5_ASAP7_75t_L g4768 ( 
.A1(n_4499),
.A2(n_1789),
.B1(n_1796),
.B2(n_1784),
.Y(n_4768)
);

HB1xp67_ASAP7_75t_L g4769 ( 
.A(n_4517),
.Y(n_4769)
);

INVx1_ASAP7_75t_SL g4770 ( 
.A(n_4378),
.Y(n_4770)
);

OR2x2_ASAP7_75t_L g4771 ( 
.A(n_4468),
.B(n_99),
.Y(n_4771)
);

BUFx2_ASAP7_75t_L g4772 ( 
.A(n_4425),
.Y(n_4772)
);

BUFx4f_ASAP7_75t_SL g4773 ( 
.A(n_4378),
.Y(n_4773)
);

BUFx3_ASAP7_75t_L g4774 ( 
.A(n_4387),
.Y(n_4774)
);

NAND2xp5_ASAP7_75t_L g4775 ( 
.A(n_4419),
.B(n_100),
.Y(n_4775)
);

INVx2_ASAP7_75t_L g4776 ( 
.A(n_4379),
.Y(n_4776)
);

INVx1_ASAP7_75t_L g4777 ( 
.A(n_4479),
.Y(n_4777)
);

NOR2xp33_ASAP7_75t_L g4778 ( 
.A(n_4445),
.B(n_102),
.Y(n_4778)
);

INVx2_ASAP7_75t_L g4779 ( 
.A(n_4379),
.Y(n_4779)
);

BUFx2_ASAP7_75t_L g4780 ( 
.A(n_4489),
.Y(n_4780)
);

A2O1A1Ixp33_ASAP7_75t_L g4781 ( 
.A1(n_4395),
.A2(n_105),
.B(n_102),
.C(n_103),
.Y(n_4781)
);

INVx1_ASAP7_75t_L g4782 ( 
.A(n_4489),
.Y(n_4782)
);

CKINVDCx20_ASAP7_75t_R g4783 ( 
.A(n_4436),
.Y(n_4783)
);

NAND2xp5_ASAP7_75t_L g4784 ( 
.A(n_4427),
.B(n_106),
.Y(n_4784)
);

INVx1_ASAP7_75t_L g4785 ( 
.A(n_4503),
.Y(n_4785)
);

INVx3_ASAP7_75t_L g4786 ( 
.A(n_4522),
.Y(n_4786)
);

BUFx12f_ASAP7_75t_L g4787 ( 
.A(n_4387),
.Y(n_4787)
);

NOR2xp33_ASAP7_75t_L g4788 ( 
.A(n_4371),
.B(n_109),
.Y(n_4788)
);

OAI21xp5_ASAP7_75t_L g4789 ( 
.A1(n_4404),
.A2(n_109),
.B(n_110),
.Y(n_4789)
);

OA21x2_ASAP7_75t_L g4790 ( 
.A1(n_4503),
.A2(n_110),
.B(n_111),
.Y(n_4790)
);

BUFx2_ASAP7_75t_L g4791 ( 
.A(n_4379),
.Y(n_4791)
);

AOI22xp5_ASAP7_75t_L g4792 ( 
.A1(n_4537),
.A2(n_4501),
.B1(n_4527),
.B2(n_4500),
.Y(n_4792)
);

INVx3_ASAP7_75t_L g4793 ( 
.A(n_4535),
.Y(n_4793)
);

BUFx6f_ASAP7_75t_L g4794 ( 
.A(n_4387),
.Y(n_4794)
);

OAI21x1_ASAP7_75t_L g4795 ( 
.A1(n_4505),
.A2(n_670),
.B(n_669),
.Y(n_4795)
);

INVx3_ASAP7_75t_SL g4796 ( 
.A(n_4535),
.Y(n_4796)
);

AND2x2_ASAP7_75t_L g4797 ( 
.A(n_4535),
.B(n_112),
.Y(n_4797)
);

INVx1_ASAP7_75t_L g4798 ( 
.A(n_4576),
.Y(n_4798)
);

OAI22xp5_ASAP7_75t_L g4799 ( 
.A1(n_4471),
.A2(n_114),
.B1(n_112),
.B2(n_113),
.Y(n_4799)
);

NAND2xp5_ASAP7_75t_L g4800 ( 
.A(n_4481),
.B(n_114),
.Y(n_4800)
);

NOR2x1_ASAP7_75t_SL g4801 ( 
.A(n_4594),
.B(n_1784),
.Y(n_4801)
);

INVx3_ASAP7_75t_L g4802 ( 
.A(n_4561),
.Y(n_4802)
);

AOI21xp5_ASAP7_75t_L g4803 ( 
.A1(n_4411),
.A2(n_1789),
.B(n_1784),
.Y(n_4803)
);

INVx1_ASAP7_75t_L g4804 ( 
.A(n_4576),
.Y(n_4804)
);

NAND2xp5_ASAP7_75t_L g4805 ( 
.A(n_4491),
.B(n_115),
.Y(n_4805)
);

BUFx6f_ASAP7_75t_L g4806 ( 
.A(n_4561),
.Y(n_4806)
);

INVx5_ASAP7_75t_L g4807 ( 
.A(n_4594),
.Y(n_4807)
);

INVx2_ASAP7_75t_SL g4808 ( 
.A(n_4561),
.Y(n_4808)
);

INVx1_ASAP7_75t_L g4809 ( 
.A(n_4576),
.Y(n_4809)
);

AND2x4_ASAP7_75t_L g4810 ( 
.A(n_4617),
.B(n_116),
.Y(n_4810)
);

INVx3_ASAP7_75t_L g4811 ( 
.A(n_4617),
.Y(n_4811)
);

NAND2xp5_ASAP7_75t_L g4812 ( 
.A(n_4510),
.B(n_117),
.Y(n_4812)
);

INVx1_ASAP7_75t_L g4813 ( 
.A(n_4480),
.Y(n_4813)
);

BUFx3_ASAP7_75t_L g4814 ( 
.A(n_4617),
.Y(n_4814)
);

INVx1_ASAP7_75t_L g4815 ( 
.A(n_4480),
.Y(n_4815)
);

NOR2x1_ASAP7_75t_L g4816 ( 
.A(n_4567),
.B(n_118),
.Y(n_4816)
);

INVx1_ASAP7_75t_L g4817 ( 
.A(n_4480),
.Y(n_4817)
);

AOI21xp5_ASAP7_75t_L g4818 ( 
.A1(n_4472),
.A2(n_1789),
.B(n_1784),
.Y(n_4818)
);

INVx1_ASAP7_75t_L g4819 ( 
.A(n_4374),
.Y(n_4819)
);

BUFx6f_ASAP7_75t_L g4820 ( 
.A(n_4502),
.Y(n_4820)
);

INVx1_ASAP7_75t_L g4821 ( 
.A(n_4374),
.Y(n_4821)
);

AOI22xp33_ASAP7_75t_L g4822 ( 
.A1(n_4428),
.A2(n_1871),
.B1(n_1875),
.B2(n_1868),
.Y(n_4822)
);

BUFx2_ASAP7_75t_L g4823 ( 
.A(n_4455),
.Y(n_4823)
);

AND2x2_ASAP7_75t_L g4824 ( 
.A(n_4518),
.B(n_4549),
.Y(n_4824)
);

A2O1A1Ixp33_ASAP7_75t_L g4825 ( 
.A1(n_4422),
.A2(n_4516),
.B(n_4525),
.C(n_4551),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4374),
.Y(n_4826)
);

AOI21xp5_ASAP7_75t_L g4827 ( 
.A1(n_4508),
.A2(n_1796),
.B(n_1789),
.Y(n_4827)
);

INVx1_ASAP7_75t_L g4828 ( 
.A(n_4485),
.Y(n_4828)
);

BUFx6f_ASAP7_75t_L g4829 ( 
.A(n_4502),
.Y(n_4829)
);

AOI21xp5_ASAP7_75t_L g4830 ( 
.A1(n_4394),
.A2(n_1820),
.B(n_1796),
.Y(n_4830)
);

BUFx6f_ASAP7_75t_L g4831 ( 
.A(n_4581),
.Y(n_4831)
);

AOI21xp5_ASAP7_75t_L g4832 ( 
.A1(n_4578),
.A2(n_1820),
.B(n_1796),
.Y(n_4832)
);

INVx2_ASAP7_75t_L g4833 ( 
.A(n_4368),
.Y(n_4833)
);

AND2x4_ASAP7_75t_L g4834 ( 
.A(n_4519),
.B(n_118),
.Y(n_4834)
);

NAND2x1p5_ASAP7_75t_L g4835 ( 
.A(n_4559),
.B(n_1820),
.Y(n_4835)
);

AND2x2_ASAP7_75t_L g4836 ( 
.A(n_4437),
.B(n_119),
.Y(n_4836)
);

O2A1O1Ixp33_ASAP7_75t_L g4837 ( 
.A1(n_4520),
.A2(n_122),
.B(n_119),
.C(n_120),
.Y(n_4837)
);

BUFx6f_ASAP7_75t_L g4838 ( 
.A(n_4564),
.Y(n_4838)
);

INVx2_ASAP7_75t_L g4839 ( 
.A(n_4368),
.Y(n_4839)
);

AND2x2_ASAP7_75t_L g4840 ( 
.A(n_4428),
.B(n_120),
.Y(n_4840)
);

AND2x4_ASAP7_75t_L g4841 ( 
.A(n_4447),
.B(n_123),
.Y(n_4841)
);

BUFx3_ASAP7_75t_L g4842 ( 
.A(n_4402),
.Y(n_4842)
);

INVx1_ASAP7_75t_SL g4843 ( 
.A(n_4372),
.Y(n_4843)
);

NAND2xp5_ASAP7_75t_L g4844 ( 
.A(n_4380),
.B(n_123),
.Y(n_4844)
);

NAND2xp5_ASAP7_75t_L g4845 ( 
.A(n_4439),
.B(n_124),
.Y(n_4845)
);

INVx1_ASAP7_75t_L g4846 ( 
.A(n_4485),
.Y(n_4846)
);

AOI21xp5_ASAP7_75t_L g4847 ( 
.A1(n_4403),
.A2(n_1823),
.B(n_1820),
.Y(n_4847)
);

INVx5_ASAP7_75t_L g4848 ( 
.A(n_4413),
.Y(n_4848)
);

AND2x2_ASAP7_75t_L g4849 ( 
.A(n_4619),
.B(n_124),
.Y(n_4849)
);

AND2x4_ASAP7_75t_L g4850 ( 
.A(n_4447),
.B(n_125),
.Y(n_4850)
);

OAI22xp5_ASAP7_75t_SL g4851 ( 
.A1(n_4431),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_4851)
);

CKINVDCx5p33_ASAP7_75t_R g4852 ( 
.A(n_4446),
.Y(n_4852)
);

INVx1_ASAP7_75t_L g4853 ( 
.A(n_4485),
.Y(n_4853)
);

AOI21xp5_ASAP7_75t_L g4854 ( 
.A1(n_4620),
.A2(n_1828),
.B(n_1823),
.Y(n_4854)
);

NOR3xp33_ASAP7_75t_L g4855 ( 
.A(n_4408),
.B(n_126),
.C(n_128),
.Y(n_4855)
);

AND2x2_ASAP7_75t_L g4856 ( 
.A(n_4447),
.B(n_130),
.Y(n_4856)
);

OAI22xp5_ASAP7_75t_L g4857 ( 
.A1(n_4412),
.A2(n_4405),
.B1(n_4507),
.B2(n_4604),
.Y(n_4857)
);

CKINVDCx20_ASAP7_75t_R g4858 ( 
.A(n_4583),
.Y(n_4858)
);

NAND2xp5_ASAP7_75t_L g4859 ( 
.A(n_4540),
.B(n_130),
.Y(n_4859)
);

OR2x6_ASAP7_75t_L g4860 ( 
.A(n_4614),
.B(n_4547),
.Y(n_4860)
);

NAND2xp5_ASAP7_75t_L g4861 ( 
.A(n_4528),
.B(n_131),
.Y(n_4861)
);

INVx2_ASAP7_75t_SL g4862 ( 
.A(n_4514),
.Y(n_4862)
);

INVx1_ASAP7_75t_L g4863 ( 
.A(n_4368),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4538),
.Y(n_4864)
);

AOI22xp5_ASAP7_75t_L g4865 ( 
.A1(n_4478),
.A2(n_1828),
.B1(n_1831),
.B2(n_1823),
.Y(n_4865)
);

NAND2xp5_ASAP7_75t_L g4866 ( 
.A(n_4584),
.B(n_131),
.Y(n_4866)
);

NAND2xp33_ASAP7_75t_L g4867 ( 
.A(n_4542),
.B(n_133),
.Y(n_4867)
);

INVx2_ASAP7_75t_L g4868 ( 
.A(n_4498),
.Y(n_4868)
);

HB1xp67_ASAP7_75t_L g4869 ( 
.A(n_4526),
.Y(n_4869)
);

INVx3_ASAP7_75t_L g4870 ( 
.A(n_4563),
.Y(n_4870)
);

NAND2xp5_ASAP7_75t_SL g4871 ( 
.A(n_4623),
.B(n_1823),
.Y(n_4871)
);

INVx2_ASAP7_75t_L g4872 ( 
.A(n_4451),
.Y(n_4872)
);

INVx2_ASAP7_75t_SL g4873 ( 
.A(n_4689),
.Y(n_4873)
);

BUFx6f_ASAP7_75t_L g4874 ( 
.A(n_4701),
.Y(n_4874)
);

INVx5_ASAP7_75t_L g4875 ( 
.A(n_4728),
.Y(n_4875)
);

AOI22xp33_ASAP7_75t_L g4876 ( 
.A1(n_4651),
.A2(n_4582),
.B1(n_4478),
.B2(n_4532),
.Y(n_4876)
);

INVx1_ASAP7_75t_L g4877 ( 
.A(n_4650),
.Y(n_4877)
);

AOI22xp33_ASAP7_75t_L g4878 ( 
.A1(n_4851),
.A2(n_4590),
.B1(n_4533),
.B2(n_4539),
.Y(n_4878)
);

OAI22xp33_ASAP7_75t_L g4879 ( 
.A1(n_4635),
.A2(n_4463),
.B1(n_4429),
.B2(n_4590),
.Y(n_4879)
);

CKINVDCx11_ASAP7_75t_R g4880 ( 
.A(n_4678),
.Y(n_4880)
);

BUFx2_ASAP7_75t_L g4881 ( 
.A(n_4629),
.Y(n_4881)
);

INVx2_ASAP7_75t_L g4882 ( 
.A(n_4674),
.Y(n_4882)
);

BUFx2_ASAP7_75t_L g4883 ( 
.A(n_4675),
.Y(n_4883)
);

CKINVDCx11_ASAP7_75t_R g4884 ( 
.A(n_4670),
.Y(n_4884)
);

INVx2_ASAP7_75t_L g4885 ( 
.A(n_4688),
.Y(n_4885)
);

INVx2_ASAP7_75t_L g4886 ( 
.A(n_4710),
.Y(n_4886)
);

OAI21xp5_ASAP7_75t_SL g4887 ( 
.A1(n_4725),
.A2(n_4611),
.B(n_4384),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4650),
.Y(n_4888)
);

INVx6_ASAP7_75t_L g4889 ( 
.A(n_4662),
.Y(n_4889)
);

AOI22xp33_ASAP7_75t_L g4890 ( 
.A1(n_4635),
.A2(n_4482),
.B1(n_4486),
.B2(n_4626),
.Y(n_4890)
);

AOI22xp33_ASAP7_75t_SL g4891 ( 
.A1(n_4683),
.A2(n_4550),
.B1(n_4461),
.B2(n_4469),
.Y(n_4891)
);

BUFx5_ASAP7_75t_L g4892 ( 
.A(n_4841),
.Y(n_4892)
);

NAND2xp5_ASAP7_75t_L g4893 ( 
.A(n_4643),
.B(n_4504),
.Y(n_4893)
);

CKINVDCx11_ASAP7_75t_R g4894 ( 
.A(n_4653),
.Y(n_4894)
);

INVx1_ASAP7_75t_L g4895 ( 
.A(n_4632),
.Y(n_4895)
);

INVx2_ASAP7_75t_L g4896 ( 
.A(n_4715),
.Y(n_4896)
);

AOI22xp33_ASAP7_75t_SL g4897 ( 
.A1(n_4683),
.A2(n_4467),
.B1(n_4414),
.B2(n_4558),
.Y(n_4897)
);

BUFx4f_ASAP7_75t_SL g4898 ( 
.A(n_4677),
.Y(n_4898)
);

NAND2xp5_ASAP7_75t_L g4899 ( 
.A(n_4764),
.B(n_4511),
.Y(n_4899)
);

INVx6_ASAP7_75t_L g4900 ( 
.A(n_4665),
.Y(n_4900)
);

OAI22xp5_ASAP7_75t_L g4901 ( 
.A1(n_4673),
.A2(n_4541),
.B1(n_4621),
.B2(n_4545),
.Y(n_4901)
);

OAI22xp5_ASAP7_75t_SL g4902 ( 
.A1(n_4718),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_4902)
);

OAI22xp5_ASAP7_75t_L g4903 ( 
.A1(n_4681),
.A2(n_4565),
.B1(n_138),
.B2(n_136),
.Y(n_4903)
);

AOI22xp33_ASAP7_75t_L g4904 ( 
.A1(n_4855),
.A2(n_4529),
.B1(n_4536),
.B2(n_4556),
.Y(n_4904)
);

INVx1_ASAP7_75t_SL g4905 ( 
.A(n_4750),
.Y(n_4905)
);

BUFx8_ASAP7_75t_SL g4906 ( 
.A(n_4652),
.Y(n_4906)
);

OAI22xp33_ASAP7_75t_L g4907 ( 
.A1(n_4641),
.A2(n_4599),
.B1(n_4588),
.B2(n_4597),
.Y(n_4907)
);

INVx1_ASAP7_75t_L g4908 ( 
.A(n_4642),
.Y(n_4908)
);

CKINVDCx20_ASAP7_75t_R g4909 ( 
.A(n_4783),
.Y(n_4909)
);

CKINVDCx20_ASAP7_75t_R g4910 ( 
.A(n_4663),
.Y(n_4910)
);

AOI22xp33_ASAP7_75t_L g4911 ( 
.A1(n_4789),
.A2(n_4557),
.B1(n_4607),
.B2(n_4610),
.Y(n_4911)
);

INVx6_ASAP7_75t_L g4912 ( 
.A(n_4787),
.Y(n_4912)
);

INVx1_ASAP7_75t_L g4913 ( 
.A(n_4654),
.Y(n_4913)
);

BUFx10_ASAP7_75t_L g4914 ( 
.A(n_4726),
.Y(n_4914)
);

BUFx10_ASAP7_75t_L g4915 ( 
.A(n_4726),
.Y(n_4915)
);

BUFx10_ASAP7_75t_L g4916 ( 
.A(n_4778),
.Y(n_4916)
);

INVx2_ASAP7_75t_L g4917 ( 
.A(n_4720),
.Y(n_4917)
);

OA21x2_ASAP7_75t_L g4918 ( 
.A1(n_4660),
.A2(n_4577),
.B(n_4407),
.Y(n_4918)
);

AND2x2_ASAP7_75t_L g4919 ( 
.A(n_4700),
.B(n_4460),
.Y(n_4919)
);

AOI22xp33_ASAP7_75t_SL g4920 ( 
.A1(n_4790),
.A2(n_4452),
.B1(n_4418),
.B2(n_4448),
.Y(n_4920)
);

INVx1_ASAP7_75t_L g4921 ( 
.A(n_4655),
.Y(n_4921)
);

BUFx2_ASAP7_75t_L g4922 ( 
.A(n_4631),
.Y(n_4922)
);

AOI22xp33_ASAP7_75t_L g4923 ( 
.A1(n_4843),
.A2(n_4385),
.B1(n_4409),
.B2(n_4417),
.Y(n_4923)
);

BUFx8_ASAP7_75t_L g4924 ( 
.A(n_4735),
.Y(n_4924)
);

AOI22xp33_ASAP7_75t_L g4925 ( 
.A1(n_4842),
.A2(n_4509),
.B1(n_4392),
.B2(n_4568),
.Y(n_4925)
);

AOI22xp33_ASAP7_75t_L g4926 ( 
.A1(n_4661),
.A2(n_4474),
.B1(n_4475),
.B2(n_1888),
.Y(n_4926)
);

OAI22xp5_ASAP7_75t_L g4927 ( 
.A1(n_4781),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.Y(n_4927)
);

CKINVDCx20_ASAP7_75t_R g4928 ( 
.A(n_4763),
.Y(n_4928)
);

CKINVDCx6p67_ASAP7_75t_R g4929 ( 
.A(n_4729),
.Y(n_4929)
);

INVx1_ASAP7_75t_L g4930 ( 
.A(n_4659),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_4666),
.Y(n_4931)
);

INVx2_ASAP7_75t_L g4932 ( 
.A(n_4724),
.Y(n_4932)
);

BUFx8_ASAP7_75t_L g4933 ( 
.A(n_4711),
.Y(n_4933)
);

AOI22xp33_ASAP7_75t_L g4934 ( 
.A1(n_4692),
.A2(n_1888),
.B1(n_1896),
.B2(n_1883),
.Y(n_4934)
);

BUFx6f_ASAP7_75t_L g4935 ( 
.A(n_4717),
.Y(n_4935)
);

HB1xp67_ASAP7_75t_L g4936 ( 
.A(n_4684),
.Y(n_4936)
);

AOI21xp5_ASAP7_75t_L g4937 ( 
.A1(n_4639),
.A2(n_4599),
.B(n_1831),
.Y(n_4937)
);

OAI22xp33_ASAP7_75t_L g4938 ( 
.A1(n_4641),
.A2(n_4599),
.B1(n_143),
.B2(n_140),
.Y(n_4938)
);

INVx1_ASAP7_75t_L g4939 ( 
.A(n_4671),
.Y(n_4939)
);

INVx1_ASAP7_75t_L g4940 ( 
.A(n_4676),
.Y(n_4940)
);

INVxp67_ASAP7_75t_SL g4941 ( 
.A(n_4698),
.Y(n_4941)
);

INVx2_ASAP7_75t_L g4942 ( 
.A(n_4733),
.Y(n_4942)
);

BUFx8_ASAP7_75t_L g4943 ( 
.A(n_4736),
.Y(n_4943)
);

BUFx4f_ASAP7_75t_SL g4944 ( 
.A(n_4668),
.Y(n_4944)
);

AOI22xp33_ASAP7_75t_L g4945 ( 
.A1(n_4799),
.A2(n_1888),
.B1(n_1896),
.B2(n_1883),
.Y(n_4945)
);

INVx4_ASAP7_75t_SL g4946 ( 
.A(n_4796),
.Y(n_4946)
);

AOI22xp33_ASAP7_75t_L g4947 ( 
.A1(n_4657),
.A2(n_1888),
.B1(n_1896),
.B2(n_1883),
.Y(n_4947)
);

BUFx8_ASAP7_75t_L g4948 ( 
.A(n_4640),
.Y(n_4948)
);

BUFx8_ASAP7_75t_L g4949 ( 
.A(n_4669),
.Y(n_4949)
);

AOI22xp33_ASAP7_75t_L g4950 ( 
.A1(n_4788),
.A2(n_1896),
.B1(n_1910),
.B2(n_1883),
.Y(n_4950)
);

INVx6_ASAP7_75t_L g4951 ( 
.A(n_4628),
.Y(n_4951)
);

INVx2_ASAP7_75t_L g4952 ( 
.A(n_4745),
.Y(n_4952)
);

OAI22xp5_ASAP7_75t_L g4953 ( 
.A1(n_4792),
.A2(n_145),
.B1(n_140),
.B2(n_142),
.Y(n_4953)
);

INVx3_ASAP7_75t_SL g4954 ( 
.A(n_4852),
.Y(n_4954)
);

INVx1_ASAP7_75t_L g4955 ( 
.A(n_4682),
.Y(n_4955)
);

INVx8_ASAP7_75t_L g4956 ( 
.A(n_4734),
.Y(n_4956)
);

INVx3_ASAP7_75t_L g4957 ( 
.A(n_4628),
.Y(n_4957)
);

INVx6_ASAP7_75t_L g4958 ( 
.A(n_4645),
.Y(n_4958)
);

OAI22xp33_ASAP7_75t_L g4959 ( 
.A1(n_4728),
.A2(n_146),
.B1(n_142),
.B2(n_145),
.Y(n_4959)
);

AOI22xp33_ASAP7_75t_SL g4960 ( 
.A1(n_4790),
.A2(n_4698),
.B1(n_4856),
.B2(n_4848),
.Y(n_4960)
);

INVx2_ASAP7_75t_L g4961 ( 
.A(n_4746),
.Y(n_4961)
);

AOI22xp33_ASAP7_75t_SL g4962 ( 
.A1(n_4848),
.A2(n_148),
.B1(n_146),
.B2(n_147),
.Y(n_4962)
);

INVx1_ASAP7_75t_L g4963 ( 
.A(n_4687),
.Y(n_4963)
);

BUFx3_ASAP7_75t_L g4964 ( 
.A(n_4645),
.Y(n_4964)
);

INVx2_ASAP7_75t_SL g4965 ( 
.A(n_4630),
.Y(n_4965)
);

BUFx10_ASAP7_75t_L g4966 ( 
.A(n_4734),
.Y(n_4966)
);

CKINVDCx11_ASAP7_75t_R g4967 ( 
.A(n_4770),
.Y(n_4967)
);

INVx1_ASAP7_75t_L g4968 ( 
.A(n_4697),
.Y(n_4968)
);

OAI22xp5_ASAP7_75t_L g4969 ( 
.A1(n_4722),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_4969)
);

OAI22xp5_ASAP7_75t_L g4970 ( 
.A1(n_4634),
.A2(n_152),
.B1(n_149),
.B2(n_150),
.Y(n_4970)
);

CKINVDCx20_ASAP7_75t_R g4971 ( 
.A(n_4773),
.Y(n_4971)
);

INVx3_ASAP7_75t_L g4972 ( 
.A(n_4820),
.Y(n_4972)
);

CKINVDCx11_ASAP7_75t_R g4973 ( 
.A(n_4717),
.Y(n_4973)
);

BUFx2_ASAP7_75t_L g4974 ( 
.A(n_4824),
.Y(n_4974)
);

OAI22xp5_ASAP7_75t_L g4975 ( 
.A1(n_4825),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_4975)
);

CKINVDCx11_ASAP7_75t_R g4976 ( 
.A(n_4739),
.Y(n_4976)
);

AOI22xp33_ASAP7_75t_SL g4977 ( 
.A1(n_4848),
.A2(n_4840),
.B1(n_4857),
.B2(n_4850),
.Y(n_4977)
);

HB1xp67_ASAP7_75t_L g4978 ( 
.A(n_4780),
.Y(n_4978)
);

CKINVDCx6p67_ASAP7_75t_R g4979 ( 
.A(n_4814),
.Y(n_4979)
);

BUFx6f_ASAP7_75t_L g4980 ( 
.A(n_4739),
.Y(n_4980)
);

INVx2_ASAP7_75t_L g4981 ( 
.A(n_4744),
.Y(n_4981)
);

BUFx8_ASAP7_75t_L g4982 ( 
.A(n_4836),
.Y(n_4982)
);

INVx5_ASAP7_75t_L g4983 ( 
.A(n_4708),
.Y(n_4983)
);

NAND2xp5_ASAP7_75t_L g4984 ( 
.A(n_4658),
.B(n_153),
.Y(n_4984)
);

OAI22xp5_ASAP7_75t_L g4985 ( 
.A1(n_4866),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_4985)
);

OAI22xp33_ASAP7_75t_L g4986 ( 
.A1(n_4691),
.A2(n_160),
.B1(n_156),
.B2(n_159),
.Y(n_4986)
);

INVx6_ASAP7_75t_L g4987 ( 
.A(n_4748),
.Y(n_4987)
);

OAI22xp33_ASAP7_75t_L g4988 ( 
.A1(n_4708),
.A2(n_161),
.B1(n_159),
.B2(n_160),
.Y(n_4988)
);

AOI22xp33_ASAP7_75t_L g4989 ( 
.A1(n_4693),
.A2(n_1922),
.B1(n_1931),
.B2(n_1910),
.Y(n_4989)
);

AOI22xp33_ASAP7_75t_SL g4990 ( 
.A1(n_4841),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.Y(n_4990)
);

BUFx6f_ASAP7_75t_L g4991 ( 
.A(n_4794),
.Y(n_4991)
);

INVx2_ASAP7_75t_L g4992 ( 
.A(n_4738),
.Y(n_4992)
);

OAI21xp5_ASAP7_75t_L g4993 ( 
.A1(n_4686),
.A2(n_164),
.B(n_165),
.Y(n_4993)
);

AOI22xp33_ASAP7_75t_L g4994 ( 
.A1(n_4767),
.A2(n_1922),
.B1(n_1931),
.B2(n_1910),
.Y(n_4994)
);

BUFx3_ASAP7_75t_L g4995 ( 
.A(n_4721),
.Y(n_4995)
);

OAI22xp33_ASAP7_75t_L g4996 ( 
.A1(n_4638),
.A2(n_167),
.B1(n_164),
.B2(n_166),
.Y(n_4996)
);

INVx1_ASAP7_75t_L g4997 ( 
.A(n_4777),
.Y(n_4997)
);

INVx2_ASAP7_75t_L g4998 ( 
.A(n_4765),
.Y(n_4998)
);

INVx1_ASAP7_75t_L g4999 ( 
.A(n_4782),
.Y(n_4999)
);

BUFx8_ASAP7_75t_L g5000 ( 
.A(n_4731),
.Y(n_5000)
);

INVx1_ASAP7_75t_L g5001 ( 
.A(n_4785),
.Y(n_5001)
);

INVx1_ASAP7_75t_SL g5002 ( 
.A(n_4762),
.Y(n_5002)
);

INVx1_ASAP7_75t_L g5003 ( 
.A(n_4780),
.Y(n_5003)
);

BUFx2_ASAP7_75t_L g5004 ( 
.A(n_4774),
.Y(n_5004)
);

AOI22xp33_ASAP7_75t_L g5005 ( 
.A1(n_4730),
.A2(n_1922),
.B1(n_1931),
.B2(n_1910),
.Y(n_5005)
);

BUFx8_ASAP7_75t_L g5006 ( 
.A(n_4705),
.Y(n_5006)
);

INVx1_ASAP7_75t_L g5007 ( 
.A(n_4769),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_4667),
.Y(n_5008)
);

BUFx8_ASAP7_75t_SL g5009 ( 
.A(n_4695),
.Y(n_5009)
);

BUFx2_ASAP7_75t_L g5010 ( 
.A(n_4702),
.Y(n_5010)
);

INVx2_ASAP7_75t_L g5011 ( 
.A(n_4850),
.Y(n_5011)
);

NAND2xp5_ASAP7_75t_L g5012 ( 
.A(n_4658),
.B(n_166),
.Y(n_5012)
);

BUFx3_ASAP7_75t_L g5013 ( 
.A(n_4737),
.Y(n_5013)
);

OAI22xp5_ASAP7_75t_L g5014 ( 
.A1(n_4627),
.A2(n_169),
.B1(n_167),
.B2(n_168),
.Y(n_5014)
);

INVx1_ASAP7_75t_L g5015 ( 
.A(n_4672),
.Y(n_5015)
);

AOI22xp33_ASAP7_75t_SL g5016 ( 
.A1(n_4703),
.A2(n_171),
.B1(n_168),
.B2(n_169),
.Y(n_5016)
);

INVx2_ASAP7_75t_L g5017 ( 
.A(n_4703),
.Y(n_5017)
);

INVx1_ASAP7_75t_L g5018 ( 
.A(n_4699),
.Y(n_5018)
);

AOI22xp33_ASAP7_75t_L g5019 ( 
.A1(n_4822),
.A2(n_4646),
.B1(n_4644),
.B2(n_4858),
.Y(n_5019)
);

NAND2xp5_ASAP7_75t_L g5020 ( 
.A(n_4704),
.B(n_4679),
.Y(n_5020)
);

AOI22xp5_ASAP7_75t_L g5021 ( 
.A1(n_4867),
.A2(n_1831),
.B1(n_1828),
.B2(n_174),
.Y(n_5021)
);

OAI22xp5_ASAP7_75t_L g5022 ( 
.A1(n_4757),
.A2(n_175),
.B1(n_171),
.B2(n_172),
.Y(n_5022)
);

CKINVDCx6p67_ASAP7_75t_R g5023 ( 
.A(n_4771),
.Y(n_5023)
);

INVx4_ASAP7_75t_L g5024 ( 
.A(n_4794),
.Y(n_5024)
);

BUFx12f_ASAP7_75t_L g5025 ( 
.A(n_4664),
.Y(n_5025)
);

AOI22xp33_ASAP7_75t_L g5026 ( 
.A1(n_4709),
.A2(n_1931),
.B1(n_1922),
.B2(n_1831),
.Y(n_5026)
);

AOI22xp33_ASAP7_75t_L g5027 ( 
.A1(n_4749),
.A2(n_1828),
.B1(n_177),
.B2(n_175),
.Y(n_5027)
);

CKINVDCx6p67_ASAP7_75t_R g5028 ( 
.A(n_4713),
.Y(n_5028)
);

INVx1_ASAP7_75t_L g5029 ( 
.A(n_4679),
.Y(n_5029)
);

OAI22xp5_ASAP7_75t_L g5030 ( 
.A1(n_4759),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_5030)
);

CKINVDCx11_ASAP7_75t_R g5031 ( 
.A(n_4806),
.Y(n_5031)
);

BUFx10_ASAP7_75t_L g5032 ( 
.A(n_4737),
.Y(n_5032)
);

INVx5_ASAP7_75t_L g5033 ( 
.A(n_4831),
.Y(n_5033)
);

AOI22xp33_ASAP7_75t_SL g5034 ( 
.A1(n_4756),
.A2(n_180),
.B1(n_178),
.B2(n_179),
.Y(n_5034)
);

INVx1_ASAP7_75t_L g5035 ( 
.A(n_4869),
.Y(n_5035)
);

AOI22xp33_ASAP7_75t_L g5036 ( 
.A1(n_4723),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_5036)
);

BUFx2_ASAP7_75t_L g5037 ( 
.A(n_4714),
.Y(n_5037)
);

INVx2_ASAP7_75t_L g5038 ( 
.A(n_4756),
.Y(n_5038)
);

BUFx4f_ASAP7_75t_SL g5039 ( 
.A(n_4690),
.Y(n_5039)
);

AOI22xp33_ASAP7_75t_L g5040 ( 
.A1(n_4637),
.A2(n_184),
.B1(n_181),
.B2(n_182),
.Y(n_5040)
);

BUFx4_ASAP7_75t_R g5041 ( 
.A(n_4801),
.Y(n_5041)
);

INVxp67_ASAP7_75t_SL g5042 ( 
.A(n_4772),
.Y(n_5042)
);

INVx1_ASAP7_75t_L g5043 ( 
.A(n_4819),
.Y(n_5043)
);

AOI22xp33_ASAP7_75t_L g5044 ( 
.A1(n_4637),
.A2(n_185),
.B1(n_182),
.B2(n_184),
.Y(n_5044)
);

AOI22xp33_ASAP7_75t_SL g5045 ( 
.A1(n_4772),
.A2(n_187),
.B1(n_185),
.B2(n_186),
.Y(n_5045)
);

INVx1_ASAP7_75t_L g5046 ( 
.A(n_4821),
.Y(n_5046)
);

INVx2_ASAP7_75t_L g5047 ( 
.A(n_4833),
.Y(n_5047)
);

CKINVDCx20_ASAP7_75t_R g5048 ( 
.A(n_4753),
.Y(n_5048)
);

INVx2_ASAP7_75t_L g5049 ( 
.A(n_4839),
.Y(n_5049)
);

INVxp67_ASAP7_75t_SL g5050 ( 
.A(n_4823),
.Y(n_5050)
);

NAND2xp5_ASAP7_75t_L g5051 ( 
.A(n_4648),
.B(n_186),
.Y(n_5051)
);

BUFx2_ASAP7_75t_SL g5052 ( 
.A(n_4751),
.Y(n_5052)
);

AOI22xp33_ASAP7_75t_L g5053 ( 
.A1(n_4845),
.A2(n_191),
.B1(n_187),
.B2(n_189),
.Y(n_5053)
);

INVx1_ASAP7_75t_L g5054 ( 
.A(n_4826),
.Y(n_5054)
);

INVx6_ASAP7_75t_L g5055 ( 
.A(n_4748),
.Y(n_5055)
);

AOI22xp33_ASAP7_75t_L g5056 ( 
.A1(n_4800),
.A2(n_192),
.B1(n_189),
.B2(n_191),
.Y(n_5056)
);

INVx5_ASAP7_75t_L g5057 ( 
.A(n_4831),
.Y(n_5057)
);

AOI22xp33_ASAP7_75t_L g5058 ( 
.A1(n_4805),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.Y(n_5058)
);

INVx2_ASAP7_75t_L g5059 ( 
.A(n_4863),
.Y(n_5059)
);

NAND2xp5_ASAP7_75t_L g5060 ( 
.A(n_4633),
.B(n_194),
.Y(n_5060)
);

NAND2xp5_ASAP7_75t_L g5061 ( 
.A(n_4716),
.B(n_197),
.Y(n_5061)
);

INVx1_ASAP7_75t_L g5062 ( 
.A(n_4828),
.Y(n_5062)
);

INVx1_ASAP7_75t_L g5063 ( 
.A(n_4846),
.Y(n_5063)
);

AOI22xp33_ASAP7_75t_SL g5064 ( 
.A1(n_4810),
.A2(n_200),
.B1(n_198),
.B2(n_199),
.Y(n_5064)
);

OA21x2_ASAP7_75t_L g5065 ( 
.A1(n_4941),
.A2(n_4823),
.B(n_4791),
.Y(n_5065)
);

NAND2xp5_ASAP7_75t_L g5066 ( 
.A(n_4968),
.B(n_5008),
.Y(n_5066)
);

NOR2x1_ASAP7_75t_SL g5067 ( 
.A(n_5052),
.B(n_4983),
.Y(n_5067)
);

AOI21xp5_ASAP7_75t_L g5068 ( 
.A1(n_4901),
.A2(n_4859),
.B(n_4861),
.Y(n_5068)
);

INVx2_ASAP7_75t_L g5069 ( 
.A(n_4998),
.Y(n_5069)
);

AOI21xp5_ASAP7_75t_L g5070 ( 
.A1(n_4938),
.A2(n_4647),
.B(n_4816),
.Y(n_5070)
);

NAND2xp5_ASAP7_75t_L g5071 ( 
.A(n_5015),
.B(n_4727),
.Y(n_5071)
);

AOI21xp5_ASAP7_75t_L g5072 ( 
.A1(n_4875),
.A2(n_4837),
.B(n_4656),
.Y(n_5072)
);

OR2x2_ASAP7_75t_L g5073 ( 
.A(n_4936),
.B(n_4853),
.Y(n_5073)
);

AND2x2_ASAP7_75t_L g5074 ( 
.A(n_4974),
.B(n_4881),
.Y(n_5074)
);

AND2x4_ASAP7_75t_L g5075 ( 
.A(n_4946),
.B(n_4820),
.Y(n_5075)
);

AND2x4_ASAP7_75t_L g5076 ( 
.A(n_4946),
.B(n_4829),
.Y(n_5076)
);

HB1xp67_ASAP7_75t_L g5077 ( 
.A(n_4978),
.Y(n_5077)
);

HB1xp67_ASAP7_75t_L g5078 ( 
.A(n_5003),
.Y(n_5078)
);

INVx1_ASAP7_75t_L g5079 ( 
.A(n_4997),
.Y(n_5079)
);

NAND2xp5_ASAP7_75t_L g5080 ( 
.A(n_5018),
.B(n_4741),
.Y(n_5080)
);

CKINVDCx20_ASAP7_75t_R g5081 ( 
.A(n_4894),
.Y(n_5081)
);

OAI22xp5_ASAP7_75t_L g5082 ( 
.A1(n_5019),
.A2(n_4755),
.B1(n_4751),
.B2(n_4860),
.Y(n_5082)
);

AOI21xp5_ASAP7_75t_L g5083 ( 
.A1(n_4875),
.A2(n_4860),
.B(n_4742),
.Y(n_5083)
);

OR2x2_ASAP7_75t_L g5084 ( 
.A(n_4886),
.B(n_4864),
.Y(n_5084)
);

AND2x2_ASAP7_75t_L g5085 ( 
.A(n_4995),
.B(n_4808),
.Y(n_5085)
);

BUFx2_ASAP7_75t_L g5086 ( 
.A(n_5009),
.Y(n_5086)
);

OAI22xp5_ASAP7_75t_L g5087 ( 
.A1(n_4875),
.A2(n_4755),
.B1(n_4810),
.B2(n_4761),
.Y(n_5087)
);

INVx1_ASAP7_75t_L g5088 ( 
.A(n_4999),
.Y(n_5088)
);

OA21x2_ASAP7_75t_L g5089 ( 
.A1(n_5050),
.A2(n_4791),
.B(n_4813),
.Y(n_5089)
);

OR2x2_ASAP7_75t_L g5090 ( 
.A(n_4965),
.B(n_4815),
.Y(n_5090)
);

INVx1_ASAP7_75t_L g5091 ( 
.A(n_5001),
.Y(n_5091)
);

OAI22xp5_ASAP7_75t_L g5092 ( 
.A1(n_4983),
.A2(n_4766),
.B1(n_4834),
.B2(n_4740),
.Y(n_5092)
);

AOI221xp5_ASAP7_75t_L g5093 ( 
.A1(n_4975),
.A2(n_4985),
.B1(n_4953),
.B2(n_4993),
.C(n_4969),
.Y(n_5093)
);

O2A1O1Ixp5_ASAP7_75t_L g5094 ( 
.A1(n_4877),
.A2(n_4812),
.B(n_4844),
.C(n_4784),
.Y(n_5094)
);

AOI21xp5_ASAP7_75t_L g5095 ( 
.A1(n_5060),
.A2(n_4871),
.B(n_4707),
.Y(n_5095)
);

CKINVDCx5p33_ASAP7_75t_R g5096 ( 
.A(n_4884),
.Y(n_5096)
);

O2A1O1Ixp5_ASAP7_75t_L g5097 ( 
.A1(n_4888),
.A2(n_4959),
.B(n_5051),
.C(n_5007),
.Y(n_5097)
);

OAI22xp5_ASAP7_75t_L g5098 ( 
.A1(n_4983),
.A2(n_4834),
.B1(n_4775),
.B2(n_4636),
.Y(n_5098)
);

NAND3xp33_ASAP7_75t_L g5099 ( 
.A(n_4960),
.B(n_4752),
.C(n_4743),
.Y(n_5099)
);

O2A1O1Ixp33_ASAP7_75t_L g5100 ( 
.A1(n_4887),
.A2(n_4996),
.B(n_5030),
.C(n_5022),
.Y(n_5100)
);

AOI21xp5_ASAP7_75t_SL g5101 ( 
.A1(n_5042),
.A2(n_4760),
.B(n_4754),
.Y(n_5101)
);

AND2x2_ASAP7_75t_L g5102 ( 
.A(n_4883),
.B(n_4719),
.Y(n_5102)
);

AND2x2_ASAP7_75t_L g5103 ( 
.A(n_4922),
.B(n_4732),
.Y(n_5103)
);

OA21x2_ASAP7_75t_L g5104 ( 
.A1(n_5017),
.A2(n_4817),
.B(n_4872),
.Y(n_5104)
);

AND2x4_ASAP7_75t_L g5105 ( 
.A(n_5011),
.B(n_4829),
.Y(n_5105)
);

NOR2xp67_ASAP7_75t_L g5106 ( 
.A(n_5038),
.B(n_4649),
.Y(n_5106)
);

O2A1O1Ixp33_ASAP7_75t_L g5107 ( 
.A1(n_4927),
.A2(n_4849),
.B(n_4797),
.C(n_4804),
.Y(n_5107)
);

INVx1_ASAP7_75t_L g5108 ( 
.A(n_4895),
.Y(n_5108)
);

AOI21x1_ASAP7_75t_SL g5109 ( 
.A1(n_5061),
.A2(n_4793),
.B(n_4786),
.Y(n_5109)
);

HB1xp67_ASAP7_75t_L g5110 ( 
.A(n_5035),
.Y(n_5110)
);

NAND2xp5_ASAP7_75t_L g5111 ( 
.A(n_4896),
.B(n_4802),
.Y(n_5111)
);

OA21x2_ASAP7_75t_L g5112 ( 
.A1(n_5062),
.A2(n_4779),
.B(n_4776),
.Y(n_5112)
);

OAI22xp5_ASAP7_75t_L g5113 ( 
.A1(n_4977),
.A2(n_4811),
.B1(n_4649),
.B2(n_4807),
.Y(n_5113)
);

AOI21x1_ASAP7_75t_SL g5114 ( 
.A1(n_4984),
.A2(n_4806),
.B(n_4862),
.Y(n_5114)
);

OR2x6_ASAP7_75t_L g5115 ( 
.A(n_4956),
.B(n_4838),
.Y(n_5115)
);

HB1xp67_ASAP7_75t_L g5116 ( 
.A(n_4899),
.Y(n_5116)
);

HB1xp67_ASAP7_75t_L g5117 ( 
.A(n_4908),
.Y(n_5117)
);

NOR2xp67_ASAP7_75t_L g5118 ( 
.A(n_4874),
.B(n_4649),
.Y(n_5118)
);

OAI22xp5_ASAP7_75t_L g5119 ( 
.A1(n_4962),
.A2(n_4807),
.B1(n_4712),
.B2(n_4838),
.Y(n_5119)
);

AND2x2_ASAP7_75t_L g5120 ( 
.A(n_5004),
.B(n_4870),
.Y(n_5120)
);

AND2x2_ASAP7_75t_L g5121 ( 
.A(n_5010),
.B(n_5037),
.Y(n_5121)
);

AND2x4_ASAP7_75t_L g5122 ( 
.A(n_5029),
.B(n_4798),
.Y(n_5122)
);

AOI21x1_ASAP7_75t_SL g5123 ( 
.A1(n_5012),
.A2(n_199),
.B(n_200),
.Y(n_5123)
);

INVx3_ASAP7_75t_L g5124 ( 
.A(n_4987),
.Y(n_5124)
);

AOI21x1_ASAP7_75t_SL g5125 ( 
.A1(n_5020),
.A2(n_202),
.B(n_203),
.Y(n_5125)
);

A2O1A1Ixp33_ASAP7_75t_L g5126 ( 
.A1(n_4905),
.A2(n_4685),
.B(n_4768),
.C(n_4865),
.Y(n_5126)
);

O2A1O1Ixp33_ASAP7_75t_L g5127 ( 
.A1(n_4988),
.A2(n_4809),
.B(n_4868),
.C(n_4706),
.Y(n_5127)
);

HB1xp67_ASAP7_75t_L g5128 ( 
.A(n_4913),
.Y(n_5128)
);

OAI22xp5_ASAP7_75t_L g5129 ( 
.A1(n_4990),
.A2(n_4807),
.B1(n_4835),
.B2(n_4694),
.Y(n_5129)
);

OAI22xp5_ASAP7_75t_SL g5130 ( 
.A1(n_4954),
.A2(n_4685),
.B1(n_206),
.B2(n_203),
.Y(n_5130)
);

BUFx3_ASAP7_75t_L g5131 ( 
.A(n_4928),
.Y(n_5131)
);

INVx3_ASAP7_75t_L g5132 ( 
.A(n_4987),
.Y(n_5132)
);

BUFx2_ASAP7_75t_L g5133 ( 
.A(n_4906),
.Y(n_5133)
);

O2A1O1Ixp5_ASAP7_75t_L g5134 ( 
.A1(n_4970),
.A2(n_4747),
.B(n_4854),
.C(n_4818),
.Y(n_5134)
);

INVx1_ASAP7_75t_L g5135 ( 
.A(n_4921),
.Y(n_5135)
);

OAI22xp5_ASAP7_75t_L g5136 ( 
.A1(n_5016),
.A2(n_5045),
.B1(n_5034),
.B2(n_5028),
.Y(n_5136)
);

HB1xp67_ASAP7_75t_L g5137 ( 
.A(n_4930),
.Y(n_5137)
);

OAI22xp5_ASAP7_75t_L g5138 ( 
.A1(n_5021),
.A2(n_4696),
.B1(n_4827),
.B2(n_4803),
.Y(n_5138)
);

AOI21x1_ASAP7_75t_SL g5139 ( 
.A1(n_4893),
.A2(n_4919),
.B(n_4898),
.Y(n_5139)
);

AOI21xp5_ASAP7_75t_L g5140 ( 
.A1(n_4903),
.A2(n_4680),
.B(n_4758),
.Y(n_5140)
);

NOR2xp33_ASAP7_75t_L g5141 ( 
.A(n_4889),
.B(n_205),
.Y(n_5141)
);

OAI22xp5_ASAP7_75t_L g5142 ( 
.A1(n_4876),
.A2(n_4902),
.B1(n_5064),
.B2(n_5036),
.Y(n_5142)
);

AOI21xp5_ASAP7_75t_L g5143 ( 
.A1(n_4907),
.A2(n_4830),
.B(n_4795),
.Y(n_5143)
);

INVx1_ASAP7_75t_L g5144 ( 
.A(n_4931),
.Y(n_5144)
);

AOI21x1_ASAP7_75t_SL g5145 ( 
.A1(n_5041),
.A2(n_205),
.B(n_207),
.Y(n_5145)
);

AOI21xp5_ASAP7_75t_L g5146 ( 
.A1(n_4879),
.A2(n_4832),
.B(n_4847),
.Y(n_5146)
);

AND2x2_ASAP7_75t_L g5147 ( 
.A(n_5013),
.B(n_207),
.Y(n_5147)
);

INVx1_ASAP7_75t_L g5148 ( 
.A(n_4939),
.Y(n_5148)
);

AND2x4_ASAP7_75t_L g5149 ( 
.A(n_4873),
.B(n_208),
.Y(n_5149)
);

HB1xp67_ASAP7_75t_L g5150 ( 
.A(n_4940),
.Y(n_5150)
);

INVx1_ASAP7_75t_L g5151 ( 
.A(n_4955),
.Y(n_5151)
);

OAI22xp5_ASAP7_75t_SL g5152 ( 
.A1(n_4971),
.A2(n_211),
.B1(n_208),
.B2(n_209),
.Y(n_5152)
);

NAND2xp5_ASAP7_75t_L g5153 ( 
.A(n_4963),
.B(n_211),
.Y(n_5153)
);

OR2x2_ASAP7_75t_L g5154 ( 
.A(n_5002),
.B(n_212),
.Y(n_5154)
);

O2A1O1Ixp33_ASAP7_75t_L g5155 ( 
.A1(n_5014),
.A2(n_214),
.B(n_212),
.C(n_213),
.Y(n_5155)
);

OA22x2_ASAP7_75t_L g5156 ( 
.A1(n_4957),
.A2(n_4972),
.B1(n_5046),
.B2(n_5043),
.Y(n_5156)
);

AND2x2_ASAP7_75t_L g5157 ( 
.A(n_4979),
.B(n_213),
.Y(n_5157)
);

AOI21x1_ASAP7_75t_L g5158 ( 
.A1(n_5063),
.A2(n_214),
.B(n_215),
.Y(n_5158)
);

OAI22xp5_ASAP7_75t_L g5159 ( 
.A1(n_5023),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_5159)
);

AOI21xp5_ASAP7_75t_L g5160 ( 
.A1(n_4937),
.A2(n_217),
.B(n_220),
.Y(n_5160)
);

INVx1_ASAP7_75t_L g5161 ( 
.A(n_5054),
.Y(n_5161)
);

INVx1_ASAP7_75t_L g5162 ( 
.A(n_4981),
.Y(n_5162)
);

NAND2xp5_ASAP7_75t_L g5163 ( 
.A(n_4892),
.B(n_220),
.Y(n_5163)
);

NOR2xp33_ASAP7_75t_R g5164 ( 
.A(n_4909),
.B(n_221),
.Y(n_5164)
);

AOI221xp5_ASAP7_75t_L g5165 ( 
.A1(n_5053),
.A2(n_223),
.B1(n_221),
.B2(n_222),
.C(n_224),
.Y(n_5165)
);

CKINVDCx5p33_ASAP7_75t_R g5166 ( 
.A(n_4880),
.Y(n_5166)
);

INVx1_ASAP7_75t_L g5167 ( 
.A(n_4992),
.Y(n_5167)
);

CKINVDCx6p67_ASAP7_75t_R g5168 ( 
.A(n_4910),
.Y(n_5168)
);

O2A1O1Ixp5_ASAP7_75t_L g5169 ( 
.A1(n_4986),
.A2(n_5024),
.B(n_5059),
.C(n_4885),
.Y(n_5169)
);

OAI22xp5_ASAP7_75t_L g5170 ( 
.A1(n_5040),
.A2(n_228),
.B1(n_224),
.B2(n_227),
.Y(n_5170)
);

AOI21xp5_ASAP7_75t_SL g5171 ( 
.A1(n_4964),
.A2(n_227),
.B(n_228),
.Y(n_5171)
);

INVx2_ASAP7_75t_SL g5172 ( 
.A(n_4900),
.Y(n_5172)
);

NAND2xp5_ASAP7_75t_L g5173 ( 
.A(n_4892),
.B(n_229),
.Y(n_5173)
);

OR2x2_ASAP7_75t_SL g5174 ( 
.A(n_4900),
.B(n_229),
.Y(n_5174)
);

AOI21xp5_ASAP7_75t_SL g5175 ( 
.A1(n_5055),
.A2(n_230),
.B(n_231),
.Y(n_5175)
);

OAI22xp5_ASAP7_75t_L g5176 ( 
.A1(n_5044),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_5176)
);

O2A1O1Ixp5_ASAP7_75t_L g5177 ( 
.A1(n_4882),
.A2(n_234),
.B(n_232),
.C(n_233),
.Y(n_5177)
);

AOI21xp5_ASAP7_75t_L g5178 ( 
.A1(n_4878),
.A2(n_234),
.B(n_235),
.Y(n_5178)
);

OR2x2_ASAP7_75t_L g5179 ( 
.A(n_4917),
.B(n_235),
.Y(n_5179)
);

OR2x2_ASAP7_75t_L g5180 ( 
.A(n_4932),
.B(n_4942),
.Y(n_5180)
);

AND2x2_ASAP7_75t_L g5181 ( 
.A(n_4929),
.B(n_236),
.Y(n_5181)
);

AND2x4_ASAP7_75t_L g5182 ( 
.A(n_5033),
.B(n_236),
.Y(n_5182)
);

INVx1_ASAP7_75t_L g5183 ( 
.A(n_4952),
.Y(n_5183)
);

AOI21x1_ASAP7_75t_SL g5184 ( 
.A1(n_4944),
.A2(n_237),
.B(n_238),
.Y(n_5184)
);

NAND2xp5_ASAP7_75t_L g5185 ( 
.A(n_4892),
.B(n_239),
.Y(n_5185)
);

CKINVDCx5p33_ASAP7_75t_R g5186 ( 
.A(n_4967),
.Y(n_5186)
);

INVx1_ASAP7_75t_L g5187 ( 
.A(n_4961),
.Y(n_5187)
);

OR2x2_ASAP7_75t_L g5188 ( 
.A(n_4892),
.B(n_4956),
.Y(n_5188)
);

INVx1_ASAP7_75t_L g5189 ( 
.A(n_5047),
.Y(n_5189)
);

INVx2_ASAP7_75t_L g5190 ( 
.A(n_5049),
.Y(n_5190)
);

AND2x4_ASAP7_75t_L g5191 ( 
.A(n_5033),
.B(n_240),
.Y(n_5191)
);

AOI21xp5_ASAP7_75t_SL g5192 ( 
.A1(n_5055),
.A2(n_240),
.B(n_241),
.Y(n_5192)
);

AND2x2_ASAP7_75t_L g5193 ( 
.A(n_4914),
.B(n_241),
.Y(n_5193)
);

AND2x2_ASAP7_75t_L g5194 ( 
.A(n_4915),
.B(n_243),
.Y(n_5194)
);

NAND2xp5_ASAP7_75t_L g5195 ( 
.A(n_5006),
.B(n_243),
.Y(n_5195)
);

OR2x2_ASAP7_75t_L g5196 ( 
.A(n_4935),
.B(n_245),
.Y(n_5196)
);

INVx1_ASAP7_75t_L g5197 ( 
.A(n_4966),
.Y(n_5197)
);

AOI221xp5_ASAP7_75t_L g5198 ( 
.A1(n_5056),
.A2(n_247),
.B1(n_245),
.B2(n_246),
.C(n_248),
.Y(n_5198)
);

OA21x2_ASAP7_75t_L g5199 ( 
.A1(n_4923),
.A2(n_249),
.B(n_251),
.Y(n_5199)
);

OAI22xp5_ASAP7_75t_L g5200 ( 
.A1(n_5048),
.A2(n_254),
.B1(n_249),
.B2(n_252),
.Y(n_5200)
);

AOI21xp5_ASAP7_75t_L g5201 ( 
.A1(n_4904),
.A2(n_254),
.B(n_255),
.Y(n_5201)
);

AND2x2_ASAP7_75t_L g5202 ( 
.A(n_5032),
.B(n_255),
.Y(n_5202)
);

NAND2xp5_ASAP7_75t_L g5203 ( 
.A(n_5006),
.B(n_256),
.Y(n_5203)
);

INVx1_ASAP7_75t_L g5204 ( 
.A(n_4918),
.Y(n_5204)
);

AOI21xp5_ASAP7_75t_L g5205 ( 
.A1(n_4890),
.A2(n_257),
.B(n_258),
.Y(n_5205)
);

BUFx6f_ASAP7_75t_L g5206 ( 
.A(n_4874),
.Y(n_5206)
);

NAND2xp5_ASAP7_75t_L g5207 ( 
.A(n_4935),
.B(n_257),
.Y(n_5207)
);

AND2x2_ASAP7_75t_L g5208 ( 
.A(n_5025),
.B(n_260),
.Y(n_5208)
);

NOR2xp67_ASAP7_75t_L g5209 ( 
.A(n_4874),
.B(n_5033),
.Y(n_5209)
);

OA21x2_ASAP7_75t_L g5210 ( 
.A1(n_4925),
.A2(n_4911),
.B(n_4926),
.Y(n_5210)
);

AND2x2_ASAP7_75t_L g5211 ( 
.A(n_4973),
.B(n_260),
.Y(n_5211)
);

AND2x4_ASAP7_75t_L g5212 ( 
.A(n_5057),
.B(n_261),
.Y(n_5212)
);

A2O1A1Ixp33_ASAP7_75t_L g5213 ( 
.A1(n_4934),
.A2(n_265),
.B(n_263),
.C(n_264),
.Y(n_5213)
);

INVx2_ASAP7_75t_L g5214 ( 
.A(n_5104),
.Y(n_5214)
);

NOR2xp33_ASAP7_75t_R g5215 ( 
.A(n_5081),
.B(n_4976),
.Y(n_5215)
);

OR2x6_ASAP7_75t_L g5216 ( 
.A(n_5209),
.B(n_4912),
.Y(n_5216)
);

BUFx3_ASAP7_75t_L g5217 ( 
.A(n_5096),
.Y(n_5217)
);

NOR2x1_ASAP7_75t_L g5218 ( 
.A(n_5124),
.B(n_5132),
.Y(n_5218)
);

AND2x4_ASAP7_75t_L g5219 ( 
.A(n_5067),
.B(n_5057),
.Y(n_5219)
);

INVxp67_ASAP7_75t_SL g5220 ( 
.A(n_5077),
.Y(n_5220)
);

INVx1_ASAP7_75t_L g5221 ( 
.A(n_5117),
.Y(n_5221)
);

INVx4_ASAP7_75t_L g5222 ( 
.A(n_5166),
.Y(n_5222)
);

NAND2xp33_ASAP7_75t_R g5223 ( 
.A(n_5164),
.B(n_5186),
.Y(n_5223)
);

INVx1_ASAP7_75t_L g5224 ( 
.A(n_5128),
.Y(n_5224)
);

NAND2x1p5_ASAP7_75t_L g5225 ( 
.A(n_5118),
.B(n_5057),
.Y(n_5225)
);

INVx3_ASAP7_75t_L g5226 ( 
.A(n_5206),
.Y(n_5226)
);

NOR2xp33_ASAP7_75t_R g5227 ( 
.A(n_5133),
.B(n_5031),
.Y(n_5227)
);

AND2x4_ASAP7_75t_L g5228 ( 
.A(n_5074),
.B(n_4935),
.Y(n_5228)
);

NOR2xp33_ASAP7_75t_R g5229 ( 
.A(n_5086),
.B(n_4924),
.Y(n_5229)
);

OR2x2_ASAP7_75t_L g5230 ( 
.A(n_5066),
.B(n_4980),
.Y(n_5230)
);

AOI22xp33_ASAP7_75t_L g5231 ( 
.A1(n_5093),
.A2(n_4916),
.B1(n_4945),
.B2(n_4950),
.Y(n_5231)
);

AND2x2_ASAP7_75t_L g5232 ( 
.A(n_5121),
.B(n_4912),
.Y(n_5232)
);

INVx5_ASAP7_75t_L g5233 ( 
.A(n_5206),
.Y(n_5233)
);

BUFx3_ASAP7_75t_L g5234 ( 
.A(n_5131),
.Y(n_5234)
);

AND2x2_ASAP7_75t_L g5235 ( 
.A(n_5102),
.B(n_4889),
.Y(n_5235)
);

AND2x4_ASAP7_75t_L g5236 ( 
.A(n_5124),
.B(n_4980),
.Y(n_5236)
);

OAI21xp5_ASAP7_75t_L g5237 ( 
.A1(n_5097),
.A2(n_5058),
.B(n_5027),
.Y(n_5237)
);

AOI22xp33_ASAP7_75t_L g5238 ( 
.A1(n_5142),
.A2(n_4989),
.B1(n_4982),
.B2(n_4891),
.Y(n_5238)
);

INVx2_ASAP7_75t_L g5239 ( 
.A(n_5104),
.Y(n_5239)
);

AOI21xp5_ASAP7_75t_L g5240 ( 
.A1(n_5083),
.A2(n_5005),
.B(n_4994),
.Y(n_5240)
);

OA21x2_ASAP7_75t_L g5241 ( 
.A1(n_5204),
.A2(n_4947),
.B(n_5026),
.Y(n_5241)
);

AOI22xp33_ASAP7_75t_SL g5242 ( 
.A1(n_5210),
.A2(n_4948),
.B1(n_5000),
.B2(n_4982),
.Y(n_5242)
);

AND2x2_ASAP7_75t_L g5243 ( 
.A(n_5103),
.B(n_4980),
.Y(n_5243)
);

INVx1_ASAP7_75t_L g5244 ( 
.A(n_5137),
.Y(n_5244)
);

OR2x2_ASAP7_75t_L g5245 ( 
.A(n_5073),
.B(n_4991),
.Y(n_5245)
);

BUFx12f_ASAP7_75t_L g5246 ( 
.A(n_5206),
.Y(n_5246)
);

INVx1_ASAP7_75t_L g5247 ( 
.A(n_5150),
.Y(n_5247)
);

AND2x2_ASAP7_75t_L g5248 ( 
.A(n_5120),
.B(n_5085),
.Y(n_5248)
);

AOI21x1_ASAP7_75t_L g5249 ( 
.A1(n_5071),
.A2(n_5080),
.B(n_5098),
.Y(n_5249)
);

NOR2x1_ASAP7_75t_L g5250 ( 
.A(n_5132),
.B(n_4991),
.Y(n_5250)
);

NOR3xp33_ASAP7_75t_SL g5251 ( 
.A(n_5100),
.B(n_5039),
.C(n_4933),
.Y(n_5251)
);

AND2x4_ASAP7_75t_L g5252 ( 
.A(n_5122),
.B(n_4991),
.Y(n_5252)
);

BUFx3_ASAP7_75t_L g5253 ( 
.A(n_5168),
.Y(n_5253)
);

INVx1_ASAP7_75t_L g5254 ( 
.A(n_5161),
.Y(n_5254)
);

BUFx3_ASAP7_75t_L g5255 ( 
.A(n_5211),
.Y(n_5255)
);

XNOR2xp5_ASAP7_75t_L g5256 ( 
.A(n_5174),
.B(n_4924),
.Y(n_5256)
);

INVx1_ASAP7_75t_L g5257 ( 
.A(n_5079),
.Y(n_5257)
);

INVx2_ASAP7_75t_L g5258 ( 
.A(n_5084),
.Y(n_5258)
);

NAND2xp5_ASAP7_75t_L g5259 ( 
.A(n_5116),
.B(n_5000),
.Y(n_5259)
);

AO31x2_ASAP7_75t_L g5260 ( 
.A1(n_5068),
.A2(n_4943),
.A3(n_4933),
.B(n_4949),
.Y(n_5260)
);

INVx1_ASAP7_75t_L g5261 ( 
.A(n_5088),
.Y(n_5261)
);

INVxp67_ASAP7_75t_L g5262 ( 
.A(n_5078),
.Y(n_5262)
);

NAND2xp5_ASAP7_75t_L g5263 ( 
.A(n_5110),
.B(n_4948),
.Y(n_5263)
);

AND2x2_ASAP7_75t_L g5264 ( 
.A(n_5197),
.B(n_4951),
.Y(n_5264)
);

NAND2xp5_ASAP7_75t_L g5265 ( 
.A(n_5091),
.B(n_4920),
.Y(n_5265)
);

HB1xp67_ASAP7_75t_L g5266 ( 
.A(n_5108),
.Y(n_5266)
);

CKINVDCx20_ASAP7_75t_R g5267 ( 
.A(n_5172),
.Y(n_5267)
);

NOR2xp33_ASAP7_75t_R g5268 ( 
.A(n_5195),
.B(n_4943),
.Y(n_5268)
);

AOI22xp33_ASAP7_75t_SL g5269 ( 
.A1(n_5210),
.A2(n_4949),
.B1(n_4958),
.B2(n_4951),
.Y(n_5269)
);

AO21x2_ASAP7_75t_L g5270 ( 
.A1(n_5153),
.A2(n_4918),
.B(n_4897),
.Y(n_5270)
);

AND2x2_ASAP7_75t_L g5271 ( 
.A(n_5156),
.B(n_5188),
.Y(n_5271)
);

INVx2_ASAP7_75t_L g5272 ( 
.A(n_5069),
.Y(n_5272)
);

AND2x4_ASAP7_75t_L g5273 ( 
.A(n_5122),
.B(n_4958),
.Y(n_5273)
);

INVx1_ASAP7_75t_L g5274 ( 
.A(n_5135),
.Y(n_5274)
);

INVx1_ASAP7_75t_L g5275 ( 
.A(n_5144),
.Y(n_5275)
);

AND2x2_ASAP7_75t_L g5276 ( 
.A(n_5075),
.B(n_263),
.Y(n_5276)
);

INVx2_ASAP7_75t_L g5277 ( 
.A(n_5180),
.Y(n_5277)
);

NAND2xp5_ASAP7_75t_L g5278 ( 
.A(n_5148),
.B(n_264),
.Y(n_5278)
);

INVx1_ASAP7_75t_L g5279 ( 
.A(n_5151),
.Y(n_5279)
);

CKINVDCx5p33_ASAP7_75t_R g5280 ( 
.A(n_5181),
.Y(n_5280)
);

NAND3xp33_ASAP7_75t_SL g5281 ( 
.A(n_5169),
.B(n_265),
.C(n_267),
.Y(n_5281)
);

BUFx10_ASAP7_75t_L g5282 ( 
.A(n_5182),
.Y(n_5282)
);

AND2x2_ASAP7_75t_L g5283 ( 
.A(n_5075),
.B(n_268),
.Y(n_5283)
);

INVx4_ASAP7_75t_L g5284 ( 
.A(n_5149),
.Y(n_5284)
);

CKINVDCx5p33_ASAP7_75t_R g5285 ( 
.A(n_5157),
.Y(n_5285)
);

NAND2xp33_ASAP7_75t_R g5286 ( 
.A(n_5182),
.B(n_5191),
.Y(n_5286)
);

CKINVDCx5p33_ASAP7_75t_R g5287 ( 
.A(n_5203),
.Y(n_5287)
);

BUFx10_ASAP7_75t_L g5288 ( 
.A(n_5191),
.Y(n_5288)
);

AO21x2_ASAP7_75t_L g5289 ( 
.A1(n_5163),
.A2(n_268),
.B(n_270),
.Y(n_5289)
);

CKINVDCx5p33_ASAP7_75t_R g5290 ( 
.A(n_5208),
.Y(n_5290)
);

OAI22xp5_ASAP7_75t_SL g5291 ( 
.A1(n_5152),
.A2(n_274),
.B1(n_271),
.B2(n_273),
.Y(n_5291)
);

AND2x2_ASAP7_75t_L g5292 ( 
.A(n_5076),
.B(n_275),
.Y(n_5292)
);

OR2x6_ASAP7_75t_L g5293 ( 
.A(n_5212),
.B(n_277),
.Y(n_5293)
);

OR2x2_ASAP7_75t_L g5294 ( 
.A(n_5111),
.B(n_5090),
.Y(n_5294)
);

CKINVDCx16_ASAP7_75t_R g5295 ( 
.A(n_5115),
.Y(n_5295)
);

INVxp67_ASAP7_75t_L g5296 ( 
.A(n_5141),
.Y(n_5296)
);

AND2x4_ASAP7_75t_L g5297 ( 
.A(n_5076),
.B(n_278),
.Y(n_5297)
);

NOR2xp33_ASAP7_75t_L g5298 ( 
.A(n_5149),
.B(n_278),
.Y(n_5298)
);

AND2x4_ASAP7_75t_L g5299 ( 
.A(n_5115),
.B(n_5212),
.Y(n_5299)
);

AOI22xp33_ASAP7_75t_L g5300 ( 
.A1(n_5099),
.A2(n_282),
.B1(n_279),
.B2(n_280),
.Y(n_5300)
);

BUFx3_ASAP7_75t_L g5301 ( 
.A(n_5147),
.Y(n_5301)
);

AOI22xp33_ASAP7_75t_L g5302 ( 
.A1(n_5199),
.A2(n_5136),
.B1(n_5070),
.B2(n_5072),
.Y(n_5302)
);

NAND2xp33_ASAP7_75t_R g5303 ( 
.A(n_5193),
.B(n_5194),
.Y(n_5303)
);

AOI22xp33_ASAP7_75t_L g5304 ( 
.A1(n_5199),
.A2(n_283),
.B1(n_279),
.B2(n_282),
.Y(n_5304)
);

AND2x2_ASAP7_75t_L g5305 ( 
.A(n_5105),
.B(n_284),
.Y(n_5305)
);

NOR2xp33_ASAP7_75t_L g5306 ( 
.A(n_5130),
.B(n_285),
.Y(n_5306)
);

O2A1O1Ixp33_ASAP7_75t_SL g5307 ( 
.A1(n_5159),
.A2(n_289),
.B(n_287),
.C(n_288),
.Y(n_5307)
);

BUFx2_ASAP7_75t_L g5308 ( 
.A(n_5065),
.Y(n_5308)
);

OAI22xp5_ASAP7_75t_L g5309 ( 
.A1(n_5082),
.A2(n_292),
.B1(n_289),
.B2(n_291),
.Y(n_5309)
);

AOI22xp5_ASAP7_75t_L g5310 ( 
.A1(n_5119),
.A2(n_295),
.B1(n_292),
.B2(n_293),
.Y(n_5310)
);

INVx1_ASAP7_75t_L g5311 ( 
.A(n_5162),
.Y(n_5311)
);

NOR2xp33_ASAP7_75t_L g5312 ( 
.A(n_5154),
.B(n_293),
.Y(n_5312)
);

AO31x2_ASAP7_75t_L g5313 ( 
.A1(n_5087),
.A2(n_301),
.A3(n_296),
.B(n_297),
.Y(n_5313)
);

OR2x2_ASAP7_75t_L g5314 ( 
.A(n_5167),
.B(n_296),
.Y(n_5314)
);

CKINVDCx5p33_ASAP7_75t_R g5315 ( 
.A(n_5202),
.Y(n_5315)
);

OR2x6_ASAP7_75t_L g5316 ( 
.A(n_5175),
.B(n_302),
.Y(n_5316)
);

INVx1_ASAP7_75t_L g5317 ( 
.A(n_5179),
.Y(n_5317)
);

AND2x4_ASAP7_75t_SL g5318 ( 
.A(n_5105),
.B(n_303),
.Y(n_5318)
);

NAND2xp5_ASAP7_75t_L g5319 ( 
.A(n_5095),
.B(n_305),
.Y(n_5319)
);

INVx2_ASAP7_75t_L g5320 ( 
.A(n_5190),
.Y(n_5320)
);

INVx1_ASAP7_75t_L g5321 ( 
.A(n_5183),
.Y(n_5321)
);

AND2x4_ASAP7_75t_L g5322 ( 
.A(n_5106),
.B(n_305),
.Y(n_5322)
);

OR2x6_ASAP7_75t_L g5323 ( 
.A(n_5192),
.B(n_307),
.Y(n_5323)
);

NOR2x1p5_ASAP7_75t_L g5324 ( 
.A(n_5173),
.B(n_307),
.Y(n_5324)
);

INVx1_ASAP7_75t_L g5325 ( 
.A(n_5187),
.Y(n_5325)
);

CKINVDCx5p33_ASAP7_75t_R g5326 ( 
.A(n_5092),
.Y(n_5326)
);

NOR3xp33_ASAP7_75t_SL g5327 ( 
.A(n_5200),
.B(n_308),
.C(n_309),
.Y(n_5327)
);

INVx2_ASAP7_75t_SL g5328 ( 
.A(n_5196),
.Y(n_5328)
);

OAI22xp5_ASAP7_75t_L g5329 ( 
.A1(n_5185),
.A2(n_310),
.B1(n_308),
.B2(n_309),
.Y(n_5329)
);

AND2x2_ASAP7_75t_L g5330 ( 
.A(n_5101),
.B(n_312),
.Y(n_5330)
);

AND2x2_ASAP7_75t_L g5331 ( 
.A(n_5094),
.B(n_5065),
.Y(n_5331)
);

AND2x4_ASAP7_75t_L g5332 ( 
.A(n_5143),
.B(n_312),
.Y(n_5332)
);

NOR2xp33_ASAP7_75t_R g5333 ( 
.A(n_5158),
.B(n_313),
.Y(n_5333)
);

NAND2xp33_ASAP7_75t_R g5334 ( 
.A(n_5089),
.B(n_313),
.Y(n_5334)
);

BUFx10_ASAP7_75t_L g5335 ( 
.A(n_5171),
.Y(n_5335)
);

CKINVDCx5p33_ASAP7_75t_R g5336 ( 
.A(n_5207),
.Y(n_5336)
);

NOR3xp33_ASAP7_75t_SL g5337 ( 
.A(n_5178),
.B(n_314),
.C(n_316),
.Y(n_5337)
);

AOI22xp33_ASAP7_75t_SL g5338 ( 
.A1(n_5113),
.A2(n_317),
.B1(n_314),
.B2(n_316),
.Y(n_5338)
);

NOR3xp33_ASAP7_75t_SL g5339 ( 
.A(n_5201),
.B(n_318),
.C(n_319),
.Y(n_5339)
);

INVx2_ASAP7_75t_L g5340 ( 
.A(n_5089),
.Y(n_5340)
);

CKINVDCx5p33_ASAP7_75t_R g5341 ( 
.A(n_5129),
.Y(n_5341)
);

INVx1_ASAP7_75t_L g5342 ( 
.A(n_5189),
.Y(n_5342)
);

AO31x2_ASAP7_75t_L g5343 ( 
.A1(n_5126),
.A2(n_320),
.A3(n_318),
.B(n_319),
.Y(n_5343)
);

INVx1_ASAP7_75t_L g5344 ( 
.A(n_5127),
.Y(n_5344)
);

HB1xp67_ASAP7_75t_L g5345 ( 
.A(n_5138),
.Y(n_5345)
);

NAND2xp33_ASAP7_75t_R g5346 ( 
.A(n_5112),
.B(n_5145),
.Y(n_5346)
);

AND2x2_ASAP7_75t_L g5347 ( 
.A(n_5139),
.B(n_320),
.Y(n_5347)
);

INVx1_ASAP7_75t_L g5348 ( 
.A(n_5107),
.Y(n_5348)
);

AND2x2_ASAP7_75t_L g5349 ( 
.A(n_5146),
.B(n_321),
.Y(n_5349)
);

OR2x6_ASAP7_75t_L g5350 ( 
.A(n_5205),
.B(n_5140),
.Y(n_5350)
);

AOI22xp5_ASAP7_75t_L g5351 ( 
.A1(n_5170),
.A2(n_324),
.B1(n_322),
.B2(n_323),
.Y(n_5351)
);

INVx2_ASAP7_75t_SL g5352 ( 
.A(n_5109),
.Y(n_5352)
);

BUFx4f_ASAP7_75t_SL g5353 ( 
.A(n_5184),
.Y(n_5353)
);

HB1xp67_ASAP7_75t_L g5354 ( 
.A(n_5160),
.Y(n_5354)
);

OAI22xp5_ASAP7_75t_L g5355 ( 
.A1(n_5165),
.A2(n_326),
.B1(n_324),
.B2(n_325),
.Y(n_5355)
);

NOR3xp33_ASAP7_75t_SL g5356 ( 
.A(n_5155),
.B(n_325),
.C(n_327),
.Y(n_5356)
);

INVx2_ASAP7_75t_L g5357 ( 
.A(n_5214),
.Y(n_5357)
);

OR2x2_ASAP7_75t_L g5358 ( 
.A(n_5221),
.B(n_5112),
.Y(n_5358)
);

BUFx6f_ASAP7_75t_L g5359 ( 
.A(n_5319),
.Y(n_5359)
);

AND2x2_ASAP7_75t_L g5360 ( 
.A(n_5271),
.B(n_5134),
.Y(n_5360)
);

INVx1_ASAP7_75t_L g5361 ( 
.A(n_5266),
.Y(n_5361)
);

INVx3_ASAP7_75t_L g5362 ( 
.A(n_5219),
.Y(n_5362)
);

AOI22xp5_ASAP7_75t_L g5363 ( 
.A1(n_5334),
.A2(n_5302),
.B1(n_5346),
.B2(n_5281),
.Y(n_5363)
);

NAND2xp5_ASAP7_75t_L g5364 ( 
.A(n_5345),
.B(n_5213),
.Y(n_5364)
);

AOI22xp33_ASAP7_75t_L g5365 ( 
.A1(n_5348),
.A2(n_5198),
.B1(n_5176),
.B2(n_5125),
.Y(n_5365)
);

BUFx6f_ASAP7_75t_L g5366 ( 
.A(n_5217),
.Y(n_5366)
);

AOI21x1_ASAP7_75t_L g5367 ( 
.A1(n_5308),
.A2(n_5114),
.B(n_5123),
.Y(n_5367)
);

AND2x2_ASAP7_75t_L g5368 ( 
.A(n_5248),
.B(n_5177),
.Y(n_5368)
);

AND2x4_ASAP7_75t_L g5369 ( 
.A(n_5219),
.B(n_328),
.Y(n_5369)
);

AND2x2_ASAP7_75t_L g5370 ( 
.A(n_5218),
.B(n_329),
.Y(n_5370)
);

INVx1_ASAP7_75t_L g5371 ( 
.A(n_5254),
.Y(n_5371)
);

NAND2xp5_ASAP7_75t_L g5372 ( 
.A(n_5344),
.B(n_329),
.Y(n_5372)
);

BUFx3_ASAP7_75t_L g5373 ( 
.A(n_5253),
.Y(n_5373)
);

INVx1_ASAP7_75t_L g5374 ( 
.A(n_5257),
.Y(n_5374)
);

INVx4_ASAP7_75t_L g5375 ( 
.A(n_5233),
.Y(n_5375)
);

AND2x2_ASAP7_75t_L g5376 ( 
.A(n_5232),
.B(n_330),
.Y(n_5376)
);

INVx1_ASAP7_75t_L g5377 ( 
.A(n_5261),
.Y(n_5377)
);

AND2x2_ASAP7_75t_L g5378 ( 
.A(n_5235),
.B(n_5243),
.Y(n_5378)
);

INVx1_ASAP7_75t_L g5379 ( 
.A(n_5274),
.Y(n_5379)
);

AO21x2_ASAP7_75t_L g5380 ( 
.A1(n_5331),
.A2(n_330),
.B(n_331),
.Y(n_5380)
);

AND2x2_ASAP7_75t_L g5381 ( 
.A(n_5284),
.B(n_5228),
.Y(n_5381)
);

INVx2_ASAP7_75t_L g5382 ( 
.A(n_5239),
.Y(n_5382)
);

AND2x2_ASAP7_75t_L g5383 ( 
.A(n_5228),
.B(n_332),
.Y(n_5383)
);

OR2x2_ASAP7_75t_L g5384 ( 
.A(n_5224),
.B(n_333),
.Y(n_5384)
);

AO21x2_ASAP7_75t_L g5385 ( 
.A1(n_5340),
.A2(n_334),
.B(n_336),
.Y(n_5385)
);

OR2x6_ASAP7_75t_L g5386 ( 
.A(n_5216),
.B(n_337),
.Y(n_5386)
);

OA21x2_ASAP7_75t_L g5387 ( 
.A1(n_5308),
.A2(n_337),
.B(n_338),
.Y(n_5387)
);

INVx1_ASAP7_75t_L g5388 ( 
.A(n_5275),
.Y(n_5388)
);

AOI22xp33_ASAP7_75t_L g5389 ( 
.A1(n_5354),
.A2(n_342),
.B1(n_338),
.B2(n_341),
.Y(n_5389)
);

INVx2_ASAP7_75t_L g5390 ( 
.A(n_5289),
.Y(n_5390)
);

INVx2_ASAP7_75t_L g5391 ( 
.A(n_5294),
.Y(n_5391)
);

OAI221xp5_ASAP7_75t_L g5392 ( 
.A1(n_5269),
.A2(n_345),
.B1(n_343),
.B2(n_344),
.C(n_346),
.Y(n_5392)
);

INVx1_ASAP7_75t_L g5393 ( 
.A(n_5279),
.Y(n_5393)
);

INVx1_ASAP7_75t_L g5394 ( 
.A(n_5244),
.Y(n_5394)
);

AND2x2_ASAP7_75t_L g5395 ( 
.A(n_5236),
.B(n_344),
.Y(n_5395)
);

NAND2xp5_ASAP7_75t_L g5396 ( 
.A(n_5332),
.B(n_5262),
.Y(n_5396)
);

HB1xp67_ASAP7_75t_L g5397 ( 
.A(n_5265),
.Y(n_5397)
);

INVx1_ASAP7_75t_L g5398 ( 
.A(n_5247),
.Y(n_5398)
);

NAND2xp5_ASAP7_75t_L g5399 ( 
.A(n_5332),
.B(n_347),
.Y(n_5399)
);

HB1xp67_ASAP7_75t_L g5400 ( 
.A(n_5270),
.Y(n_5400)
);

AO21x2_ASAP7_75t_L g5401 ( 
.A1(n_5278),
.A2(n_347),
.B(n_348),
.Y(n_5401)
);

NAND2xp5_ASAP7_75t_L g5402 ( 
.A(n_5220),
.B(n_348),
.Y(n_5402)
);

INVx1_ASAP7_75t_L g5403 ( 
.A(n_5311),
.Y(n_5403)
);

INVx2_ASAP7_75t_SL g5404 ( 
.A(n_5282),
.Y(n_5404)
);

INVx1_ASAP7_75t_L g5405 ( 
.A(n_5321),
.Y(n_5405)
);

NAND2xp5_ASAP7_75t_L g5406 ( 
.A(n_5349),
.B(n_350),
.Y(n_5406)
);

HB1xp67_ASAP7_75t_L g5407 ( 
.A(n_5350),
.Y(n_5407)
);

AND2x2_ASAP7_75t_L g5408 ( 
.A(n_5236),
.B(n_351),
.Y(n_5408)
);

OA21x2_ASAP7_75t_L g5409 ( 
.A1(n_5237),
.A2(n_351),
.B(n_352),
.Y(n_5409)
);

INVx2_ASAP7_75t_L g5410 ( 
.A(n_5272),
.Y(n_5410)
);

INVx1_ASAP7_75t_L g5411 ( 
.A(n_5325),
.Y(n_5411)
);

NOR2xp33_ASAP7_75t_SL g5412 ( 
.A(n_5222),
.B(n_353),
.Y(n_5412)
);

INVx1_ASAP7_75t_L g5413 ( 
.A(n_5342),
.Y(n_5413)
);

INVx1_ASAP7_75t_L g5414 ( 
.A(n_5317),
.Y(n_5414)
);

OR2x6_ASAP7_75t_L g5415 ( 
.A(n_5216),
.B(n_354),
.Y(n_5415)
);

INVxp67_ASAP7_75t_L g5416 ( 
.A(n_5350),
.Y(n_5416)
);

HB1xp67_ASAP7_75t_L g5417 ( 
.A(n_5352),
.Y(n_5417)
);

INVx1_ASAP7_75t_L g5418 ( 
.A(n_5314),
.Y(n_5418)
);

NOR2x1_ASAP7_75t_L g5419 ( 
.A(n_5293),
.B(n_354),
.Y(n_5419)
);

NOR2xp33_ASAP7_75t_SL g5420 ( 
.A(n_5295),
.B(n_355),
.Y(n_5420)
);

INVx1_ASAP7_75t_L g5421 ( 
.A(n_5258),
.Y(n_5421)
);

OAI21xp33_ASAP7_75t_L g5422 ( 
.A1(n_5306),
.A2(n_356),
.B(n_357),
.Y(n_5422)
);

BUFx3_ASAP7_75t_L g5423 ( 
.A(n_5255),
.Y(n_5423)
);

AO21x2_ASAP7_75t_L g5424 ( 
.A1(n_5249),
.A2(n_356),
.B(n_357),
.Y(n_5424)
);

INVx2_ASAP7_75t_L g5425 ( 
.A(n_5277),
.Y(n_5425)
);

OAI21xp5_ASAP7_75t_SL g5426 ( 
.A1(n_5242),
.A2(n_361),
.B(n_362),
.Y(n_5426)
);

OR2x2_ASAP7_75t_L g5427 ( 
.A(n_5230),
.B(n_361),
.Y(n_5427)
);

AND2x4_ASAP7_75t_L g5428 ( 
.A(n_5299),
.B(n_362),
.Y(n_5428)
);

INVx2_ASAP7_75t_L g5429 ( 
.A(n_5313),
.Y(n_5429)
);

INVx3_ASAP7_75t_L g5430 ( 
.A(n_5260),
.Y(n_5430)
);

AND2x4_ASAP7_75t_L g5431 ( 
.A(n_5299),
.B(n_363),
.Y(n_5431)
);

INVx2_ASAP7_75t_L g5432 ( 
.A(n_5313),
.Y(n_5432)
);

BUFx2_ASAP7_75t_L g5433 ( 
.A(n_5227),
.Y(n_5433)
);

NAND2xp5_ASAP7_75t_L g5434 ( 
.A(n_5330),
.B(n_363),
.Y(n_5434)
);

AO21x2_ASAP7_75t_L g5435 ( 
.A1(n_5333),
.A2(n_365),
.B(n_366),
.Y(n_5435)
);

OAI21x1_ASAP7_75t_L g5436 ( 
.A1(n_5250),
.A2(n_5259),
.B(n_5263),
.Y(n_5436)
);

AND2x2_ASAP7_75t_L g5437 ( 
.A(n_5226),
.B(n_365),
.Y(n_5437)
);

INVx1_ASAP7_75t_L g5438 ( 
.A(n_5328),
.Y(n_5438)
);

AOI22xp33_ASAP7_75t_L g5439 ( 
.A1(n_5291),
.A2(n_368),
.B1(n_366),
.B2(n_367),
.Y(n_5439)
);

INVx2_ASAP7_75t_L g5440 ( 
.A(n_5320),
.Y(n_5440)
);

AO21x2_ASAP7_75t_L g5441 ( 
.A1(n_5312),
.A2(n_5310),
.B(n_5347),
.Y(n_5441)
);

INVx2_ASAP7_75t_L g5442 ( 
.A(n_5343),
.Y(n_5442)
);

INVx1_ASAP7_75t_L g5443 ( 
.A(n_5245),
.Y(n_5443)
);

INVx2_ASAP7_75t_L g5444 ( 
.A(n_5343),
.Y(n_5444)
);

INVxp67_ASAP7_75t_SL g5445 ( 
.A(n_5324),
.Y(n_5445)
);

AND2x2_ASAP7_75t_L g5446 ( 
.A(n_5264),
.B(n_367),
.Y(n_5446)
);

INVx1_ASAP7_75t_L g5447 ( 
.A(n_5301),
.Y(n_5447)
);

INVx1_ASAP7_75t_L g5448 ( 
.A(n_5305),
.Y(n_5448)
);

INVx2_ASAP7_75t_L g5449 ( 
.A(n_5293),
.Y(n_5449)
);

AND2x2_ASAP7_75t_L g5450 ( 
.A(n_5233),
.B(n_369),
.Y(n_5450)
);

AO21x2_ASAP7_75t_L g5451 ( 
.A1(n_5329),
.A2(n_369),
.B(n_370),
.Y(n_5451)
);

INVx2_ASAP7_75t_SL g5452 ( 
.A(n_5288),
.Y(n_5452)
);

INVx2_ASAP7_75t_L g5453 ( 
.A(n_5241),
.Y(n_5453)
);

AND2x2_ASAP7_75t_L g5454 ( 
.A(n_5233),
.B(n_370),
.Y(n_5454)
);

OA21x2_ASAP7_75t_L g5455 ( 
.A1(n_5341),
.A2(n_371),
.B(n_372),
.Y(n_5455)
);

AND2x2_ASAP7_75t_L g5456 ( 
.A(n_5273),
.B(n_374),
.Y(n_5456)
);

INVx2_ASAP7_75t_L g5457 ( 
.A(n_5241),
.Y(n_5457)
);

NAND2xp5_ASAP7_75t_L g5458 ( 
.A(n_5326),
.B(n_374),
.Y(n_5458)
);

AND2x2_ASAP7_75t_L g5459 ( 
.A(n_5273),
.B(n_375),
.Y(n_5459)
);

INVx1_ASAP7_75t_L g5460 ( 
.A(n_5336),
.Y(n_5460)
);

AND2x2_ASAP7_75t_L g5461 ( 
.A(n_5252),
.B(n_376),
.Y(n_5461)
);

AND2x2_ASAP7_75t_L g5462 ( 
.A(n_5252),
.B(n_377),
.Y(n_5462)
);

INVx2_ASAP7_75t_L g5463 ( 
.A(n_5335),
.Y(n_5463)
);

HB1xp67_ASAP7_75t_L g5464 ( 
.A(n_5286),
.Y(n_5464)
);

BUFx3_ASAP7_75t_L g5465 ( 
.A(n_5246),
.Y(n_5465)
);

INVxp67_ASAP7_75t_SL g5466 ( 
.A(n_5300),
.Y(n_5466)
);

AND2x2_ASAP7_75t_L g5467 ( 
.A(n_5407),
.B(n_5260),
.Y(n_5467)
);

NOR2xp33_ASAP7_75t_L g5468 ( 
.A(n_5433),
.B(n_5256),
.Y(n_5468)
);

INVx2_ASAP7_75t_L g5469 ( 
.A(n_5387),
.Y(n_5469)
);

INVx1_ASAP7_75t_L g5470 ( 
.A(n_5371),
.Y(n_5470)
);

INVx1_ASAP7_75t_L g5471 ( 
.A(n_5374),
.Y(n_5471)
);

INVx1_ASAP7_75t_L g5472 ( 
.A(n_5377),
.Y(n_5472)
);

INVx5_ASAP7_75t_L g5473 ( 
.A(n_5375),
.Y(n_5473)
);

HB1xp67_ASAP7_75t_L g5474 ( 
.A(n_5387),
.Y(n_5474)
);

OR2x2_ASAP7_75t_L g5475 ( 
.A(n_5391),
.B(n_5238),
.Y(n_5475)
);

AND2x2_ASAP7_75t_L g5476 ( 
.A(n_5407),
.B(n_5251),
.Y(n_5476)
);

INVx1_ASAP7_75t_L g5477 ( 
.A(n_5379),
.Y(n_5477)
);

INVx2_ASAP7_75t_SL g5478 ( 
.A(n_5373),
.Y(n_5478)
);

NAND2xp5_ASAP7_75t_L g5479 ( 
.A(n_5359),
.B(n_5298),
.Y(n_5479)
);

AND2x2_ASAP7_75t_L g5480 ( 
.A(n_5423),
.B(n_5234),
.Y(n_5480)
);

INVx1_ASAP7_75t_L g5481 ( 
.A(n_5388),
.Y(n_5481)
);

OR2x2_ASAP7_75t_L g5482 ( 
.A(n_5391),
.B(n_5309),
.Y(n_5482)
);

OR2x2_ASAP7_75t_L g5483 ( 
.A(n_5414),
.B(n_5296),
.Y(n_5483)
);

NAND2xp5_ASAP7_75t_L g5484 ( 
.A(n_5359),
.B(n_5297),
.Y(n_5484)
);

INVx2_ASAP7_75t_L g5485 ( 
.A(n_5387),
.Y(n_5485)
);

OR2x2_ASAP7_75t_L g5486 ( 
.A(n_5361),
.B(n_5438),
.Y(n_5486)
);

NAND2xp5_ASAP7_75t_L g5487 ( 
.A(n_5359),
.B(n_5297),
.Y(n_5487)
);

INVx2_ASAP7_75t_L g5488 ( 
.A(n_5455),
.Y(n_5488)
);

AND2x2_ASAP7_75t_L g5489 ( 
.A(n_5362),
.B(n_5229),
.Y(n_5489)
);

AND2x2_ASAP7_75t_L g5490 ( 
.A(n_5362),
.B(n_5280),
.Y(n_5490)
);

INVx2_ASAP7_75t_L g5491 ( 
.A(n_5455),
.Y(n_5491)
);

INVx2_ASAP7_75t_L g5492 ( 
.A(n_5455),
.Y(n_5492)
);

AND2x2_ASAP7_75t_L g5493 ( 
.A(n_5417),
.B(n_5285),
.Y(n_5493)
);

INVx2_ASAP7_75t_L g5494 ( 
.A(n_5424),
.Y(n_5494)
);

NOR2x1_ASAP7_75t_L g5495 ( 
.A(n_5386),
.B(n_5276),
.Y(n_5495)
);

INVx1_ASAP7_75t_L g5496 ( 
.A(n_5393),
.Y(n_5496)
);

INVx1_ASAP7_75t_L g5497 ( 
.A(n_5403),
.Y(n_5497)
);

INVx1_ASAP7_75t_L g5498 ( 
.A(n_5405),
.Y(n_5498)
);

AND2x2_ASAP7_75t_L g5499 ( 
.A(n_5417),
.B(n_5267),
.Y(n_5499)
);

AND2x2_ASAP7_75t_L g5500 ( 
.A(n_5360),
.B(n_5268),
.Y(n_5500)
);

BUFx2_ASAP7_75t_L g5501 ( 
.A(n_5373),
.Y(n_5501)
);

AOI22xp33_ASAP7_75t_L g5502 ( 
.A1(n_5359),
.A2(n_5353),
.B1(n_5304),
.B2(n_5355),
.Y(n_5502)
);

BUFx3_ASAP7_75t_L g5503 ( 
.A(n_5366),
.Y(n_5503)
);

NAND2xp5_ASAP7_75t_L g5504 ( 
.A(n_5364),
.B(n_5368),
.Y(n_5504)
);

NOR3xp33_ASAP7_75t_L g5505 ( 
.A(n_5430),
.B(n_5338),
.C(n_5307),
.Y(n_5505)
);

INVx3_ASAP7_75t_L g5506 ( 
.A(n_5375),
.Y(n_5506)
);

NOR2xp33_ASAP7_75t_L g5507 ( 
.A(n_5366),
.B(n_5287),
.Y(n_5507)
);

HB1xp67_ASAP7_75t_L g5508 ( 
.A(n_5380),
.Y(n_5508)
);

AND2x2_ASAP7_75t_L g5509 ( 
.A(n_5423),
.B(n_5215),
.Y(n_5509)
);

AND2x2_ASAP7_75t_L g5510 ( 
.A(n_5378),
.B(n_5283),
.Y(n_5510)
);

OR2x2_ASAP7_75t_L g5511 ( 
.A(n_5394),
.B(n_5231),
.Y(n_5511)
);

AND2x2_ASAP7_75t_L g5512 ( 
.A(n_5381),
.B(n_5292),
.Y(n_5512)
);

OAI22xp5_ASAP7_75t_L g5513 ( 
.A1(n_5363),
.A2(n_5464),
.B1(n_5416),
.B2(n_5426),
.Y(n_5513)
);

INVx1_ASAP7_75t_L g5514 ( 
.A(n_5411),
.Y(n_5514)
);

INVx2_ASAP7_75t_L g5515 ( 
.A(n_5424),
.Y(n_5515)
);

AND2x2_ASAP7_75t_L g5516 ( 
.A(n_5404),
.B(n_5315),
.Y(n_5516)
);

INVx2_ASAP7_75t_L g5517 ( 
.A(n_5409),
.Y(n_5517)
);

INVx1_ASAP7_75t_L g5518 ( 
.A(n_5413),
.Y(n_5518)
);

AND2x2_ASAP7_75t_L g5519 ( 
.A(n_5375),
.B(n_5225),
.Y(n_5519)
);

INVx1_ASAP7_75t_L g5520 ( 
.A(n_5398),
.Y(n_5520)
);

INVx2_ASAP7_75t_SL g5521 ( 
.A(n_5366),
.Y(n_5521)
);

OAI221xp5_ASAP7_75t_L g5522 ( 
.A1(n_5464),
.A2(n_5397),
.B1(n_5400),
.B2(n_5409),
.C(n_5429),
.Y(n_5522)
);

AND2x2_ASAP7_75t_L g5523 ( 
.A(n_5416),
.B(n_5322),
.Y(n_5523)
);

INVx2_ASAP7_75t_L g5524 ( 
.A(n_5409),
.Y(n_5524)
);

INVx2_ASAP7_75t_L g5525 ( 
.A(n_5385),
.Y(n_5525)
);

AND2x4_ASAP7_75t_L g5526 ( 
.A(n_5463),
.B(n_5322),
.Y(n_5526)
);

AND2x4_ASAP7_75t_L g5527 ( 
.A(n_5463),
.B(n_5318),
.Y(n_5527)
);

INVx1_ASAP7_75t_L g5528 ( 
.A(n_5418),
.Y(n_5528)
);

INVx1_ASAP7_75t_L g5529 ( 
.A(n_5421),
.Y(n_5529)
);

NAND2x1p5_ASAP7_75t_SL g5530 ( 
.A(n_5419),
.B(n_5356),
.Y(n_5530)
);

BUFx2_ASAP7_75t_L g5531 ( 
.A(n_5465),
.Y(n_5531)
);

AND2x2_ASAP7_75t_L g5532 ( 
.A(n_5380),
.B(n_5290),
.Y(n_5532)
);

AND2x2_ASAP7_75t_L g5533 ( 
.A(n_5404),
.B(n_5316),
.Y(n_5533)
);

INVx1_ASAP7_75t_L g5534 ( 
.A(n_5372),
.Y(n_5534)
);

AND2x2_ASAP7_75t_L g5535 ( 
.A(n_5452),
.B(n_5316),
.Y(n_5535)
);

AND2x4_ASAP7_75t_L g5536 ( 
.A(n_5452),
.B(n_5323),
.Y(n_5536)
);

INVxp67_ASAP7_75t_SL g5537 ( 
.A(n_5400),
.Y(n_5537)
);

INVx1_ASAP7_75t_L g5538 ( 
.A(n_5429),
.Y(n_5538)
);

OR2x2_ASAP7_75t_L g5539 ( 
.A(n_5443),
.B(n_5240),
.Y(n_5539)
);

INVx1_ASAP7_75t_L g5540 ( 
.A(n_5432),
.Y(n_5540)
);

AND2x2_ASAP7_75t_L g5541 ( 
.A(n_5447),
.B(n_5327),
.Y(n_5541)
);

AOI211xp5_ASAP7_75t_SL g5542 ( 
.A1(n_5513),
.A2(n_5392),
.B(n_5412),
.C(n_5422),
.Y(n_5542)
);

OAI221xp5_ASAP7_75t_L g5543 ( 
.A1(n_5474),
.A2(n_5397),
.B1(n_5432),
.B2(n_5457),
.C(n_5453),
.Y(n_5543)
);

NAND2xp5_ASAP7_75t_L g5544 ( 
.A(n_5474),
.B(n_5466),
.Y(n_5544)
);

AOI221xp5_ASAP7_75t_L g5545 ( 
.A1(n_5508),
.A2(n_5466),
.B1(n_5457),
.B2(n_5453),
.C(n_5390),
.Y(n_5545)
);

OAI22xp5_ASAP7_75t_L g5546 ( 
.A1(n_5504),
.A2(n_5445),
.B1(n_5365),
.B2(n_5389),
.Y(n_5546)
);

INVx1_ASAP7_75t_L g5547 ( 
.A(n_5508),
.Y(n_5547)
);

OAI21xp5_ASAP7_75t_L g5548 ( 
.A1(n_5505),
.A2(n_5445),
.B(n_5458),
.Y(n_5548)
);

INVx1_ASAP7_75t_L g5549 ( 
.A(n_5528),
.Y(n_5549)
);

INVx2_ASAP7_75t_L g5550 ( 
.A(n_5501),
.Y(n_5550)
);

AND2x2_ASAP7_75t_L g5551 ( 
.A(n_5509),
.B(n_5369),
.Y(n_5551)
);

AOI33xp33_ASAP7_75t_L g5552 ( 
.A1(n_5502),
.A2(n_5365),
.A3(n_5439),
.B1(n_5389),
.B2(n_5390),
.B3(n_5370),
.Y(n_5552)
);

AND2x2_ASAP7_75t_L g5553 ( 
.A(n_5499),
.B(n_5369),
.Y(n_5553)
);

INVx1_ASAP7_75t_L g5554 ( 
.A(n_5470),
.Y(n_5554)
);

AND4x1_ASAP7_75t_L g5555 ( 
.A(n_5468),
.B(n_5420),
.C(n_5439),
.D(n_5337),
.Y(n_5555)
);

AOI211xp5_ASAP7_75t_L g5556 ( 
.A1(n_5522),
.A2(n_5430),
.B(n_5434),
.C(n_5369),
.Y(n_5556)
);

NAND4xp25_ASAP7_75t_L g5557 ( 
.A(n_5476),
.B(n_5430),
.C(n_5396),
.D(n_5465),
.Y(n_5557)
);

AND2x2_ASAP7_75t_L g5558 ( 
.A(n_5499),
.B(n_5366),
.Y(n_5558)
);

NAND4xp25_ASAP7_75t_SL g5559 ( 
.A(n_5476),
.B(n_5402),
.C(n_5406),
.D(n_5376),
.Y(n_5559)
);

HB1xp67_ASAP7_75t_L g5560 ( 
.A(n_5478),
.Y(n_5560)
);

INVx2_ASAP7_75t_L g5561 ( 
.A(n_5478),
.Y(n_5561)
);

HB1xp67_ASAP7_75t_L g5562 ( 
.A(n_5531),
.Y(n_5562)
);

A2O1A1Ixp33_ASAP7_75t_L g5563 ( 
.A1(n_5532),
.A2(n_5442),
.B(n_5444),
.C(n_5339),
.Y(n_5563)
);

INVx1_ASAP7_75t_L g5564 ( 
.A(n_5471),
.Y(n_5564)
);

INVx1_ASAP7_75t_L g5565 ( 
.A(n_5472),
.Y(n_5565)
);

NOR3xp33_ASAP7_75t_SL g5566 ( 
.A(n_5468),
.B(n_5223),
.C(n_5460),
.Y(n_5566)
);

INVx1_ASAP7_75t_L g5567 ( 
.A(n_5477),
.Y(n_5567)
);

BUFx2_ASAP7_75t_L g5568 ( 
.A(n_5480),
.Y(n_5568)
);

INVx1_ASAP7_75t_L g5569 ( 
.A(n_5481),
.Y(n_5569)
);

INVxp33_ASAP7_75t_L g5570 ( 
.A(n_5507),
.Y(n_5570)
);

CKINVDCx5p33_ASAP7_75t_R g5571 ( 
.A(n_5503),
.Y(n_5571)
);

NAND3xp33_ASAP7_75t_L g5572 ( 
.A(n_5469),
.B(n_5444),
.C(n_5442),
.Y(n_5572)
);

AOI22xp33_ASAP7_75t_L g5573 ( 
.A1(n_5488),
.A2(n_5435),
.B1(n_5441),
.B2(n_5382),
.Y(n_5573)
);

OAI21xp5_ASAP7_75t_SL g5574 ( 
.A1(n_5500),
.A2(n_5367),
.B(n_5428),
.Y(n_5574)
);

INVx1_ASAP7_75t_L g5575 ( 
.A(n_5496),
.Y(n_5575)
);

AOI22xp5_ASAP7_75t_L g5576 ( 
.A1(n_5532),
.A2(n_5435),
.B1(n_5441),
.B2(n_5451),
.Y(n_5576)
);

INVx2_ASAP7_75t_L g5577 ( 
.A(n_5503),
.Y(n_5577)
);

BUFx3_ASAP7_75t_L g5578 ( 
.A(n_5493),
.Y(n_5578)
);

NAND2xp33_ASAP7_75t_R g5579 ( 
.A(n_5536),
.B(n_5386),
.Y(n_5579)
);

NAND2xp5_ASAP7_75t_L g5580 ( 
.A(n_5469),
.B(n_5401),
.Y(n_5580)
);

AOI22xp5_ASAP7_75t_L g5581 ( 
.A1(n_5488),
.A2(n_5451),
.B1(n_5303),
.B2(n_5401),
.Y(n_5581)
);

NOR2xp33_ASAP7_75t_L g5582 ( 
.A(n_5507),
.B(n_5428),
.Y(n_5582)
);

AOI21xp5_ASAP7_75t_L g5583 ( 
.A1(n_5491),
.A2(n_5492),
.B(n_5485),
.Y(n_5583)
);

AOI22xp33_ASAP7_75t_L g5584 ( 
.A1(n_5491),
.A2(n_5357),
.B1(n_5382),
.B2(n_5425),
.Y(n_5584)
);

OAI31xp33_ASAP7_75t_L g5585 ( 
.A1(n_5492),
.A2(n_5358),
.A3(n_5399),
.B(n_5450),
.Y(n_5585)
);

AOI22xp33_ASAP7_75t_L g5586 ( 
.A1(n_5517),
.A2(n_5357),
.B1(n_5425),
.B2(n_5410),
.Y(n_5586)
);

OAI221xp5_ASAP7_75t_L g5587 ( 
.A1(n_5485),
.A2(n_5386),
.B1(n_5415),
.B2(n_5323),
.C(n_5449),
.Y(n_5587)
);

NAND2xp33_ASAP7_75t_SL g5588 ( 
.A(n_5500),
.B(n_5383),
.Y(n_5588)
);

INVx2_ASAP7_75t_L g5589 ( 
.A(n_5510),
.Y(n_5589)
);

INVx5_ASAP7_75t_L g5590 ( 
.A(n_5473),
.Y(n_5590)
);

AND2x2_ASAP7_75t_L g5591 ( 
.A(n_5558),
.B(n_5489),
.Y(n_5591)
);

INVx1_ASAP7_75t_L g5592 ( 
.A(n_5562),
.Y(n_5592)
);

NOR2xp67_ASAP7_75t_L g5593 ( 
.A(n_5574),
.B(n_5559),
.Y(n_5593)
);

AND2x2_ASAP7_75t_L g5594 ( 
.A(n_5553),
.B(n_5493),
.Y(n_5594)
);

NAND2xp5_ASAP7_75t_L g5595 ( 
.A(n_5552),
.B(n_5534),
.Y(n_5595)
);

OR2x2_ASAP7_75t_L g5596 ( 
.A(n_5544),
.B(n_5483),
.Y(n_5596)
);

INVx1_ASAP7_75t_L g5597 ( 
.A(n_5547),
.Y(n_5597)
);

INVx1_ASAP7_75t_L g5598 ( 
.A(n_5580),
.Y(n_5598)
);

INVx2_ASAP7_75t_L g5599 ( 
.A(n_5568),
.Y(n_5599)
);

AND2x2_ASAP7_75t_L g5600 ( 
.A(n_5551),
.B(n_5490),
.Y(n_5600)
);

INVx1_ASAP7_75t_L g5601 ( 
.A(n_5580),
.Y(n_5601)
);

OR2x2_ASAP7_75t_L g5602 ( 
.A(n_5544),
.B(n_5486),
.Y(n_5602)
);

INVx1_ASAP7_75t_L g5603 ( 
.A(n_5572),
.Y(n_5603)
);

OR2x2_ASAP7_75t_L g5604 ( 
.A(n_5550),
.B(n_5511),
.Y(n_5604)
);

INVx2_ASAP7_75t_SL g5605 ( 
.A(n_5590),
.Y(n_5605)
);

AND2x4_ASAP7_75t_SL g5606 ( 
.A(n_5560),
.B(n_5490),
.Y(n_5606)
);

INVx1_ASAP7_75t_L g5607 ( 
.A(n_5554),
.Y(n_5607)
);

NAND2xp5_ASAP7_75t_L g5608 ( 
.A(n_5546),
.B(n_5539),
.Y(n_5608)
);

AND2x2_ASAP7_75t_L g5609 ( 
.A(n_5578),
.B(n_5489),
.Y(n_5609)
);

AND2x4_ASAP7_75t_L g5610 ( 
.A(n_5589),
.B(n_5521),
.Y(n_5610)
);

OR2x2_ASAP7_75t_L g5611 ( 
.A(n_5546),
.B(n_5521),
.Y(n_5611)
);

AND2x2_ASAP7_75t_L g5612 ( 
.A(n_5566),
.B(n_5516),
.Y(n_5612)
);

NAND2xp5_ASAP7_75t_SL g5613 ( 
.A(n_5548),
.B(n_5473),
.Y(n_5613)
);

INVx2_ASAP7_75t_L g5614 ( 
.A(n_5576),
.Y(n_5614)
);

INVx1_ASAP7_75t_L g5615 ( 
.A(n_5564),
.Y(n_5615)
);

INVx1_ASAP7_75t_L g5616 ( 
.A(n_5565),
.Y(n_5616)
);

NAND2xp5_ASAP7_75t_SL g5617 ( 
.A(n_5548),
.B(n_5473),
.Y(n_5617)
);

NAND2xp5_ASAP7_75t_L g5618 ( 
.A(n_5542),
.B(n_5482),
.Y(n_5618)
);

INVx2_ASAP7_75t_L g5619 ( 
.A(n_5561),
.Y(n_5619)
);

INVx1_ASAP7_75t_L g5620 ( 
.A(n_5567),
.Y(n_5620)
);

NAND2x1p5_ASAP7_75t_L g5621 ( 
.A(n_5590),
.B(n_5473),
.Y(n_5621)
);

INVx1_ASAP7_75t_L g5622 ( 
.A(n_5569),
.Y(n_5622)
);

AND2x4_ASAP7_75t_L g5623 ( 
.A(n_5590),
.B(n_5523),
.Y(n_5623)
);

AND2x2_ASAP7_75t_L g5624 ( 
.A(n_5570),
.B(n_5512),
.Y(n_5624)
);

HB1xp67_ASAP7_75t_L g5625 ( 
.A(n_5577),
.Y(n_5625)
);

OR2x2_ASAP7_75t_L g5626 ( 
.A(n_5599),
.B(n_5557),
.Y(n_5626)
);

OR2x2_ASAP7_75t_L g5627 ( 
.A(n_5599),
.B(n_5549),
.Y(n_5627)
);

INVx1_ASAP7_75t_L g5628 ( 
.A(n_5625),
.Y(n_5628)
);

INVx2_ASAP7_75t_L g5629 ( 
.A(n_5591),
.Y(n_5629)
);

NAND2xp5_ASAP7_75t_L g5630 ( 
.A(n_5624),
.B(n_5542),
.Y(n_5630)
);

NAND2xp5_ASAP7_75t_L g5631 ( 
.A(n_5625),
.B(n_5563),
.Y(n_5631)
);

INVx2_ASAP7_75t_L g5632 ( 
.A(n_5591),
.Y(n_5632)
);

INVx1_ASAP7_75t_L g5633 ( 
.A(n_5592),
.Y(n_5633)
);

OR2x2_ASAP7_75t_L g5634 ( 
.A(n_5596),
.B(n_5602),
.Y(n_5634)
);

OR2x2_ASAP7_75t_L g5635 ( 
.A(n_5611),
.B(n_5588),
.Y(n_5635)
);

INVx1_ASAP7_75t_L g5636 ( 
.A(n_5604),
.Y(n_5636)
);

AND2x2_ASAP7_75t_L g5637 ( 
.A(n_5594),
.B(n_5533),
.Y(n_5637)
);

OR2x2_ASAP7_75t_L g5638 ( 
.A(n_5608),
.B(n_5520),
.Y(n_5638)
);

OR2x6_ASAP7_75t_L g5639 ( 
.A(n_5619),
.B(n_5583),
.Y(n_5639)
);

NAND2xp5_ASAP7_75t_L g5640 ( 
.A(n_5610),
.B(n_5571),
.Y(n_5640)
);

INVx1_ASAP7_75t_L g5641 ( 
.A(n_5619),
.Y(n_5641)
);

AOI21xp33_ASAP7_75t_SL g5642 ( 
.A1(n_5613),
.A2(n_5530),
.B(n_5579),
.Y(n_5642)
);

NAND2xp5_ASAP7_75t_L g5643 ( 
.A(n_5610),
.B(n_5609),
.Y(n_5643)
);

HB1xp67_ASAP7_75t_L g5644 ( 
.A(n_5610),
.Y(n_5644)
);

NAND2xp5_ASAP7_75t_L g5645 ( 
.A(n_5603),
.B(n_5537),
.Y(n_5645)
);

BUFx2_ASAP7_75t_L g5646 ( 
.A(n_5623),
.Y(n_5646)
);

AND2x2_ASAP7_75t_L g5647 ( 
.A(n_5600),
.B(n_5533),
.Y(n_5647)
);

INVx1_ASAP7_75t_L g5648 ( 
.A(n_5597),
.Y(n_5648)
);

NAND2xp5_ASAP7_75t_L g5649 ( 
.A(n_5606),
.B(n_5585),
.Y(n_5649)
);

INVx1_ASAP7_75t_SL g5650 ( 
.A(n_5635),
.Y(n_5650)
);

INVx2_ASAP7_75t_L g5651 ( 
.A(n_5639),
.Y(n_5651)
);

INVx2_ASAP7_75t_L g5652 ( 
.A(n_5639),
.Y(n_5652)
);

INVx2_ASAP7_75t_L g5653 ( 
.A(n_5639),
.Y(n_5653)
);

NOR2xp33_ASAP7_75t_L g5654 ( 
.A(n_5644),
.B(n_5606),
.Y(n_5654)
);

AND2x2_ASAP7_75t_L g5655 ( 
.A(n_5647),
.B(n_5535),
.Y(n_5655)
);

AND2x2_ASAP7_75t_L g5656 ( 
.A(n_5637),
.B(n_5535),
.Y(n_5656)
);

INVx1_ASAP7_75t_L g5657 ( 
.A(n_5629),
.Y(n_5657)
);

INVx4_ASAP7_75t_L g5658 ( 
.A(n_5646),
.Y(n_5658)
);

INVx2_ASAP7_75t_L g5659 ( 
.A(n_5632),
.Y(n_5659)
);

INVx1_ASAP7_75t_L g5660 ( 
.A(n_5636),
.Y(n_5660)
);

INVx1_ASAP7_75t_L g5661 ( 
.A(n_5628),
.Y(n_5661)
);

NAND2xp5_ASAP7_75t_L g5662 ( 
.A(n_5634),
.B(n_5623),
.Y(n_5662)
);

NAND2x1p5_ASAP7_75t_L g5663 ( 
.A(n_5641),
.B(n_5590),
.Y(n_5663)
);

INVx1_ASAP7_75t_L g5664 ( 
.A(n_5627),
.Y(n_5664)
);

INVx1_ASAP7_75t_L g5665 ( 
.A(n_5643),
.Y(n_5665)
);

INVx1_ASAP7_75t_L g5666 ( 
.A(n_5645),
.Y(n_5666)
);

AND2x2_ASAP7_75t_L g5667 ( 
.A(n_5640),
.B(n_5612),
.Y(n_5667)
);

INVx1_ASAP7_75t_SL g5668 ( 
.A(n_5631),
.Y(n_5668)
);

NOR2xp67_ASAP7_75t_L g5669 ( 
.A(n_5642),
.B(n_5582),
.Y(n_5669)
);

NOR2xp67_ASAP7_75t_L g5670 ( 
.A(n_5642),
.B(n_5623),
.Y(n_5670)
);

INVx2_ASAP7_75t_L g5671 ( 
.A(n_5638),
.Y(n_5671)
);

NOR2xp33_ASAP7_75t_SL g5672 ( 
.A(n_5626),
.B(n_5630),
.Y(n_5672)
);

NOR2xp33_ASAP7_75t_L g5673 ( 
.A(n_5649),
.B(n_5618),
.Y(n_5673)
);

AOI21xp5_ASAP7_75t_L g5674 ( 
.A1(n_5673),
.A2(n_5593),
.B(n_5613),
.Y(n_5674)
);

INVx2_ASAP7_75t_L g5675 ( 
.A(n_5658),
.Y(n_5675)
);

OAI22xp33_ASAP7_75t_SL g5676 ( 
.A1(n_5672),
.A2(n_5614),
.B1(n_5543),
.B2(n_5581),
.Y(n_5676)
);

NAND2xp5_ASAP7_75t_L g5677 ( 
.A(n_5658),
.B(n_5523),
.Y(n_5677)
);

INVxp67_ASAP7_75t_SL g5678 ( 
.A(n_5670),
.Y(n_5678)
);

AOI32xp33_ASAP7_75t_L g5679 ( 
.A1(n_5673),
.A2(n_5556),
.A3(n_5617),
.B1(n_5595),
.B2(n_5545),
.Y(n_5679)
);

OAI21xp5_ASAP7_75t_L g5680 ( 
.A1(n_5669),
.A2(n_5617),
.B(n_5654),
.Y(n_5680)
);

NAND2xp5_ASAP7_75t_L g5681 ( 
.A(n_5671),
.B(n_5648),
.Y(n_5681)
);

INVx2_ASAP7_75t_L g5682 ( 
.A(n_5655),
.Y(n_5682)
);

NAND2xp5_ASAP7_75t_L g5683 ( 
.A(n_5671),
.B(n_5607),
.Y(n_5683)
);

OAI21xp33_ASAP7_75t_SL g5684 ( 
.A1(n_5650),
.A2(n_5645),
.B(n_5605),
.Y(n_5684)
);

INVx2_ASAP7_75t_L g5685 ( 
.A(n_5656),
.Y(n_5685)
);

NAND2xp5_ASAP7_75t_L g5686 ( 
.A(n_5654),
.B(n_5615),
.Y(n_5686)
);

INVx1_ASAP7_75t_L g5687 ( 
.A(n_5659),
.Y(n_5687)
);

AOI22xp5_ASAP7_75t_L g5688 ( 
.A1(n_5668),
.A2(n_5614),
.B1(n_5573),
.B2(n_5494),
.Y(n_5688)
);

INVx1_ASAP7_75t_L g5689 ( 
.A(n_5659),
.Y(n_5689)
);

AOI22xp5_ASAP7_75t_L g5690 ( 
.A1(n_5651),
.A2(n_5494),
.B1(n_5515),
.B2(n_5587),
.Y(n_5690)
);

INVx1_ASAP7_75t_L g5691 ( 
.A(n_5677),
.Y(n_5691)
);

OR2x2_ASAP7_75t_L g5692 ( 
.A(n_5682),
.B(n_5664),
.Y(n_5692)
);

INVx1_ASAP7_75t_L g5693 ( 
.A(n_5685),
.Y(n_5693)
);

OR2x2_ASAP7_75t_L g5694 ( 
.A(n_5681),
.B(n_5662),
.Y(n_5694)
);

AND2x2_ASAP7_75t_L g5695 ( 
.A(n_5678),
.B(n_5667),
.Y(n_5695)
);

INVx1_ASAP7_75t_L g5696 ( 
.A(n_5687),
.Y(n_5696)
);

AND2x2_ASAP7_75t_L g5697 ( 
.A(n_5680),
.B(n_5665),
.Y(n_5697)
);

AND2x2_ASAP7_75t_L g5698 ( 
.A(n_5675),
.B(n_5657),
.Y(n_5698)
);

OR2x2_ASAP7_75t_L g5699 ( 
.A(n_5683),
.B(n_5660),
.Y(n_5699)
);

OAI31xp33_ASAP7_75t_SL g5700 ( 
.A1(n_5689),
.A2(n_5598),
.A3(n_5601),
.B(n_5666),
.Y(n_5700)
);

INVx1_ASAP7_75t_SL g5701 ( 
.A(n_5686),
.Y(n_5701)
);

NOR2xp33_ASAP7_75t_L g5702 ( 
.A(n_5684),
.B(n_5526),
.Y(n_5702)
);

INVx1_ASAP7_75t_L g5703 ( 
.A(n_5694),
.Y(n_5703)
);

INVx1_ASAP7_75t_L g5704 ( 
.A(n_5695),
.Y(n_5704)
);

INVx1_ASAP7_75t_L g5705 ( 
.A(n_5692),
.Y(n_5705)
);

INVx1_ASAP7_75t_L g5706 ( 
.A(n_5698),
.Y(n_5706)
);

AOI22xp5_ASAP7_75t_L g5707 ( 
.A1(n_5702),
.A2(n_5676),
.B1(n_5688),
.B2(n_5651),
.Y(n_5707)
);

INVx1_ASAP7_75t_L g5708 ( 
.A(n_5699),
.Y(n_5708)
);

NAND2xp5_ASAP7_75t_L g5709 ( 
.A(n_5701),
.B(n_5684),
.Y(n_5709)
);

NAND2x1_ASAP7_75t_L g5710 ( 
.A(n_5693),
.B(n_5605),
.Y(n_5710)
);

INVx1_ASAP7_75t_L g5711 ( 
.A(n_5697),
.Y(n_5711)
);

AND2x2_ASAP7_75t_L g5712 ( 
.A(n_5691),
.B(n_5674),
.Y(n_5712)
);

AOI322xp5_ASAP7_75t_L g5713 ( 
.A1(n_5696),
.A2(n_5652),
.A3(n_5653),
.B1(n_5690),
.B2(n_5515),
.C1(n_5584),
.C2(n_5586),
.Y(n_5713)
);

NAND2xp5_ASAP7_75t_SL g5714 ( 
.A(n_5700),
.B(n_5679),
.Y(n_5714)
);

NAND2xp5_ASAP7_75t_L g5715 ( 
.A(n_5691),
.B(n_5661),
.Y(n_5715)
);

NAND2xp5_ASAP7_75t_SL g5716 ( 
.A(n_5702),
.B(n_5506),
.Y(n_5716)
);

INVx1_ASAP7_75t_L g5717 ( 
.A(n_5712),
.Y(n_5717)
);

AND2x2_ASAP7_75t_SL g5718 ( 
.A(n_5709),
.B(n_5652),
.Y(n_5718)
);

O2A1O1Ixp33_ASAP7_75t_L g5719 ( 
.A1(n_5714),
.A2(n_5653),
.B(n_5663),
.C(n_5633),
.Y(n_5719)
);

A2O1A1Ixp33_ASAP7_75t_L g5720 ( 
.A1(n_5713),
.A2(n_5620),
.B(n_5622),
.C(n_5616),
.Y(n_5720)
);

NOR2xp33_ASAP7_75t_L g5721 ( 
.A(n_5703),
.B(n_5663),
.Y(n_5721)
);

NAND2xp5_ASAP7_75t_L g5722 ( 
.A(n_5705),
.B(n_5575),
.Y(n_5722)
);

AOI22x1_ASAP7_75t_L g5723 ( 
.A1(n_5704),
.A2(n_5621),
.B1(n_5506),
.B2(n_5467),
.Y(n_5723)
);

AND2x2_ASAP7_75t_L g5724 ( 
.A(n_5711),
.B(n_5467),
.Y(n_5724)
);

INVx1_ASAP7_75t_L g5725 ( 
.A(n_5706),
.Y(n_5725)
);

A2O1A1Ixp33_ASAP7_75t_L g5726 ( 
.A1(n_5707),
.A2(n_5524),
.B(n_5517),
.C(n_5525),
.Y(n_5726)
);

INVx1_ASAP7_75t_L g5727 ( 
.A(n_5708),
.Y(n_5727)
);

INVx1_ASAP7_75t_SL g5728 ( 
.A(n_5724),
.Y(n_5728)
);

AND2x2_ASAP7_75t_L g5729 ( 
.A(n_5717),
.B(n_5710),
.Y(n_5729)
);

INVx1_ASAP7_75t_L g5730 ( 
.A(n_5718),
.Y(n_5730)
);

INVx1_ASAP7_75t_L g5731 ( 
.A(n_5727),
.Y(n_5731)
);

AOI22xp33_ASAP7_75t_L g5732 ( 
.A1(n_5725),
.A2(n_5524),
.B1(n_5525),
.B2(n_5716),
.Y(n_5732)
);

INVx1_ASAP7_75t_L g5733 ( 
.A(n_5726),
.Y(n_5733)
);

NAND2xp5_ASAP7_75t_L g5734 ( 
.A(n_5721),
.B(n_5715),
.Y(n_5734)
);

AOI22xp33_ASAP7_75t_L g5735 ( 
.A1(n_5722),
.A2(n_5715),
.B1(n_5538),
.B2(n_5540),
.Y(n_5735)
);

INVx1_ASAP7_75t_L g5736 ( 
.A(n_5719),
.Y(n_5736)
);

OAI21xp33_ASAP7_75t_L g5737 ( 
.A1(n_5720),
.A2(n_5621),
.B(n_5506),
.Y(n_5737)
);

INVxp67_ASAP7_75t_SL g5738 ( 
.A(n_5723),
.Y(n_5738)
);

NAND2xp5_ASAP7_75t_L g5739 ( 
.A(n_5730),
.B(n_5555),
.Y(n_5739)
);

NAND2xp5_ASAP7_75t_L g5740 ( 
.A(n_5729),
.B(n_5541),
.Y(n_5740)
);

NOR2xp33_ASAP7_75t_L g5741 ( 
.A(n_5728),
.B(n_5479),
.Y(n_5741)
);

NOR3x1_ASAP7_75t_L g5742 ( 
.A(n_5738),
.B(n_5436),
.C(n_5484),
.Y(n_5742)
);

NOR4xp25_ASAP7_75t_L g5743 ( 
.A(n_5736),
.B(n_5449),
.C(n_5487),
.D(n_5497),
.Y(n_5743)
);

INVx1_ASAP7_75t_L g5744 ( 
.A(n_5734),
.Y(n_5744)
);

OAI21xp5_ASAP7_75t_L g5745 ( 
.A1(n_5731),
.A2(n_5495),
.B(n_5526),
.Y(n_5745)
);

INVxp67_ASAP7_75t_SL g5746 ( 
.A(n_5738),
.Y(n_5746)
);

NOR4xp25_ASAP7_75t_L g5747 ( 
.A(n_5733),
.B(n_5498),
.C(n_5518),
.D(n_5514),
.Y(n_5747)
);

NOR2x1_ASAP7_75t_L g5748 ( 
.A(n_5737),
.B(n_5536),
.Y(n_5748)
);

O2A1O1Ixp33_ASAP7_75t_L g5749 ( 
.A1(n_5732),
.A2(n_5536),
.B(n_5415),
.C(n_5526),
.Y(n_5749)
);

OAI21xp33_ASAP7_75t_L g5750 ( 
.A1(n_5735),
.A2(n_5415),
.B(n_5519),
.Y(n_5750)
);

NOR3xp33_ASAP7_75t_L g5751 ( 
.A(n_5730),
.B(n_5475),
.C(n_5527),
.Y(n_5751)
);

NOR3xp33_ASAP7_75t_L g5752 ( 
.A(n_5730),
.B(n_5527),
.C(n_5454),
.Y(n_5752)
);

OAI21xp33_ASAP7_75t_L g5753 ( 
.A1(n_5734),
.A2(n_5519),
.B(n_5431),
.Y(n_5753)
);

AOI21xp5_ASAP7_75t_L g5754 ( 
.A1(n_5734),
.A2(n_5527),
.B(n_5446),
.Y(n_5754)
);

NAND2xp5_ASAP7_75t_L g5755 ( 
.A(n_5730),
.B(n_5428),
.Y(n_5755)
);

AOI22xp5_ASAP7_75t_L g5756 ( 
.A1(n_5730),
.A2(n_5431),
.B1(n_5529),
.B2(n_5384),
.Y(n_5756)
);

HB1xp67_ASAP7_75t_L g5757 ( 
.A(n_5730),
.Y(n_5757)
);

NAND3xp33_ASAP7_75t_L g5758 ( 
.A(n_5730),
.B(n_5502),
.C(n_5431),
.Y(n_5758)
);

AOI211xp5_ASAP7_75t_L g5759 ( 
.A1(n_5746),
.A2(n_5395),
.B(n_5408),
.C(n_5437),
.Y(n_5759)
);

AOI221xp5_ASAP7_75t_L g5760 ( 
.A1(n_5757),
.A2(n_5530),
.B1(n_5459),
.B2(n_5456),
.C(n_5462),
.Y(n_5760)
);

AND2x4_ASAP7_75t_L g5761 ( 
.A(n_5745),
.B(n_5436),
.Y(n_5761)
);

NOR2x1_ASAP7_75t_L g5762 ( 
.A(n_5744),
.B(n_5461),
.Y(n_5762)
);

OR2x2_ASAP7_75t_L g5763 ( 
.A(n_5743),
.B(n_5755),
.Y(n_5763)
);

NOR3xp33_ASAP7_75t_L g5764 ( 
.A(n_5740),
.B(n_5427),
.C(n_5448),
.Y(n_5764)
);

NAND5xp2_ASAP7_75t_L g5765 ( 
.A(n_5751),
.B(n_5351),
.C(n_382),
.D(n_378),
.E(n_381),
.Y(n_5765)
);

NAND2xp5_ASAP7_75t_L g5766 ( 
.A(n_5754),
.B(n_5385),
.Y(n_5766)
);

AOI21xp33_ASAP7_75t_SL g5767 ( 
.A1(n_5739),
.A2(n_381),
.B(n_382),
.Y(n_5767)
);

NOR3xp33_ASAP7_75t_L g5768 ( 
.A(n_5741),
.B(n_5440),
.C(n_5410),
.Y(n_5768)
);

OAI21xp5_ASAP7_75t_L g5769 ( 
.A1(n_5758),
.A2(n_5748),
.B(n_5749),
.Y(n_5769)
);

NAND3xp33_ASAP7_75t_SL g5770 ( 
.A(n_5752),
.B(n_5440),
.C(n_383),
.Y(n_5770)
);

NAND3xp33_ASAP7_75t_L g5771 ( 
.A(n_5750),
.B(n_5747),
.C(n_5753),
.Y(n_5771)
);

INVx1_ASAP7_75t_L g5772 ( 
.A(n_5742),
.Y(n_5772)
);

INVx1_ASAP7_75t_L g5773 ( 
.A(n_5756),
.Y(n_5773)
);

AND2x2_ASAP7_75t_L g5774 ( 
.A(n_5745),
.B(n_383),
.Y(n_5774)
);

NOR2xp33_ASAP7_75t_L g5775 ( 
.A(n_5746),
.B(n_385),
.Y(n_5775)
);

NOR2xp33_ASAP7_75t_L g5776 ( 
.A(n_5746),
.B(n_386),
.Y(n_5776)
);

OAI21xp33_ASAP7_75t_L g5777 ( 
.A1(n_5753),
.A2(n_386),
.B(n_387),
.Y(n_5777)
);

NOR2x1_ASAP7_75t_L g5778 ( 
.A(n_5744),
.B(n_388),
.Y(n_5778)
);

INVxp67_ASAP7_75t_SL g5779 ( 
.A(n_5757),
.Y(n_5779)
);

NOR4xp25_ASAP7_75t_L g5780 ( 
.A(n_5746),
.B(n_390),
.C(n_388),
.D(n_389),
.Y(n_5780)
);

NAND2xp5_ASAP7_75t_L g5781 ( 
.A(n_5754),
.B(n_391),
.Y(n_5781)
);

NOR3x1_ASAP7_75t_SL g5782 ( 
.A(n_5757),
.B(n_391),
.C(n_392),
.Y(n_5782)
);

HB1xp67_ASAP7_75t_L g5783 ( 
.A(n_5748),
.Y(n_5783)
);

NAND4xp25_ASAP7_75t_SL g5784 ( 
.A(n_5771),
.B(n_5762),
.C(n_5781),
.D(n_5772),
.Y(n_5784)
);

OAI22xp5_ASAP7_75t_L g5785 ( 
.A1(n_5779),
.A2(n_395),
.B1(n_393),
.B2(n_394),
.Y(n_5785)
);

NOR4xp25_ASAP7_75t_L g5786 ( 
.A(n_5763),
.B(n_398),
.C(n_393),
.D(n_397),
.Y(n_5786)
);

NOR2x1p5_ASAP7_75t_L g5787 ( 
.A(n_5770),
.B(n_397),
.Y(n_5787)
);

NOR2xp33_ASAP7_75t_L g5788 ( 
.A(n_5783),
.B(n_398),
.Y(n_5788)
);

AOI22xp5_ASAP7_75t_L g5789 ( 
.A1(n_5766),
.A2(n_401),
.B1(n_399),
.B2(n_400),
.Y(n_5789)
);

NOR2x1_ASAP7_75t_L g5790 ( 
.A(n_5775),
.B(n_399),
.Y(n_5790)
);

AOI211xp5_ASAP7_75t_L g5791 ( 
.A1(n_5769),
.A2(n_403),
.B(n_400),
.C(n_402),
.Y(n_5791)
);

NOR3xp33_ASAP7_75t_L g5792 ( 
.A(n_5776),
.B(n_402),
.C(n_403),
.Y(n_5792)
);

INVx2_ASAP7_75t_L g5793 ( 
.A(n_5778),
.Y(n_5793)
);

NOR3x1_ASAP7_75t_L g5794 ( 
.A(n_5773),
.B(n_404),
.C(n_405),
.Y(n_5794)
);

INVx1_ASAP7_75t_L g5795 ( 
.A(n_5782),
.Y(n_5795)
);

NOR2x1_ASAP7_75t_L g5796 ( 
.A(n_5774),
.B(n_5765),
.Y(n_5796)
);

NAND2xp5_ASAP7_75t_L g5797 ( 
.A(n_5760),
.B(n_406),
.Y(n_5797)
);

INVx1_ASAP7_75t_L g5798 ( 
.A(n_5767),
.Y(n_5798)
);

OAI211xp5_ASAP7_75t_L g5799 ( 
.A1(n_5780),
.A2(n_408),
.B(n_406),
.C(n_407),
.Y(n_5799)
);

NAND3xp33_ASAP7_75t_L g5800 ( 
.A(n_5777),
.B(n_410),
.C(n_411),
.Y(n_5800)
);

OAI211xp5_ASAP7_75t_SL g5801 ( 
.A1(n_5768),
.A2(n_415),
.B(n_412),
.C(n_414),
.Y(n_5801)
);

A2O1A1Ixp33_ASAP7_75t_L g5802 ( 
.A1(n_5761),
.A2(n_417),
.B(n_415),
.C(n_416),
.Y(n_5802)
);

NOR2xp33_ASAP7_75t_L g5803 ( 
.A(n_5761),
.B(n_417),
.Y(n_5803)
);

NOR3xp33_ASAP7_75t_L g5804 ( 
.A(n_5759),
.B(n_418),
.C(n_419),
.Y(n_5804)
);

OAI211xp5_ASAP7_75t_L g5805 ( 
.A1(n_5764),
.A2(n_421),
.B(n_419),
.C(n_420),
.Y(n_5805)
);

NAND2xp5_ASAP7_75t_L g5806 ( 
.A(n_5779),
.B(n_423),
.Y(n_5806)
);

OAI21xp5_ASAP7_75t_L g5807 ( 
.A1(n_5779),
.A2(n_424),
.B(n_425),
.Y(n_5807)
);

OAI211xp5_ASAP7_75t_SL g5808 ( 
.A1(n_5772),
.A2(n_426),
.B(n_424),
.C(n_425),
.Y(n_5808)
);

NOR2xp33_ASAP7_75t_L g5809 ( 
.A(n_5779),
.B(n_426),
.Y(n_5809)
);

NOR4xp25_ASAP7_75t_L g5810 ( 
.A(n_5772),
.B(n_431),
.C(n_428),
.D(n_429),
.Y(n_5810)
);

AOI211xp5_ASAP7_75t_L g5811 ( 
.A1(n_5779),
.A2(n_433),
.B(n_429),
.C(n_432),
.Y(n_5811)
);

NAND3xp33_ASAP7_75t_SL g5812 ( 
.A(n_5763),
.B(n_434),
.C(n_437),
.Y(n_5812)
);

OAI211xp5_ASAP7_75t_L g5813 ( 
.A1(n_5810),
.A2(n_440),
.B(n_437),
.C(n_438),
.Y(n_5813)
);

NAND3xp33_ASAP7_75t_L g5814 ( 
.A(n_5795),
.B(n_5788),
.C(n_5793),
.Y(n_5814)
);

NOR3xp33_ASAP7_75t_L g5815 ( 
.A(n_5784),
.B(n_438),
.C(n_441),
.Y(n_5815)
);

AOI211xp5_ASAP7_75t_L g5816 ( 
.A1(n_5786),
.A2(n_443),
.B(n_441),
.C(n_442),
.Y(n_5816)
);

NOR3xp33_ASAP7_75t_L g5817 ( 
.A(n_5806),
.B(n_443),
.C(n_444),
.Y(n_5817)
);

NAND3xp33_ASAP7_75t_SL g5818 ( 
.A(n_5791),
.B(n_445),
.C(n_446),
.Y(n_5818)
);

AND2x2_ASAP7_75t_L g5819 ( 
.A(n_5796),
.B(n_447),
.Y(n_5819)
);

AOI22xp5_ASAP7_75t_L g5820 ( 
.A1(n_5803),
.A2(n_449),
.B1(n_447),
.B2(n_448),
.Y(n_5820)
);

NAND3x1_ASAP7_75t_L g5821 ( 
.A(n_5809),
.B(n_448),
.C(n_449),
.Y(n_5821)
);

NOR2xp33_ASAP7_75t_L g5822 ( 
.A(n_5799),
.B(n_450),
.Y(n_5822)
);

AOI311xp33_ASAP7_75t_L g5823 ( 
.A1(n_5804),
.A2(n_451),
.A3(n_452),
.B(n_453),
.C(n_454),
.Y(n_5823)
);

NAND4xp25_ASAP7_75t_L g5824 ( 
.A(n_5794),
.B(n_455),
.C(n_452),
.D(n_454),
.Y(n_5824)
);

OAI211xp5_ASAP7_75t_L g5825 ( 
.A1(n_5789),
.A2(n_457),
.B(n_455),
.C(n_456),
.Y(n_5825)
);

OAI221xp5_ASAP7_75t_L g5826 ( 
.A1(n_5802),
.A2(n_456),
.B1(n_457),
.B2(n_458),
.C(n_459),
.Y(n_5826)
);

NAND3xp33_ASAP7_75t_SL g5827 ( 
.A(n_5792),
.B(n_458),
.C(n_459),
.Y(n_5827)
);

NAND2xp5_ASAP7_75t_L g5828 ( 
.A(n_5790),
.B(n_460),
.Y(n_5828)
);

NAND4xp25_ASAP7_75t_L g5829 ( 
.A(n_5798),
.B(n_464),
.C(n_460),
.D(n_463),
.Y(n_5829)
);

OAI211xp5_ASAP7_75t_SL g5830 ( 
.A1(n_5797),
.A2(n_466),
.B(n_467),
.C(n_468),
.Y(n_5830)
);

NAND2xp5_ASAP7_75t_L g5831 ( 
.A(n_5787),
.B(n_467),
.Y(n_5831)
);

OA211x2_ASAP7_75t_L g5832 ( 
.A1(n_5807),
.A2(n_468),
.B(n_469),
.C(n_470),
.Y(n_5832)
);

NAND3xp33_ASAP7_75t_SL g5833 ( 
.A(n_5811),
.B(n_470),
.C(n_473),
.Y(n_5833)
);

AND4x2_ASAP7_75t_L g5834 ( 
.A(n_5812),
.B(n_473),
.C(n_474),
.D(n_475),
.Y(n_5834)
);

NOR2x1_ASAP7_75t_L g5835 ( 
.A(n_5785),
.B(n_475),
.Y(n_5835)
);

NOR3xp33_ASAP7_75t_L g5836 ( 
.A(n_5808),
.B(n_478),
.C(n_481),
.Y(n_5836)
);

NOR4xp25_ASAP7_75t_L g5837 ( 
.A(n_5805),
.B(n_478),
.C(n_481),
.D(n_482),
.Y(n_5837)
);

CKINVDCx5p33_ASAP7_75t_R g5838 ( 
.A(n_5819),
.Y(n_5838)
);

OR2x2_ASAP7_75t_L g5839 ( 
.A(n_5824),
.B(n_5800),
.Y(n_5839)
);

AOI22xp5_ASAP7_75t_L g5840 ( 
.A1(n_5814),
.A2(n_5801),
.B1(n_483),
.B2(n_484),
.Y(n_5840)
);

NAND2xp5_ASAP7_75t_L g5841 ( 
.A(n_5816),
.B(n_482),
.Y(n_5841)
);

INVx1_ASAP7_75t_L g5842 ( 
.A(n_5834),
.Y(n_5842)
);

NOR2x1_ASAP7_75t_L g5843 ( 
.A(n_5829),
.B(n_483),
.Y(n_5843)
);

NAND2xp5_ASAP7_75t_L g5844 ( 
.A(n_5821),
.B(n_484),
.Y(n_5844)
);

INVx1_ASAP7_75t_L g5845 ( 
.A(n_5828),
.Y(n_5845)
);

OAI21xp33_ASAP7_75t_L g5846 ( 
.A1(n_5822),
.A2(n_485),
.B(n_486),
.Y(n_5846)
);

AOI21xp33_ASAP7_75t_SL g5847 ( 
.A1(n_5815),
.A2(n_485),
.B(n_486),
.Y(n_5847)
);

AOI221xp5_ASAP7_75t_L g5848 ( 
.A1(n_5837),
.A2(n_487),
.B1(n_488),
.B2(n_489),
.C(n_491),
.Y(n_5848)
);

NOR2x1_ASAP7_75t_L g5849 ( 
.A(n_5831),
.B(n_487),
.Y(n_5849)
);

NOR2xp67_ASAP7_75t_L g5850 ( 
.A(n_5813),
.B(n_489),
.Y(n_5850)
);

INVx2_ASAP7_75t_SL g5851 ( 
.A(n_5835),
.Y(n_5851)
);

NAND2xp5_ASAP7_75t_L g5852 ( 
.A(n_5836),
.B(n_491),
.Y(n_5852)
);

OR2x2_ASAP7_75t_L g5853 ( 
.A(n_5827),
.B(n_492),
.Y(n_5853)
);

XOR2xp5_ASAP7_75t_L g5854 ( 
.A(n_5832),
.B(n_493),
.Y(n_5854)
);

NOR2x1p5_ASAP7_75t_L g5855 ( 
.A(n_5833),
.B(n_495),
.Y(n_5855)
);

HB1xp67_ASAP7_75t_L g5856 ( 
.A(n_5817),
.Y(n_5856)
);

INVx2_ASAP7_75t_L g5857 ( 
.A(n_5855),
.Y(n_5857)
);

NAND4xp75_ASAP7_75t_L g5858 ( 
.A(n_5849),
.B(n_5820),
.C(n_5823),
.D(n_5830),
.Y(n_5858)
);

NAND2x1p5_ASAP7_75t_L g5859 ( 
.A(n_5842),
.B(n_5818),
.Y(n_5859)
);

AND2x2_ASAP7_75t_L g5860 ( 
.A(n_5843),
.B(n_5825),
.Y(n_5860)
);

NOR3xp33_ASAP7_75t_L g5861 ( 
.A(n_5838),
.B(n_5826),
.C(n_495),
.Y(n_5861)
);

INVxp67_ASAP7_75t_SL g5862 ( 
.A(n_5844),
.Y(n_5862)
);

NAND2xp5_ASAP7_75t_L g5863 ( 
.A(n_5851),
.B(n_5850),
.Y(n_5863)
);

INVxp67_ASAP7_75t_L g5864 ( 
.A(n_5854),
.Y(n_5864)
);

NOR2xp67_ASAP7_75t_L g5865 ( 
.A(n_5847),
.B(n_497),
.Y(n_5865)
);

NOR2x1_ASAP7_75t_L g5866 ( 
.A(n_5853),
.B(n_497),
.Y(n_5866)
);

XNOR2xp5_ASAP7_75t_L g5867 ( 
.A(n_5856),
.B(n_498),
.Y(n_5867)
);

INVx1_ASAP7_75t_L g5868 ( 
.A(n_5841),
.Y(n_5868)
);

NOR4xp75_ASAP7_75t_L g5869 ( 
.A(n_5846),
.B(n_498),
.C(n_499),
.D(n_500),
.Y(n_5869)
);

NAND2xp5_ASAP7_75t_L g5870 ( 
.A(n_5845),
.B(n_500),
.Y(n_5870)
);

OR2x2_ASAP7_75t_L g5871 ( 
.A(n_5852),
.B(n_501),
.Y(n_5871)
);

AND3x4_ASAP7_75t_L g5872 ( 
.A(n_5848),
.B(n_501),
.C(n_502),
.Y(n_5872)
);

NAND3x1_ASAP7_75t_L g5873 ( 
.A(n_5866),
.B(n_5870),
.C(n_5863),
.Y(n_5873)
);

NAND5xp2_ASAP7_75t_L g5874 ( 
.A(n_5859),
.B(n_5840),
.C(n_5839),
.D(n_506),
.E(n_507),
.Y(n_5874)
);

NAND4xp75_ASAP7_75t_L g5875 ( 
.A(n_5865),
.B(n_504),
.C(n_505),
.D(n_507),
.Y(n_5875)
);

NOR4xp25_ASAP7_75t_L g5876 ( 
.A(n_5864),
.B(n_504),
.C(n_505),
.D(n_509),
.Y(n_5876)
);

NAND3xp33_ASAP7_75t_SL g5877 ( 
.A(n_5857),
.B(n_509),
.C(n_510),
.Y(n_5877)
);

INVx1_ASAP7_75t_L g5878 ( 
.A(n_5867),
.Y(n_5878)
);

NOR3xp33_ASAP7_75t_L g5879 ( 
.A(n_5862),
.B(n_510),
.C(n_511),
.Y(n_5879)
);

NAND3x1_ASAP7_75t_L g5880 ( 
.A(n_5869),
.B(n_511),
.C(n_512),
.Y(n_5880)
);

OA22x2_ASAP7_75t_L g5881 ( 
.A1(n_5872),
.A2(n_512),
.B1(n_513),
.B2(n_514),
.Y(n_5881)
);

NOR4xp25_ASAP7_75t_L g5882 ( 
.A(n_5868),
.B(n_513),
.C(n_514),
.D(n_515),
.Y(n_5882)
);

NOR3xp33_ASAP7_75t_L g5883 ( 
.A(n_5871),
.B(n_515),
.C(n_516),
.Y(n_5883)
);

NAND4xp25_ASAP7_75t_L g5884 ( 
.A(n_5860),
.B(n_5861),
.C(n_5858),
.D(n_520),
.Y(n_5884)
);

OR5x1_ASAP7_75t_L g5885 ( 
.A(n_5872),
.B(n_517),
.C(n_518),
.D(n_520),
.E(n_521),
.Y(n_5885)
);

NAND2xp5_ASAP7_75t_L g5886 ( 
.A(n_5862),
.B(n_517),
.Y(n_5886)
);

NOR2x2_ASAP7_75t_L g5887 ( 
.A(n_5858),
.B(n_521),
.Y(n_5887)
);

NOR4xp25_ASAP7_75t_L g5888 ( 
.A(n_5863),
.B(n_522),
.C(n_523),
.D(n_524),
.Y(n_5888)
);

AOI211xp5_ASAP7_75t_SL g5889 ( 
.A1(n_5864),
.A2(n_523),
.B(n_524),
.C(n_526),
.Y(n_5889)
);

NOR2xp67_ASAP7_75t_L g5890 ( 
.A(n_5867),
.B(n_529),
.Y(n_5890)
);

CKINVDCx5p33_ASAP7_75t_R g5891 ( 
.A(n_5878),
.Y(n_5891)
);

INVx1_ASAP7_75t_L g5892 ( 
.A(n_5890),
.Y(n_5892)
);

INVx1_ASAP7_75t_L g5893 ( 
.A(n_5881),
.Y(n_5893)
);

A2O1A1Ixp33_ASAP7_75t_L g5894 ( 
.A1(n_5889),
.A2(n_529),
.B(n_530),
.C(n_531),
.Y(n_5894)
);

OAI322xp33_ASAP7_75t_L g5895 ( 
.A1(n_5886),
.A2(n_532),
.A3(n_533),
.B1(n_534),
.B2(n_536),
.C1(n_537),
.C2(n_538),
.Y(n_5895)
);

CKINVDCx5p33_ASAP7_75t_R g5896 ( 
.A(n_5873),
.Y(n_5896)
);

CKINVDCx5p33_ASAP7_75t_R g5897 ( 
.A(n_5887),
.Y(n_5897)
);

CKINVDCx5p33_ASAP7_75t_R g5898 ( 
.A(n_5877),
.Y(n_5898)
);

AOI22xp33_ASAP7_75t_SL g5899 ( 
.A1(n_5885),
.A2(n_538),
.B1(n_539),
.B2(n_540),
.Y(n_5899)
);

INVx1_ASAP7_75t_L g5900 ( 
.A(n_5880),
.Y(n_5900)
);

INVx1_ASAP7_75t_L g5901 ( 
.A(n_5875),
.Y(n_5901)
);

INVx1_ASAP7_75t_L g5902 ( 
.A(n_5874),
.Y(n_5902)
);

CKINVDCx20_ASAP7_75t_R g5903 ( 
.A(n_5884),
.Y(n_5903)
);

INVx1_ASAP7_75t_L g5904 ( 
.A(n_5883),
.Y(n_5904)
);

NOR2x1p5_ASAP7_75t_L g5905 ( 
.A(n_5896),
.B(n_5876),
.Y(n_5905)
);

CKINVDCx20_ASAP7_75t_R g5906 ( 
.A(n_5891),
.Y(n_5906)
);

NAND3xp33_ASAP7_75t_SL g5907 ( 
.A(n_5897),
.B(n_5879),
.C(n_5888),
.Y(n_5907)
);

AOI22xp5_ASAP7_75t_L g5908 ( 
.A1(n_5903),
.A2(n_5882),
.B1(n_541),
.B2(n_542),
.Y(n_5908)
);

OAI22xp5_ASAP7_75t_L g5909 ( 
.A1(n_5902),
.A2(n_539),
.B1(n_542),
.B2(n_543),
.Y(n_5909)
);

OAI221xp5_ASAP7_75t_L g5910 ( 
.A1(n_5899),
.A2(n_544),
.B1(n_545),
.B2(n_546),
.C(n_548),
.Y(n_5910)
);

AND2x4_ASAP7_75t_L g5911 ( 
.A(n_5892),
.B(n_544),
.Y(n_5911)
);

AOI322xp5_ASAP7_75t_L g5912 ( 
.A1(n_5900),
.A2(n_549),
.A3(n_550),
.B1(n_551),
.B2(n_552),
.C1(n_553),
.C2(n_555),
.Y(n_5912)
);

INVx2_ASAP7_75t_L g5913 ( 
.A(n_5906),
.Y(n_5913)
);

INVx1_ASAP7_75t_L g5914 ( 
.A(n_5905),
.Y(n_5914)
);

INVx2_ASAP7_75t_L g5915 ( 
.A(n_5911),
.Y(n_5915)
);

INVx1_ASAP7_75t_L g5916 ( 
.A(n_5907),
.Y(n_5916)
);

OAI22xp5_ASAP7_75t_L g5917 ( 
.A1(n_5910),
.A2(n_5893),
.B1(n_5894),
.B2(n_5898),
.Y(n_5917)
);

AOI22xp5_ASAP7_75t_L g5918 ( 
.A1(n_5908),
.A2(n_5901),
.B1(n_5904),
.B2(n_5895),
.Y(n_5918)
);

AOI22xp33_ASAP7_75t_SL g5919 ( 
.A1(n_5909),
.A2(n_549),
.B1(n_550),
.B2(n_553),
.Y(n_5919)
);

CKINVDCx20_ASAP7_75t_R g5920 ( 
.A(n_5912),
.Y(n_5920)
);

OAI22xp5_ASAP7_75t_L g5921 ( 
.A1(n_5913),
.A2(n_555),
.B1(n_556),
.B2(n_558),
.Y(n_5921)
);

AOI221xp5_ASAP7_75t_L g5922 ( 
.A1(n_5916),
.A2(n_5914),
.B1(n_5917),
.B2(n_5915),
.C(n_5920),
.Y(n_5922)
);

AOI22xp33_ASAP7_75t_L g5923 ( 
.A1(n_5919),
.A2(n_559),
.B1(n_560),
.B2(n_563),
.Y(n_5923)
);

XNOR2x1_ASAP7_75t_L g5924 ( 
.A(n_5918),
.B(n_560),
.Y(n_5924)
);

NAND3xp33_ASAP7_75t_L g5925 ( 
.A(n_5913),
.B(n_563),
.C(n_564),
.Y(n_5925)
);

AND4x1_ASAP7_75t_L g5926 ( 
.A(n_5914),
.B(n_564),
.C(n_565),
.D(n_566),
.Y(n_5926)
);

XNOR2xp5_ASAP7_75t_L g5927 ( 
.A(n_5922),
.B(n_565),
.Y(n_5927)
);

AOI22x1_ASAP7_75t_L g5928 ( 
.A1(n_5924),
.A2(n_567),
.B1(n_568),
.B2(n_569),
.Y(n_5928)
);

OAI22xp33_ASAP7_75t_L g5929 ( 
.A1(n_5925),
.A2(n_568),
.B1(n_569),
.B2(n_571),
.Y(n_5929)
);

OAI22xp5_ASAP7_75t_L g5930 ( 
.A1(n_5923),
.A2(n_571),
.B1(n_572),
.B2(n_573),
.Y(n_5930)
);

AOI22xp33_ASAP7_75t_L g5931 ( 
.A1(n_5921),
.A2(n_574),
.B1(n_575),
.B2(n_576),
.Y(n_5931)
);

INVxp67_ASAP7_75t_SL g5932 ( 
.A(n_5927),
.Y(n_5932)
);

AOI22xp33_ASAP7_75t_L g5933 ( 
.A1(n_5928),
.A2(n_5926),
.B1(n_577),
.B2(n_578),
.Y(n_5933)
);

OAI22xp5_ASAP7_75t_SL g5934 ( 
.A1(n_5931),
.A2(n_574),
.B1(n_577),
.B2(n_578),
.Y(n_5934)
);

HB1xp67_ASAP7_75t_L g5935 ( 
.A(n_5930),
.Y(n_5935)
);

OAI22xp33_ASAP7_75t_L g5936 ( 
.A1(n_5932),
.A2(n_5929),
.B1(n_580),
.B2(n_581),
.Y(n_5936)
);

AOI21xp5_ASAP7_75t_L g5937 ( 
.A1(n_5935),
.A2(n_579),
.B(n_580),
.Y(n_5937)
);

OAI21x1_ASAP7_75t_SL g5938 ( 
.A1(n_5933),
.A2(n_5934),
.B(n_582),
.Y(n_5938)
);

INVx1_ASAP7_75t_L g5939 ( 
.A(n_5932),
.Y(n_5939)
);

OAI22xp5_ASAP7_75t_L g5940 ( 
.A1(n_5933),
.A2(n_579),
.B1(n_583),
.B2(n_584),
.Y(n_5940)
);

OAI21xp5_ASAP7_75t_L g5941 ( 
.A1(n_5939),
.A2(n_583),
.B(n_585),
.Y(n_5941)
);

AOI21xp5_ASAP7_75t_L g5942 ( 
.A1(n_5938),
.A2(n_5940),
.B(n_5936),
.Y(n_5942)
);

OAI21xp33_ASAP7_75t_SL g5943 ( 
.A1(n_5937),
.A2(n_587),
.B(n_588),
.Y(n_5943)
);

AOI21xp5_ASAP7_75t_L g5944 ( 
.A1(n_5939),
.A2(n_588),
.B(n_589),
.Y(n_5944)
);

AOI221xp5_ASAP7_75t_L g5945 ( 
.A1(n_5939),
.A2(n_590),
.B1(n_591),
.B2(n_592),
.C(n_593),
.Y(n_5945)
);

AOI21xp5_ASAP7_75t_L g5946 ( 
.A1(n_5939),
.A2(n_590),
.B(n_591),
.Y(n_5946)
);

NOR2x1_ASAP7_75t_L g5947 ( 
.A(n_5939),
.B(n_595),
.Y(n_5947)
);

INVx1_ASAP7_75t_L g5948 ( 
.A(n_5939),
.Y(n_5948)
);

XNOR2xp5_ASAP7_75t_L g5949 ( 
.A(n_5939),
.B(n_595),
.Y(n_5949)
);

INVx1_ASAP7_75t_L g5950 ( 
.A(n_5939),
.Y(n_5950)
);

AOI22xp5_ASAP7_75t_L g5951 ( 
.A1(n_5948),
.A2(n_596),
.B1(n_598),
.B2(n_599),
.Y(n_5951)
);

AO22x1_ASAP7_75t_L g5952 ( 
.A1(n_5950),
.A2(n_598),
.B1(n_599),
.B2(n_600),
.Y(n_5952)
);

AOI22xp5_ASAP7_75t_L g5953 ( 
.A1(n_5947),
.A2(n_600),
.B1(n_602),
.B2(n_603),
.Y(n_5953)
);

OAI22xp5_ASAP7_75t_L g5954 ( 
.A1(n_5949),
.A2(n_5946),
.B1(n_5944),
.B2(n_5942),
.Y(n_5954)
);

AO22x2_ASAP7_75t_L g5955 ( 
.A1(n_5941),
.A2(n_602),
.B1(n_603),
.B2(n_604),
.Y(n_5955)
);

AOI22xp5_ASAP7_75t_L g5956 ( 
.A1(n_5943),
.A2(n_604),
.B1(n_605),
.B2(n_606),
.Y(n_5956)
);

AOI22xp5_ASAP7_75t_L g5957 ( 
.A1(n_5945),
.A2(n_606),
.B1(n_607),
.B2(n_608),
.Y(n_5957)
);

AOI22xp5_ASAP7_75t_L g5958 ( 
.A1(n_5948),
.A2(n_607),
.B1(n_609),
.B2(n_611),
.Y(n_5958)
);

OAI22xp5_ASAP7_75t_L g5959 ( 
.A1(n_5948),
.A2(n_609),
.B1(n_612),
.B2(n_613),
.Y(n_5959)
);

OAI22xp33_ASAP7_75t_L g5960 ( 
.A1(n_5948),
.A2(n_612),
.B1(n_614),
.B2(n_615),
.Y(n_5960)
);

AOI21xp5_ASAP7_75t_L g5961 ( 
.A1(n_5954),
.A2(n_614),
.B(n_616),
.Y(n_5961)
);

OAI21xp5_ASAP7_75t_L g5962 ( 
.A1(n_5956),
.A2(n_616),
.B(n_617),
.Y(n_5962)
);

NAND2xp5_ASAP7_75t_L g5963 ( 
.A(n_5955),
.B(n_617),
.Y(n_5963)
);

AOI21xp5_ASAP7_75t_L g5964 ( 
.A1(n_5952),
.A2(n_5960),
.B(n_5953),
.Y(n_5964)
);

AND2x2_ASAP7_75t_L g5965 ( 
.A(n_5957),
.B(n_5951),
.Y(n_5965)
);

XNOR2xp5_ASAP7_75t_L g5966 ( 
.A(n_5958),
.B(n_618),
.Y(n_5966)
);

OAI21xp5_ASAP7_75t_SL g5967 ( 
.A1(n_5959),
.A2(n_618),
.B(n_620),
.Y(n_5967)
);

OR2x2_ASAP7_75t_L g5968 ( 
.A(n_5956),
.B(n_620),
.Y(n_5968)
);

OAI22xp33_ASAP7_75t_L g5969 ( 
.A1(n_5963),
.A2(n_622),
.B1(n_623),
.B2(n_624),
.Y(n_5969)
);

OAI22xp5_ASAP7_75t_SL g5970 ( 
.A1(n_5966),
.A2(n_622),
.B1(n_626),
.B2(n_627),
.Y(n_5970)
);

HB1xp67_ASAP7_75t_L g5971 ( 
.A(n_5968),
.Y(n_5971)
);

INVx1_ASAP7_75t_L g5972 ( 
.A(n_5965),
.Y(n_5972)
);

OAI22xp33_ASAP7_75t_L g5973 ( 
.A1(n_5967),
.A2(n_626),
.B1(n_627),
.B2(n_633),
.Y(n_5973)
);

AOI221xp5_ASAP7_75t_L g5974 ( 
.A1(n_5972),
.A2(n_5964),
.B1(n_5961),
.B2(n_5962),
.C(n_636),
.Y(n_5974)
);

AOI221xp5_ASAP7_75t_L g5975 ( 
.A1(n_5974),
.A2(n_5971),
.B1(n_5969),
.B2(n_5973),
.C(n_5970),
.Y(n_5975)
);

AOI211xp5_ASAP7_75t_L g5976 ( 
.A1(n_5975),
.A2(n_633),
.B(n_634),
.C(n_635),
.Y(n_5976)
);


endmodule