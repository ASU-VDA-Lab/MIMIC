module fake_jpeg_25326_n_307 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_307);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_307;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_44),
.Y(n_62)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_24),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_45),
.B(n_47),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_24),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_22),
.B1(n_18),
.B2(n_17),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_51),
.A2(n_52),
.B1(n_57),
.B2(n_61),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_26),
.B1(n_17),
.B2(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_53),
.B(n_55),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_33),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_34),
.B1(n_24),
.B2(n_16),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_59),
.B1(n_60),
.B2(n_41),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_18),
.B1(n_30),
.B2(n_26),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_58),
.B(n_66),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_34),
.B1(n_16),
.B2(n_28),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_38),
.A2(n_34),
.B1(n_16),
.B2(n_28),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_30),
.B1(n_26),
.B2(n_17),
.Y(n_61)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_39),
.B(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_20),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_67),
.B(n_35),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_20),
.B(n_19),
.C(n_28),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_68),
.B(n_85),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_71),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_72),
.B(n_75),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_73),
.A2(n_82),
.B1(n_27),
.B2(n_63),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_20),
.B1(n_19),
.B2(n_31),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_74),
.A2(n_83),
.B1(n_92),
.B2(n_97),
.Y(n_115)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

AO22x1_ASAP7_75t_SL g76 ( 
.A1(n_55),
.A2(n_37),
.B1(n_39),
.B2(n_41),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_76),
.A2(n_90),
.B1(n_21),
.B2(n_33),
.Y(n_134)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_77),
.B(n_80),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_78),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_41),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_81),
.A2(n_99),
.B1(n_32),
.B2(n_25),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_57),
.A2(n_37),
.B1(n_27),
.B2(n_23),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_84),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_29),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_62),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_91),
.Y(n_129)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

AO22x1_ASAP7_75t_SL g90 ( 
.A1(n_55),
.A2(n_37),
.B1(n_39),
.B2(n_21),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_67),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_50),
.A2(n_35),
.B1(n_31),
.B2(n_30),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_93),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_58),
.B(n_29),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_102),
.Y(n_109)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_56),
.Y(n_99)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_101),
.A2(n_105),
.B1(n_64),
.B2(n_54),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_53),
.B(n_29),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_15),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_59),
.B(n_31),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_27),
.Y(n_118)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_100),
.B(n_55),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_107),
.A2(n_90),
.B(n_93),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_94),
.B(n_55),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_108),
.B(n_112),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_110),
.B(n_12),
.Y(n_158)
);

NAND2x1_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_51),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_106),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_116),
.A2(n_118),
.B(n_21),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_117),
.Y(n_145)
);

FAx1_ASAP7_75t_SL g121 ( 
.A(n_106),
.B(n_63),
.CI(n_49),
.CON(n_121),
.SN(n_121)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_76),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_75),
.A2(n_63),
.B1(n_64),
.B2(n_32),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_122),
.A2(n_134),
.B1(n_81),
.B2(n_80),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_126),
.A2(n_101),
.B1(n_105),
.B2(n_86),
.Y(n_152)
);

OAI22x1_ASAP7_75t_L g130 ( 
.A1(n_76),
.A2(n_29),
.B1(n_25),
.B2(n_32),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_130),
.A2(n_124),
.B1(n_123),
.B2(n_115),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_94),
.B(n_32),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_90),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_136),
.A2(n_163),
.B1(n_165),
.B2(n_166),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_137),
.A2(n_130),
.B(n_121),
.C(n_107),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_112),
.A2(n_68),
.B(n_98),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_138),
.A2(n_153),
.B(n_167),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_129),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_139),
.B(n_158),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_98),
.B1(n_81),
.B2(n_71),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_140),
.A2(n_142),
.B1(n_155),
.B2(n_124),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_88),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_143),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_134),
.A2(n_107),
.B1(n_125),
.B2(n_116),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_135),
.B(n_131),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_146),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_111),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_89),
.Y(n_147)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_150),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_131),
.B(n_116),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_151),
.B(n_164),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_152),
.A2(n_154),
.B1(n_156),
.B2(n_153),
.Y(n_168)
);

NOR2x1_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_77),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_126),
.A2(n_72),
.B1(n_69),
.B2(n_83),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_107),
.A2(n_69),
.B1(n_32),
.B2(n_23),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_109),
.B(n_84),
.Y(n_159)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_109),
.B(n_78),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_160),
.Y(n_195)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

INVx5_ASAP7_75t_SL g179 ( 
.A(n_162),
.Y(n_179)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_118),
.B(n_21),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_168),
.A2(n_190),
.B(n_149),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_169),
.B(n_155),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_108),
.C(n_133),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_170),
.B(n_176),
.C(n_182),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_188),
.Y(n_206)
);

INVxp33_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_174),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_132),
.C(n_127),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_178),
.A2(n_181),
.B1(n_186),
.B2(n_194),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_163),
.A2(n_120),
.B1(n_132),
.B2(n_114),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_127),
.C(n_114),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_147),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_184),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_165),
.A2(n_120),
.B1(n_113),
.B2(n_123),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_159),
.Y(n_188)
);

AOI322xp5_ASAP7_75t_L g189 ( 
.A1(n_150),
.A2(n_110),
.A3(n_25),
.B1(n_23),
.B2(n_113),
.C1(n_119),
.C2(n_123),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_189),
.B(n_192),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_139),
.B(n_119),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_146),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_110),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_196),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_136),
.A2(n_119),
.B1(n_23),
.B2(n_25),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_142),
.B(n_15),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_200),
.A2(n_202),
.B(n_207),
.Y(n_239)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_201),
.B(n_204),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_137),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_143),
.Y(n_203)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_179),
.A2(n_145),
.B1(n_197),
.B2(n_183),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_205),
.A2(n_217),
.B1(n_220),
.B2(n_183),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_140),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_178),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_211),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_180),
.A2(n_166),
.B1(n_153),
.B2(n_152),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_210),
.A2(n_222),
.B1(n_185),
.B2(n_195),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_172),
.B(n_158),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_168),
.A2(n_138),
.B1(n_148),
.B2(n_151),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_213),
.A2(n_185),
.B1(n_169),
.B2(n_190),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_190),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_174),
.Y(n_233)
);

XNOR2x1_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_138),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_219),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_179),
.A2(n_144),
.B1(n_162),
.B2(n_157),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_187),
.A2(n_154),
.B1(n_167),
.B2(n_15),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_170),
.B(n_182),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_171),
.C(n_193),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_173),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_206),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_226),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_229),
.Y(n_246)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_228),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_208),
.A2(n_213),
.B1(n_216),
.B2(n_198),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_230),
.A2(n_232),
.B1(n_237),
.B2(n_241),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_202),
.A2(n_187),
.B1(n_177),
.B2(n_196),
.Y(n_232)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_199),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_191),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_235),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_221),
.C(n_171),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_238),
.C(n_215),
.Y(n_245)
);

OAI22x1_ASAP7_75t_L g237 ( 
.A1(n_200),
.A2(n_187),
.B1(n_191),
.B2(n_2),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_14),
.C(n_13),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_202),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_222),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_242),
.B(n_220),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_235),
.C(n_228),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_240),
.Y(n_247)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_247),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_231),
.Y(n_248)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_248),
.Y(n_262)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_238),
.B(n_212),
.Y(n_250)
);

OAI322xp33_ASAP7_75t_L g263 ( 
.A1(n_250),
.A2(n_251),
.A3(n_237),
.B1(n_252),
.B2(n_223),
.C1(n_232),
.C2(n_246),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_223),
.B(n_207),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_215),
.C(n_219),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_256),
.C(n_258),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_226),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_243),
.C(n_230),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_218),
.C(n_199),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_214),
.C(n_13),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_225),
.C(n_239),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_263),
.A2(n_244),
.B1(n_259),
.B2(n_257),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_268),
.C(n_269),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_239),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_267),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_12),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_9),
.C(n_1),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_273),
.C(n_260),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_258),
.B(n_9),
.Y(n_271)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_271),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_9),
.C(n_1),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_267),
.A2(n_255),
.B1(n_246),
.B2(n_259),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_274),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_289)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_277),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_278),
.A2(n_280),
.B(n_284),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_265),
.A2(n_257),
.B1(n_1),
.B2(n_2),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_279),
.A2(n_282),
.B1(n_0),
.B2(n_5),
.Y(n_292)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_271),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_7),
.C(n_1),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_269),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_272),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_282)
);

AO21x1_ASAP7_75t_L g284 ( 
.A1(n_261),
.A2(n_0),
.B(n_3),
.Y(n_284)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_286),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_264),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_287),
.B(n_289),
.Y(n_295)
);

OA21x2_ASAP7_75t_L g288 ( 
.A1(n_274),
.A2(n_262),
.B(n_4),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_290),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_280),
.A2(n_275),
.B(n_283),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_279),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_296),
.B(n_297),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_285),
.B(n_286),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_295),
.A2(n_291),
.B(n_287),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_298),
.B(n_299),
.Y(n_301)
);

AOI21xp33_ASAP7_75t_L g300 ( 
.A1(n_293),
.A2(n_290),
.B(n_288),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_288),
.C(n_294),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_301),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_303),
.A2(n_302),
.B1(n_282),
.B2(n_281),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_304),
.A2(n_284),
.B(n_276),
.Y(n_305)
);

AOI221xp5_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_277),
.B1(n_6),
.B2(n_7),
.C(n_5),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_7),
.Y(n_307)
);


endmodule