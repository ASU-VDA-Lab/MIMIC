module fake_jpeg_23793_n_178 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_178);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_31),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_18),
.A2(n_0),
.B(n_1),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_18),
.B1(n_22),
.B2(n_13),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_13),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_33),
.B(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_47),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_48),
.B1(n_17),
.B2(n_28),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_30),
.B(n_14),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_22),
.C(n_13),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_16),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_22),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_28),
.A2(n_17),
.B1(n_16),
.B2(n_24),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_26),
.Y(n_50)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_53),
.B(n_67),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_55),
.B(n_58),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_56),
.A2(n_57),
.B1(n_52),
.B2(n_44),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_29),
.B1(n_17),
.B2(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_21),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_45),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_59),
.B(n_61),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_1),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_49),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_64),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_49),
.B(n_24),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_23),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_19),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_69),
.B(n_71),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_52),
.B1(n_51),
.B2(n_39),
.Y(n_74)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_41),
.Y(n_75)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_58),
.A2(n_39),
.B1(n_44),
.B2(n_43),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_79),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_59),
.A2(n_19),
.B1(n_26),
.B2(n_23),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_80),
.A2(n_83),
.B(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_41),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_81),
.B(n_54),
.Y(n_86)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

OAI32xp33_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_36),
.A3(n_34),
.B1(n_27),
.B2(n_21),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_86),
.B(n_88),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_72),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_87),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_73),
.Y(n_88)
);

CKINVDCx10_ASAP7_75t_R g89 ( 
.A(n_82),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_89),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_60),
.B(n_66),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_69),
.B(n_25),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_83),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_97),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_65),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_101),
.C(n_84),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_14),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_98),
.B(n_84),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_63),
.C(n_68),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_112),
.C(n_115),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_105),
.Y(n_127)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_99),
.A2(n_71),
.B1(n_74),
.B2(n_78),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_111),
.B1(n_116),
.B2(n_94),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_89),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_108),
.A2(n_110),
.B(n_114),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_115),
.B1(n_94),
.B2(n_25),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_99),
.A2(n_54),
.B(n_68),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_97),
.A2(n_63),
.B1(n_40),
.B2(n_36),
.Y(n_111)
);

XOR2x2_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_69),
.Y(n_112)
);

OA21x2_ASAP7_75t_SL g130 ( 
.A1(n_112),
.A2(n_92),
.B(n_25),
.Y(n_130)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_95),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_90),
.A2(n_36),
.B(n_34),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_119),
.C(n_123),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_91),
.C(n_96),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_120),
.Y(n_138)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_125),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_104),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_129),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_114),
.Y(n_142)
);

NAND3xp33_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_92),
.C(n_7),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_102),
.C(n_110),
.Y(n_140)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_127),
.B(n_117),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_134),
.B(n_121),
.Y(n_148)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_137),
.A2(n_142),
.B(n_143),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_119),
.C(n_123),
.Y(n_146)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_141),
.B(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_152),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_118),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_146),
.C(n_147),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_124),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_153),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_107),
.C(n_15),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_151),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_15),
.C(n_21),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_15),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_15),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_150),
.A2(n_138),
.B1(n_143),
.B2(n_136),
.Y(n_154)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_154),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_133),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_160),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_136),
.B1(n_135),
.B2(n_142),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_147),
.B(n_132),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_2),
.Y(n_167)
);

AOI21xp33_ASAP7_75t_L g163 ( 
.A1(n_159),
.A2(n_135),
.B(n_12),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_163),
.A2(n_165),
.B(n_166),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_157),
.A2(n_10),
.B(n_6),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g166 ( 
.A(n_155),
.B(n_6),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_158),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_164),
.B(n_156),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_168),
.B(n_169),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_155),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_166),
.C(n_3),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_2),
.C(n_3),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_170),
.A2(n_2),
.B(n_3),
.Y(n_173)
);

AOI322xp5_ASAP7_75t_L g176 ( 
.A1(n_173),
.A2(n_4),
.A3(n_21),
.B1(n_27),
.B2(n_34),
.C1(n_40),
.C2(n_174),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_176),
.Y(n_177)
);

FAx1_ASAP7_75t_SL g178 ( 
.A(n_177),
.B(n_4),
.CI(n_40),
.CON(n_178),
.SN(n_178)
);


endmodule