module fake_jpeg_2510_n_500 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_500);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_500;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_7),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_15),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_56),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_57),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_58),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_26),
.B(n_7),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_59),
.B(n_71),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_60),
.Y(n_185)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx11_ASAP7_75t_L g173 ( 
.A(n_62),
.Y(n_173)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_64),
.Y(n_198)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx11_ASAP7_75t_L g192 ( 
.A(n_65),
.Y(n_192)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_47),
.Y(n_66)
);

CKINVDCx6p67_ASAP7_75t_R g139 ( 
.A(n_66),
.Y(n_139)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_68),
.Y(n_151)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_69),
.Y(n_143)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_70),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_26),
.B(n_6),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_72),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_73),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_28),
.B(n_10),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_74),
.B(n_93),
.Y(n_123)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_75),
.Y(n_180)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_76),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_78),
.Y(n_186)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_79),
.Y(n_160)
);

BUFx24_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_80),
.Y(n_130)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g183 ( 
.A(n_81),
.Y(n_183)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_83),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_84),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVxp33_ASAP7_75t_L g167 ( 
.A(n_86),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_87),
.Y(n_152)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_88),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_89),
.Y(n_194)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_21),
.Y(n_90)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_91),
.Y(n_196)
);

BUFx4f_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_27),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_94),
.Y(n_164)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_95),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_96),
.Y(n_206)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_97),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_21),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_98),
.B(n_99),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_21),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_101),
.Y(n_131)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_23),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_103),
.Y(n_140)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_SL g162 ( 
.A1(n_104),
.A2(n_113),
.B(n_39),
.Y(n_162)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_106),
.Y(n_150)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_41),
.Y(n_106)
);

BUFx24_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_107),
.B(n_119),
.Y(n_175)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_41),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_111),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_109),
.B(n_24),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_46),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_110),
.B(n_112),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_39),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_46),
.Y(n_112)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_25),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_54),
.B(n_10),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_115),
.Y(n_166)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_22),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_22),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_116),
.B(n_117),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_37),
.B(n_18),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_28),
.B(n_5),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_121),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_29),
.B(n_5),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_37),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_120),
.B(n_2),
.Y(n_184)
);

CKINVDCx9p33_ASAP7_75t_R g121 ( 
.A(n_39),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_42),
.A2(n_5),
.B1(n_15),
.B2(n_12),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_122),
.A2(n_34),
.B1(n_51),
.B2(n_36),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_133),
.A2(n_163),
.B1(n_193),
.B2(n_198),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_59),
.B(n_34),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_135),
.B(n_136),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_71),
.B(n_32),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_74),
.B(n_32),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_138),
.B(n_148),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_109),
.A2(n_25),
.B1(n_54),
.B2(n_36),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_141),
.A2(n_145),
.B1(n_146),
.B2(n_155),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_111),
.A2(n_31),
.B1(n_51),
.B2(n_29),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_111),
.A2(n_31),
.B1(n_53),
.B2(n_42),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_52),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_64),
.A2(n_77),
.B1(n_85),
.B2(n_91),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_149),
.A2(n_161),
.B1(n_178),
.B2(n_182),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_92),
.A2(n_53),
.B1(n_52),
.B2(n_50),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_93),
.A2(n_50),
.B1(n_49),
.B2(n_45),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_156),
.B(n_157),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_49),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_158),
.B(n_169),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_57),
.A2(n_58),
.B1(n_60),
.B2(n_89),
.Y(n_161)
);

INVx3_ASAP7_75t_SL g274 ( 
.A(n_162),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_87),
.A2(n_45),
.B1(n_43),
.B2(n_30),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_120),
.B(n_43),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_84),
.A2(n_30),
.B1(n_24),
.B2(n_3),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_170),
.A2(n_181),
.B1(n_195),
.B2(n_197),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_56),
.B(n_12),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_174),
.B(n_176),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_63),
.B(n_12),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_96),
.A2(n_16),
.B1(n_2),
.B2(n_3),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_105),
.B(n_1),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_179),
.B(n_188),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_88),
.A2(n_80),
.B1(n_110),
.B2(n_112),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_98),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_184),
.B(n_201),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_100),
.B(n_2),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_102),
.B(n_4),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_190),
.B(n_191),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_107),
.B(n_4),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_121),
.A2(n_4),
.B1(n_23),
.B2(n_25),
.Y(n_195)
);

AND2x4_ASAP7_75t_L g197 ( 
.A(n_66),
.B(n_101),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_197),
.Y(n_229)
);

AO22x1_ASAP7_75t_SL g201 ( 
.A1(n_106),
.A2(n_103),
.B1(n_101),
.B2(n_61),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_57),
.A2(n_58),
.B1(n_60),
.B2(n_85),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_203),
.A2(n_205),
.B1(n_161),
.B2(n_145),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_114),
.B(n_59),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_204),
.B(n_150),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_114),
.A2(n_122),
.B1(n_119),
.B2(n_71),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_144),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_167),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_208),
.Y(n_303)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_151),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_211),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_139),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_212),
.B(n_244),
.Y(n_283)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_213),
.Y(n_278)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_142),
.Y(n_214)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_214),
.Y(n_287)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_154),
.Y(n_215)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_215),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_217),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_177),
.B(n_128),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_218),
.B(n_219),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_166),
.B(n_123),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_126),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_221),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_197),
.A2(n_195),
.B1(n_180),
.B2(n_181),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_223),
.A2(n_232),
.B1(n_236),
.B2(n_240),
.Y(n_314)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_224),
.Y(n_291)
);

INVx11_ASAP7_75t_L g227 ( 
.A(n_139),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_227),
.Y(n_292)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_134),
.Y(n_228)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_228),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_123),
.B(n_172),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_230),
.B(n_233),
.Y(n_321)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_171),
.Y(n_231)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_231),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_187),
.A2(n_153),
.B1(n_200),
.B2(n_144),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_175),
.B(n_139),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_175),
.B(n_125),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_235),
.B(n_242),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_187),
.A2(n_200),
.B1(n_165),
.B2(n_202),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_127),
.Y(n_237)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_237),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_165),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_238),
.B(n_275),
.Y(n_294)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_143),
.Y(n_239)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_239),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_202),
.A2(n_160),
.B1(n_170),
.B2(n_141),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_143),
.Y(n_241)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_241),
.Y(n_324)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_173),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_168),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_243),
.B(n_245),
.Y(n_280)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_173),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_130),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_246),
.B(n_254),
.Y(n_315)
);

NOR2x1_ASAP7_75t_L g322 ( 
.A(n_247),
.B(n_270),
.Y(n_322)
);

INVx8_ASAP7_75t_L g248 ( 
.A(n_206),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_248),
.B(n_250),
.Y(n_281)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_183),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_206),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_253),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_131),
.B(n_140),
.Y(n_252)
);

MAJx2_ASAP7_75t_L g317 ( 
.A(n_252),
.B(n_273),
.C(n_238),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_183),
.B(n_167),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_129),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_198),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_256),
.Y(n_284)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_201),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_164),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_263),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_258),
.A2(n_225),
.B1(n_274),
.B2(n_247),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_203),
.A2(n_159),
.B1(n_185),
.B2(n_137),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_260),
.A2(n_266),
.B1(n_232),
.B2(n_236),
.Y(n_323)
);

O2A1O1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_146),
.A2(n_155),
.B(n_192),
.C(n_129),
.Y(n_262)
);

OA21x2_ASAP7_75t_L g312 ( 
.A1(n_262),
.A2(n_223),
.B(n_267),
.Y(n_312)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_132),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_132),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_267),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_137),
.A2(n_185),
.B1(n_159),
.B2(n_192),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_186),
.B(n_147),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_186),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_268),
.B(n_276),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_147),
.B(n_152),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_271),
.Y(n_289)
);

AND2x4_ASAP7_75t_L g270 ( 
.A(n_152),
.B(n_194),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_194),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_124),
.B(n_196),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_272),
.B(n_275),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_196),
.B(n_124),
.Y(n_273)
);

INVx4_ASAP7_75t_SL g275 ( 
.A(n_139),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_139),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_273),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_277),
.B(n_296),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_261),
.B(n_226),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_288),
.B(n_309),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_234),
.B(n_265),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_265),
.B(n_209),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_300),
.B(n_302),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_301),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_209),
.B(n_222),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_304),
.A2(n_300),
.B1(n_312),
.B2(n_296),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_274),
.B(n_229),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_305),
.B(n_307),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_259),
.B(n_249),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g354 ( 
.A(n_306),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_220),
.B(n_270),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_270),
.B(n_269),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_270),
.B(n_231),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_310),
.B(n_311),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_210),
.B(n_221),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_312),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_208),
.B(n_207),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_320),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_317),
.B(n_254),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_228),
.B(n_241),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_323),
.A2(n_242),
.B1(n_245),
.B2(n_314),
.Y(n_343)
);

MAJx2_ASAP7_75t_L g325 ( 
.A(n_240),
.B(n_216),
.C(n_217),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_325),
.B(n_314),
.C(n_312),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_285),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_328),
.B(n_331),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_288),
.B(n_224),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_329),
.B(n_361),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_239),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_330),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_227),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_313),
.Y(n_332)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_332),
.Y(n_366)
);

INVx2_ASAP7_75t_SL g333 ( 
.A(n_294),
.Y(n_333)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_333),
.Y(n_390)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_313),
.Y(n_334)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_334),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_284),
.A2(n_262),
.B1(n_216),
.B2(n_271),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_335),
.A2(n_343),
.B1(n_348),
.B2(n_360),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_336),
.B(n_342),
.C(n_351),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_305),
.A2(n_255),
.B(n_248),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_337),
.A2(n_282),
.B(n_280),
.Y(n_364)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_313),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_338),
.Y(n_392)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_311),
.Y(n_340)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_340),
.Y(n_374)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_287),
.Y(n_341)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_341),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_277),
.B(n_251),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_319),
.B(n_283),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_345),
.B(n_350),
.Y(n_373)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_278),
.Y(n_346)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_346),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_304),
.A2(n_297),
.B1(n_325),
.B2(n_290),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_349),
.B(n_359),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_294),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_294),
.A2(n_322),
.B(n_310),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_352),
.A2(n_355),
.B(n_319),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_322),
.A2(n_309),
.B(n_307),
.Y(n_355)
);

NOR2x1_ASAP7_75t_L g358 ( 
.A(n_302),
.B(n_290),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_358),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_303),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_322),
.A2(n_323),
.B1(n_317),
.B2(n_289),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_278),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_293),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_362),
.B(n_292),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_318),
.Y(n_363)
);

CKINVDCx14_ASAP7_75t_R g393 ( 
.A(n_363),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_364),
.A2(n_391),
.B(n_333),
.Y(n_404)
);

OA21x2_ASAP7_75t_L g375 ( 
.A1(n_352),
.A2(n_279),
.B(n_315),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_375),
.B(n_377),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_340),
.B(n_286),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_326),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_378),
.B(n_327),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_342),
.B(n_298),
.C(n_299),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_379),
.B(n_381),
.C(n_388),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_336),
.B(n_298),
.C(n_293),
.Y(n_381)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_383),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_358),
.B(n_281),
.Y(n_384)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_384),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_339),
.B(n_291),
.Y(n_385)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_385),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_386),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_348),
.A2(n_291),
.B1(n_295),
.B2(n_292),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_387),
.A2(n_350),
.B1(n_343),
.B2(n_333),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_347),
.B(n_324),
.C(n_299),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_353),
.B(n_295),
.Y(n_389)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_389),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_344),
.A2(n_303),
.B(n_324),
.Y(n_391)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_392),
.Y(n_395)
);

INVx2_ASAP7_75t_SL g437 ( 
.A(n_395),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_369),
.A2(n_349),
.B1(n_344),
.B2(n_360),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_397),
.A2(n_398),
.B1(n_415),
.B2(n_374),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_369),
.A2(n_387),
.B1(n_372),
.B2(n_368),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g399 ( 
.A(n_370),
.B(n_347),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_399),
.B(n_405),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_393),
.B(n_354),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_400),
.B(n_402),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_393),
.B(n_328),
.Y(n_402)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_403),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_404),
.A2(n_410),
.B(n_390),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_370),
.B(n_356),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_392),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_407),
.B(n_413),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_378),
.B(n_329),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_409),
.B(n_417),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_386),
.A2(n_351),
.B(n_355),
.Y(n_410)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_411),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_372),
.A2(n_356),
.B1(n_357),
.B2(n_327),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_412),
.A2(n_385),
.B1(n_373),
.B2(n_382),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_392),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_391),
.Y(n_414)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_414),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_368),
.A2(n_357),
.B1(n_337),
.B2(n_346),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_373),
.B(n_359),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_371),
.B(n_308),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g432 ( 
.A(n_418),
.B(n_365),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_399),
.B(n_379),
.C(n_381),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_420),
.B(n_423),
.C(n_424),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_405),
.B(n_379),
.C(n_388),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_401),
.B(n_375),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_425),
.B(n_434),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_426),
.B(n_428),
.Y(n_451)
);

AOI322xp5_ASAP7_75t_L g427 ( 
.A1(n_396),
.A2(n_406),
.A3(n_419),
.B1(n_416),
.B2(n_384),
.C1(n_408),
.C2(n_394),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_427),
.B(n_416),
.Y(n_454)
);

AOI321xp33_ASAP7_75t_L g429 ( 
.A1(n_406),
.A2(n_375),
.A3(n_365),
.B1(n_374),
.B2(n_364),
.C(n_388),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_429),
.A2(n_435),
.B(n_438),
.Y(n_455)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_432),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_401),
.B(n_375),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_408),
.A2(n_390),
.B(n_382),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_396),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_436),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_397),
.A2(n_389),
.B1(n_377),
.B2(n_383),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_439),
.B(n_419),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_410),
.B(n_367),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_440),
.B(n_415),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_431),
.B(n_412),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_443),
.B(n_449),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_432),
.Y(n_444)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_444),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_445),
.B(n_452),
.C(n_420),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_446),
.B(n_450),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_422),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_424),
.B(n_398),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_425),
.B(n_394),
.C(n_404),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_453),
.B(n_454),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_421),
.B(n_366),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_456),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_421),
.Y(n_457)
);

NOR3xp33_ASAP7_75t_L g464 ( 
.A(n_457),
.B(n_441),
.C(n_435),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_426),
.B(n_366),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_458),
.B(n_430),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_461),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_451),
.A2(n_430),
.B1(n_428),
.B2(n_439),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_463),
.A2(n_467),
.B1(n_469),
.B2(n_447),
.Y(n_476)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_464),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_445),
.B(n_434),
.C(n_423),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_465),
.B(n_442),
.C(n_450),
.Y(n_479)
);

INVx11_ASAP7_75t_L g466 ( 
.A(n_444),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_466),
.B(n_457),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_455),
.A2(n_438),
.B(n_433),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_468),
.A2(n_446),
.B(n_440),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_455),
.A2(n_433),
.B(n_414),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_471),
.A2(n_456),
.B(n_447),
.Y(n_474)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_472),
.Y(n_488)
);

OAI221xp5_ASAP7_75t_L g473 ( 
.A1(n_462),
.A2(n_429),
.B1(n_453),
.B2(n_458),
.C(n_448),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_473),
.A2(n_474),
.B(n_481),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_476),
.B(n_477),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_470),
.B(n_449),
.Y(n_477)
);

A2O1A1O1Ixp25_ASAP7_75t_L g482 ( 
.A1(n_479),
.A2(n_461),
.B(n_470),
.C(n_451),
.D(n_459),
.Y(n_482)
);

OAI321xp33_ASAP7_75t_L g486 ( 
.A1(n_480),
.A2(n_466),
.A3(n_460),
.B1(n_463),
.B2(n_413),
.C(n_407),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_465),
.B(n_442),
.C(n_452),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_482),
.B(n_479),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_478),
.A2(n_468),
.B(n_471),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_484),
.A2(n_485),
.B(n_486),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_474),
.A2(n_459),
.B(n_469),
.Y(n_485)
);

AOI21x1_ASAP7_75t_L g489 ( 
.A1(n_488),
.A2(n_481),
.B(n_475),
.Y(n_489)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_489),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_490),
.B(n_492),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_487),
.B(n_460),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_491),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_483),
.B(n_361),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_494),
.A2(n_493),
.B1(n_491),
.B2(n_437),
.Y(n_497)
);

AO21x1_ASAP7_75t_L g499 ( 
.A1(n_497),
.A2(n_498),
.B(n_495),
.Y(n_499)
);

NAND3xp33_ASAP7_75t_L g498 ( 
.A(n_496),
.B(n_376),
.C(n_380),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_499),
.B(n_380),
.Y(n_500)
);


endmodule