module fake_jpeg_26292_n_107 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_107);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_107;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_22),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_23),
.B(n_1),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_29),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_1),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

NAND2xp33_ASAP7_75t_SL g33 ( 
.A(n_31),
.B(n_32),
.Y(n_33)
);

BUFx12f_ASAP7_75t_SL g32 ( 
.A(n_22),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_23),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_18),
.Y(n_38)
);

AO22x1_ASAP7_75t_SL g40 ( 
.A1(n_32),
.A2(n_20),
.B1(n_16),
.B2(n_18),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_41),
.B1(n_13),
.B2(n_12),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_24),
.A2(n_11),
.B1(n_13),
.B2(n_12),
.Y(n_41)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_34),
.B(n_28),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_45),
.B(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx2_ASAP7_75t_SL g47 ( 
.A(n_42),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_11),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_49),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_15),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_53),
.B(n_55),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_15),
.Y(n_53)
);

O2A1O1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_33),
.A2(n_32),
.B(n_27),
.C(n_30),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_21),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_57),
.C(n_58),
.Y(n_60)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_57),
.A2(n_33),
.B1(n_40),
.B2(n_30),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_40),
.C(n_25),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_67),
.C(n_36),
.Y(n_76)
);

AO22x1_ASAP7_75t_SL g65 ( 
.A1(n_55),
.A2(n_40),
.B1(n_54),
.B2(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

MAJx2_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_25),
.C(n_26),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_19),
.B(n_21),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_19),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_26),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_76),
.C(n_66),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_73),
.Y(n_83)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_61),
.B(n_68),
.C(n_59),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_74),
.B(n_78),
.Y(n_87)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_60),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_80),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_77),
.A2(n_65),
.B1(n_67),
.B2(n_51),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_75),
.B1(n_31),
.B2(n_16),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_76),
.C(n_71),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_77),
.A2(n_14),
.B1(n_43),
.B2(n_20),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_SL g89 ( 
.A1(n_84),
.A2(n_31),
.B(n_73),
.C(n_49),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_91),
.Y(n_94)
);

AOI21x1_ASAP7_75t_SL g95 ( 
.A1(n_89),
.A2(n_84),
.B(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_92),
.B(n_8),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_1),
.B(n_3),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_96),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_86),
.B(n_3),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_97),
.A2(n_5),
.B(n_6),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_100),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_5),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_10),
.Y(n_104)
);

OAI21x1_ASAP7_75t_L g102 ( 
.A1(n_99),
.A2(n_7),
.B(n_8),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

AOI21x1_ASAP7_75t_L g106 ( 
.A1(n_104),
.A2(n_105),
.B(n_103),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_3),
.Y(n_107)
);


endmodule