module real_jpeg_26563_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_166;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_255;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_228;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_244;
wire n_179;
wire n_216;
wire n_202;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

INVx5_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_1),
.A2(n_43),
.B1(n_44),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_51),
.Y(n_98)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_2),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_3),
.A2(n_74),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_3),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_3),
.A2(n_56),
.B1(n_58),
.B2(n_80),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_3),
.A2(n_43),
.B1(n_44),
.B2(n_80),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_80),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_4),
.A2(n_74),
.B1(n_79),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_4),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_4),
.A2(n_56),
.B1(n_58),
.B2(n_137),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_4),
.A2(n_43),
.B1(n_44),
.B2(n_137),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_137),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_6),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_7),
.A2(n_34),
.B1(n_56),
.B2(n_58),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_7),
.A2(n_34),
.B1(n_43),
.B2(n_44),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_8),
.A2(n_74),
.B1(n_79),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_8),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_8),
.A2(n_56),
.B1(n_58),
.B2(n_112),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_8),
.A2(n_43),
.B1(n_44),
.B2(n_112),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_112),
.Y(n_220)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_9),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_9),
.B(n_77),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_9),
.B(n_58),
.Y(n_179)
);

AOI21xp33_ASAP7_75t_L g183 ( 
.A1(n_9),
.A2(n_58),
.B(n_179),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_9),
.A2(n_43),
.B1(n_44),
.B2(n_126),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_9),
.A2(n_28),
.B(n_47),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_9),
.B(n_59),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_9),
.A2(n_37),
.B1(n_87),
.B2(n_228),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_10),
.A2(n_43),
.B1(n_44),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_10),
.A2(n_49),
.B1(n_56),
.B2(n_58),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_49),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_11),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_12),
.A2(n_39),
.B1(n_74),
.B2(n_79),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_12),
.A2(n_39),
.B1(n_56),
.B2(n_58),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_12),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_149)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_14),
.A2(n_43),
.B1(n_44),
.B2(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_15),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_140),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_138),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_114),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_19),
.B(n_114),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_95),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_83),
.B2(n_84),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_52),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_40),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_24),
.B(n_40),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_35),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_25),
.A2(n_37),
.B(n_128),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_26),
.A2(n_38),
.B(n_100),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_26),
.A2(n_36),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_27),
.A2(n_28),
.B1(n_45),
.B2(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_27),
.B(n_233),
.Y(n_232)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_33),
.B(n_37),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_35),
.A2(n_87),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

INVx5_ASAP7_75t_SL g88 ( 
.A(n_36),
.Y(n_88)
);

INVx11_ASAP7_75t_L g229 ( 
.A(n_36),
.Y(n_229)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_37),
.B(n_126),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_41),
.A2(n_50),
.B(n_91),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_41),
.A2(n_91),
.B(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_41),
.A2(n_46),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_41),
.A2(n_187),
.B(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_41),
.A2(n_46),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_41),
.A2(n_46),
.B1(n_186),
.B2(n_205),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_46),
.Y(n_41)
);

AOI32xp33_ASAP7_75t_L g177 ( 
.A1(n_43),
.A2(n_56),
.A3(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp33_ASAP7_75t_SL g180 ( 
.A(n_44),
.B(n_66),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_L g206 ( 
.A1(n_44),
.A2(n_45),
.B(n_126),
.C(n_207),
.Y(n_206)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_46),
.A2(n_48),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_46),
.B(n_126),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_68),
.B2(n_69),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_59),
.B(n_62),
.Y(n_54)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_58),
.B1(n_61),
.B2(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_58),
.B1(n_72),
.B2(n_73),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_56),
.A2(n_76),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_58),
.B(n_72),
.Y(n_124)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_63),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_60),
.B(n_107),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_60),
.A2(n_64),
.B1(n_131),
.B2(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_60),
.A2(n_64),
.B1(n_152),
.B2(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_60),
.A2(n_64),
.B1(n_165),
.B2(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_66),
.Y(n_178)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_78),
.B(n_81),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_70),
.A2(n_78),
.B1(n_111),
.B2(n_113),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_70),
.A2(n_111),
.B1(n_113),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_71),
.A2(n_77),
.B1(n_125),
.B2(n_136),
.Y(n_153)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_74),
.B(n_76),
.C(n_77),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_74),
.Y(n_76)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

HAxp5_ASAP7_75t_SL g125 ( 
.A(n_74),
.B(n_126),
.CON(n_125),
.SN(n_125)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_77),
.B(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_90),
.B2(n_94),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B(n_89),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_87),
.A2(n_88),
.B1(n_98),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_87),
.A2(n_220),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_90),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_92),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_93),
.B(n_149),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_104),
.C(n_109),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_101),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_97),
.B(n_101),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_104),
.A2(n_109),
.B1(n_110),
.B2(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_104),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B(n_108),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_130),
.B(n_132),
.Y(n_129)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.C(n_120),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_115),
.A2(n_118),
.B1(n_119),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_115),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_120),
.A2(n_121),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_129),
.C(n_133),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_122),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_127),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_129),
.A2(n_133),
.B1(n_134),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_129),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_169),
.B(n_252),
.C(n_258),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_157),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_142),
.B(n_157),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_154),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_144),
.B(n_145),
.C(n_154),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.C(n_153),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_146),
.A2(n_147),
.B1(n_150),
.B2(n_151),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_153),
.B(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.C(n_163),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_158),
.A2(n_159),
.B1(n_247),
.B2(n_249),
.Y(n_246)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_248),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_163),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.C(n_168),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_168),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_251),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_244),
.B(n_250),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_198),
.B(n_243),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_188),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_173),
.B(n_188),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_181),
.C(n_184),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_174),
.A2(n_175),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_177),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_181),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_193),
.B2(n_194),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_189),
.B(n_195),
.C(n_196),
.Y(n_245)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_237),
.B(n_242),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_216),
.B(n_236),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_208),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_201),
.B(n_208),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_206),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_202),
.A2(n_203),
.B1(n_206),
.B2(n_223),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_206),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_214),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_213),
.C(n_214),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_215),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_224),
.B(n_235),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_218),
.B(n_222),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_230),
.B(n_234),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_226),
.B(n_227),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_238),
.B(n_239),
.Y(n_242)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_245),
.B(n_246),
.Y(n_250)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_247),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_253),
.B(n_254),
.Y(n_258)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);


endmodule