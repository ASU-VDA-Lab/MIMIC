module fake_jpeg_14578_n_70 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_70);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_70;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_24;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_67;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_4),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx4f_ASAP7_75t_SL g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_21),
.Y(n_27)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_23),
.Y(n_25)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_18),
.A2(n_13),
.B1(n_9),
.B2(n_10),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_34),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_15),
.C(n_12),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_15),
.C(n_16),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_17),
.Y(n_32)
);

BUFx24_ASAP7_75t_SL g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_10),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_36),
.C(n_15),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_12),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_30),
.A2(n_23),
.B1(n_22),
.B2(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_40),
.Y(n_46)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_43),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_29),
.C(n_20),
.Y(n_50)
);

XNOR2x1_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_19),
.Y(n_47)
);

OA21x2_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_49),
.B(n_46),
.Y(n_54)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_24),
.B(n_16),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_48),
.B(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_53),
.Y(n_58)
);

INVxp33_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_55),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_60),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_51),
.C(n_29),
.Y(n_60)
);

AOI21xp33_ASAP7_75t_SL g61 ( 
.A1(n_57),
.A2(n_56),
.B(n_37),
.Y(n_61)
);

OAI21x1_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_7),
.B(n_2),
.Y(n_64)
);

AO22x1_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_60),
.B1(n_1),
.B2(n_23),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_1),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_64),
.B(n_3),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_2),
.Y(n_66)
);

AO221x1_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_67),
.B1(n_5),
.B2(n_8),
.C(n_29),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_5),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_62),
.Y(n_70)
);


endmodule