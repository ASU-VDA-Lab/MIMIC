module real_jpeg_27437_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_215;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_205;
wire n_110;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_216;
wire n_128;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_0),
.A2(n_35),
.B1(n_41),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_0),
.A2(n_45),
.B1(n_53),
.B2(n_54),
.Y(n_126)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_3),
.A2(n_53),
.B1(n_54),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_3),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_3),
.A2(n_29),
.B1(n_57),
.B2(n_86),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_3),
.A2(n_35),
.B1(n_41),
.B2(n_86),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_5),
.A2(n_35),
.B1(n_41),
.B2(n_124),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_5),
.Y(n_124)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_7),
.A2(n_35),
.B1(n_41),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_7),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_8),
.A2(n_29),
.B1(n_57),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_8),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_8),
.A2(n_30),
.B1(n_60),
.B2(n_70),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_8),
.A2(n_35),
.B1(n_41),
.B2(n_60),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_8),
.A2(n_53),
.B1(n_54),
.B2(n_60),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_9),
.A2(n_27),
.B(n_29),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_9),
.A2(n_25),
.B1(n_30),
.B2(n_70),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_9),
.B(n_54),
.Y(n_153)
);

A2O1A1O1Ixp25_ASAP7_75t_L g155 ( 
.A1(n_9),
.A2(n_54),
.B(n_88),
.C(n_153),
.D(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_9),
.B(n_51),
.Y(n_160)
);

OAI21xp33_ASAP7_75t_L g184 ( 
.A1(n_9),
.A2(n_34),
.B(n_166),
.Y(n_184)
);

A2O1A1O1Ixp25_ASAP7_75t_L g194 ( 
.A1(n_9),
.A2(n_50),
.B(n_57),
.C(n_62),
.D(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_9),
.B(n_57),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_10),
.A2(n_30),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_10),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_10),
.A2(n_29),
.B1(n_57),
.B2(n_69),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_10),
.A2(n_53),
.B1(n_54),
.B2(n_69),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_10),
.A2(n_35),
.B1(n_41),
.B2(n_69),
.Y(n_173)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_11),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_12),
.A2(n_29),
.B1(n_57),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_12),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_12),
.A2(n_30),
.B1(n_64),
.B2(n_70),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_12),
.A2(n_53),
.B1(n_54),
.B2(n_64),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_12),
.A2(n_35),
.B1(n_41),
.B2(n_64),
.Y(n_168)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_14),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_14),
.A2(n_29),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_15),
.A2(n_35),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_15),
.A2(n_42),
.B1(n_53),
.B2(n_54),
.Y(n_93)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_16),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_132),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_130),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_108),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_20),
.B(n_108),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_78),
.C(n_95),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_21),
.B(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_46),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_22),
.B(n_47),
.C(n_77),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_31),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_23),
.A2(n_24),
.B1(n_31),
.B2(n_32),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B(n_28),
.C(n_30),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_25),
.B(n_71),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_25),
.B(n_94),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_25),
.B(n_38),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_57),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_26),
.A2(n_27),
.B1(n_30),
.B2(n_70),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

AOI32xp33_ASAP7_75t_L g202 ( 
.A1(n_29),
.A2(n_54),
.A3(n_195),
.B1(n_203),
.B2(n_205),
.Y(n_202)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_33),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_34),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_34),
.A2(n_81),
.B1(n_82),
.B2(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_34),
.A2(n_40),
.B1(n_81),
.B2(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_34),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_34),
.B(n_168),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_35),
.A2(n_41),
.B1(n_89),
.B2(n_90),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_35),
.B(n_89),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI32xp33_ASAP7_75t_L g152 ( 
.A1(n_41),
.A2(n_53),
.A3(n_90),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_41),
.B(n_186),
.Y(n_185)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_43),
.B(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_44),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_66),
.B2(n_77),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_58),
.B(n_61),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_50),
.A2(n_51),
.B1(n_59),
.B2(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_50),
.B(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_55),
.Y(n_50)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_52),
.Y(n_204)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

NAND2xp33_ASAP7_75t_SL g205 ( 
.A(n_53),
.B(n_204),
.Y(n_205)
);

O2A1O1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_54),
.A2(n_89),
.B(n_91),
.C(n_92),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_54),
.B(n_89),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_65),
.A2(n_118),
.B(n_119),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_65),
.A2(n_107),
.B(n_119),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_66),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_71),
.B(n_73),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_68),
.A2(n_72),
.B1(n_74),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_72),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_72),
.B(n_76),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_76),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_74),
.A2(n_102),
.B(n_103),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_78),
.B(n_95),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_84),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_84),
.Y(n_111)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_81),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_81),
.A2(n_173),
.B(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_87),
.B1(n_93),
.B2(n_94),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_85),
.A2(n_94),
.B(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_87),
.A2(n_93),
.B1(n_94),
.B2(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_87),
.A2(n_215),
.B(n_216),
.Y(n_214)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_88),
.B(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_88),
.A2(n_92),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_94),
.B(n_100),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_94),
.A2(n_98),
.B(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_101),
.C(n_105),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_96),
.A2(n_97),
.B1(n_105),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_101),
.B(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_108)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_121),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_116),
.B2(n_117),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_125),
.Y(n_121)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_127),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_146),
.B(n_223),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_144),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_134),
.B(n_144),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.C(n_139),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_135),
.B(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_138),
.B(n_139),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.C(n_143),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_140),
.B(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_141),
.B(n_143),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_142),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_218),
.B(n_222),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_207),
.B(n_217),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_190),
.B(n_206),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_169),
.B(n_189),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_157),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_151),
.B(n_157),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_155),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_156),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_164),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_159),
.B(n_162),
.C(n_164),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_163),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_165),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_177),
.B(n_188),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_176),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_171),
.B(n_176),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_175),
.A2(n_182),
.B(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_183),
.B(n_187),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_179),
.B(n_180),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_191),
.B(n_192),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_199),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_196),
.C(n_199),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_198),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_202),
.Y(n_213)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_208),
.B(n_209),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_213),
.C(n_214),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_219),
.B(n_220),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);


endmodule