module fake_jpeg_17181_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_10),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_24),
.Y(n_42)
);

AO22x1_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_24),
.B1(n_31),
.B2(n_18),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_16),
.B(n_8),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_16),
.Y(n_45)
);

NAND3xp33_ASAP7_75t_L g93 ( 
.A(n_45),
.B(n_31),
.C(n_32),
.Y(n_93)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_34),
.B1(n_17),
.B2(n_20),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_51),
.A2(n_53),
.B1(n_62),
.B2(n_42),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_34),
.B1(n_24),
.B2(n_18),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_35),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_59),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_34),
.B1(n_20),
.B2(n_18),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_57),
.A2(n_42),
.B1(n_27),
.B2(n_31),
.Y(n_75)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_41),
.B(n_24),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_20),
.B1(n_24),
.B2(n_28),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_30),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_23),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_27),
.Y(n_69)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_69),
.B(n_70),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_28),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_71),
.B(n_76),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_72),
.Y(n_126)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_75),
.A2(n_100),
.B1(n_103),
.B2(n_58),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_56),
.B(n_19),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_49),
.Y(n_80)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_19),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_82),
.Y(n_119)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_35),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_84),
.B(n_91),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_85),
.B(n_90),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_87),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_88),
.Y(n_123)
);

OR2x2_ASAP7_75t_SL g90 ( 
.A(n_59),
.B(n_31),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_35),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_48),
.A2(n_31),
.B(n_26),
.C(n_27),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_92),
.A2(n_99),
.B(n_101),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_93),
.Y(n_127)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_50),
.B(n_26),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_97),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_48),
.A2(n_40),
.B1(n_38),
.B2(n_36),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_52),
.A2(n_33),
.B1(n_32),
.B2(n_22),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_54),
.A2(n_40),
.B1(n_38),
.B2(n_21),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_25),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_102),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_52),
.A2(n_33),
.B1(n_22),
.B2(n_7),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_53),
.A2(n_40),
.B1(n_38),
.B2(n_25),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

FAx1_ASAP7_75t_SL g105 ( 
.A(n_46),
.B(n_43),
.CI(n_23),
.CON(n_105),
.SN(n_105)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_66),
.C(n_43),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_108),
.Y(n_157)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_80),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_111),
.B(n_124),
.Y(n_139)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_116),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_84),
.B(n_43),
.C(n_46),
.Y(n_124)
);

O2A1O1Ixp33_ASAP7_75t_SL g125 ( 
.A1(n_71),
.A2(n_73),
.B(n_91),
.C(n_105),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_125),
.A2(n_83),
.B(n_79),
.Y(n_151)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_86),
.B(n_23),
.C(n_25),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_82),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_120),
.A2(n_73),
.B(n_69),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_130),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_121),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_136),
.B(n_140),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_112),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_106),
.A2(n_86),
.B1(n_87),
.B2(n_105),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_141),
.A2(n_145),
.B1(n_154),
.B2(n_165),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_112),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_163),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_106),
.A2(n_58),
.B1(n_67),
.B2(n_61),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_143),
.A2(n_108),
.B1(n_128),
.B2(n_123),
.Y(n_178)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_122),
.A2(n_86),
.B1(n_104),
.B2(n_90),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_95),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_146),
.B(n_152),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_127),
.A2(n_122),
.B1(n_129),
.B2(n_120),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_148),
.A2(n_166),
.B1(n_109),
.B2(n_113),
.Y(n_188)
);

AOI22x1_ASAP7_75t_SL g150 ( 
.A1(n_125),
.A2(n_92),
.B1(n_70),
.B2(n_97),
.Y(n_150)
);

OAI211xp5_ASAP7_75t_L g175 ( 
.A1(n_150),
.A2(n_145),
.B(n_141),
.C(n_165),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_151),
.B(n_117),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_110),
.B(n_78),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_99),
.B1(n_101),
.B2(n_79),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_153),
.A2(n_160),
.B1(n_123),
.B2(n_132),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_111),
.A2(n_83),
.B1(n_85),
.B2(n_96),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_89),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_156),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_89),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_94),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_161),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_127),
.A2(n_29),
.B(n_25),
.C(n_14),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_114),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_88),
.Y(n_164)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_125),
.A2(n_77),
.B1(n_63),
.B2(n_88),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_134),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_170),
.B(n_171),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_151),
.A2(n_113),
.B(n_121),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_173),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_110),
.C(n_126),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_174),
.B(n_29),
.C(n_157),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_154),
.Y(n_209)
);

BUFx8_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_176),
.Y(n_203)
);

NOR2x1_ASAP7_75t_R g177 ( 
.A(n_150),
.B(n_129),
.Y(n_177)
);

MAJx2_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_139),
.C(n_160),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_191),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_158),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_179),
.B(n_180),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_152),
.B(n_118),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_158),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_183),
.B(n_188),
.Y(n_225)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_138),
.Y(n_185)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_190),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_149),
.Y(n_191)
);

BUFx24_ASAP7_75t_SL g192 ( 
.A(n_156),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_193),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_149),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_196),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_148),
.B(n_114),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_155),
.Y(n_205)
);

NAND3xp33_ASAP7_75t_SL g196 ( 
.A(n_166),
.B(n_135),
.C(n_161),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_147),
.A2(n_116),
.B1(n_118),
.B2(n_25),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_198),
.A2(n_137),
.B1(n_116),
.B2(n_157),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_153),
.B1(n_147),
.B2(n_160),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_200),
.A2(n_212),
.B1(n_219),
.B2(n_181),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_201),
.A2(n_216),
.B1(n_188),
.B2(n_179),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_205),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_163),
.Y(n_207)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_170),
.Y(n_231)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_187),
.A2(n_136),
.B1(n_142),
.B2(n_140),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_226),
.C(n_168),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_186),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_217),
.B(n_224),
.Y(n_239)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_169),
.Y(n_218)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_187),
.A2(n_137),
.B1(n_1),
.B2(n_2),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_168),
.B(n_29),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_171),
.B(n_30),
.Y(n_226)
);

AOI22x1_ASAP7_75t_L g227 ( 
.A1(n_220),
.A2(n_173),
.B1(n_177),
.B2(n_195),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_227),
.A2(n_234),
.B1(n_241),
.B2(n_221),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_223),
.A2(n_194),
.B1(n_182),
.B2(n_197),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_228),
.A2(n_205),
.B1(n_204),
.B2(n_201),
.Y(n_249)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_229),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_206),
.Y(n_230)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_230),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_209),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_167),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_235),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_174),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_244),
.C(n_245),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_207),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_206),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_238),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_182),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_225),
.A2(n_202),
.B1(n_200),
.B2(n_212),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_210),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_243),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_172),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_181),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_246),
.A2(n_248),
.B1(n_239),
.B2(n_238),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_183),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_249),
.B(n_236),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_0),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_247),
.A2(n_214),
.B1(n_204),
.B2(n_208),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_253),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_213),
.C(n_226),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_260),
.C(n_262),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_261),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_227),
.A2(n_211),
.B1(n_208),
.B2(n_216),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_258),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_211),
.C(n_190),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_198),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_228),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_227),
.B(n_189),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_266),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_185),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_268),
.A2(n_274),
.B1(n_276),
.B2(n_279),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_251),
.A2(n_236),
.B(n_242),
.Y(n_270)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_270),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_242),
.Y(n_271)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_255),
.A2(n_243),
.B1(n_240),
.B2(n_176),
.Y(n_274)
);

A2O1A1O1Ixp25_ASAP7_75t_L g275 ( 
.A1(n_265),
.A2(n_240),
.B(n_176),
.C(n_30),
.D(n_9),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_266),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_7),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_278),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_257),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_264),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_281),
.A2(n_10),
.B1(n_13),
.B2(n_12),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_274),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_284),
.Y(n_295)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_283),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_252),
.C(n_260),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_256),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_286),
.C(n_294),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

OAI21xp33_ASAP7_75t_L g287 ( 
.A1(n_272),
.A2(n_262),
.B(n_261),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_287),
.A2(n_9),
.B(n_11),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_290),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_252),
.C(n_254),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_9),
.Y(n_294)
);

OAI21x1_ASAP7_75t_L g296 ( 
.A1(n_287),
.A2(n_280),
.B(n_269),
.Y(n_296)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_296),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_282),
.A2(n_278),
.B1(n_272),
.B2(n_269),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_297),
.Y(n_307)
);

OAI21x1_ASAP7_75t_L g304 ( 
.A1(n_298),
.A2(n_286),
.B(n_289),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_291),
.A2(n_11),
.B1(n_3),
.B2(n_4),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_302),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_0),
.C(n_3),
.Y(n_302)
);

NOR3x1_ASAP7_75t_SL g310 ( 
.A(n_304),
.B(n_297),
.C(n_299),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_293),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_309),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_292),
.Y(n_309)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_310),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_299),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_312),
.C(n_294),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_306),
.B(n_302),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_314),
.A2(n_313),
.B(n_307),
.Y(n_316)
);

A2O1A1Ixp33_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_315),
.B(n_303),
.C(n_5),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_3),
.B(n_4),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_5),
.Y(n_319)
);

AOI21x1_ASAP7_75t_SL g320 ( 
.A1(n_319),
.A2(n_5),
.B(n_310),
.Y(n_320)
);


endmodule