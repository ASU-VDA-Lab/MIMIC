module real_jpeg_17313_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_578;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_525;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_599;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_325;
wire n_594;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_0),
.A2(n_21),
.B(n_609),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_0),
.B(n_610),
.Y(n_609)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_1),
.Y(n_106)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_1),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_1),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g338 ( 
.A(n_1),
.Y(n_338)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_2),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_2),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_2),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_2),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g188 ( 
.A(n_3),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_3),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g211 ( 
.A(n_3),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_3),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_4),
.A2(n_122),
.B1(n_126),
.B2(n_131),
.Y(n_121)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_4),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_4),
.A2(n_131),
.B1(n_194),
.B2(n_196),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_4),
.A2(n_131),
.B1(n_370),
.B2(n_372),
.Y(n_369)
);

OAI22xp33_ASAP7_75t_SL g593 ( 
.A1(n_4),
.A2(n_131),
.B1(n_245),
.B2(n_594),
.Y(n_593)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_5),
.A2(n_226),
.B1(n_230),
.B2(n_231),
.Y(n_225)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_5),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_5),
.A2(n_230),
.B1(n_250),
.B2(n_255),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_5),
.A2(n_230),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_5),
.A2(n_149),
.B1(n_230),
.B2(n_243),
.Y(n_391)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_6),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_6),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_6),
.Y(n_119)
);

BUFx4f_ASAP7_75t_L g125 ( 
.A(n_6),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_7),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_7),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_7),
.A2(n_72),
.B1(n_280),
.B2(n_282),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_7),
.A2(n_72),
.B1(n_345),
.B2(n_347),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_7),
.A2(n_72),
.B1(n_439),
.B2(n_442),
.Y(n_438)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_8),
.A2(n_112),
.B1(n_115),
.B2(n_116),
.Y(n_111)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_8),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_8),
.A2(n_115),
.B1(n_214),
.B2(n_218),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g350 ( 
.A1(n_8),
.A2(n_115),
.B1(n_351),
.B2(n_354),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g568 ( 
.A1(n_8),
.A2(n_115),
.B1(n_569),
.B2(n_570),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_9),
.A2(n_168),
.B1(n_169),
.B2(n_171),
.Y(n_167)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_9),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_9),
.A2(n_171),
.B1(n_326),
.B2(n_329),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_9),
.A2(n_171),
.B1(n_574),
.B2(n_578),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_10),
.A2(n_156),
.B1(n_160),
.B2(n_161),
.Y(n_155)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_10),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_10),
.A2(n_74),
.B1(n_160),
.B2(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_10),
.A2(n_160),
.B1(n_448),
.B2(n_450),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_SL g459 ( 
.A1(n_10),
.A2(n_160),
.B1(n_460),
.B2(n_463),
.Y(n_459)
);

OAI22xp33_ASAP7_75t_L g30 ( 
.A1(n_11),
.A2(n_31),
.B1(n_36),
.B2(n_37),
.Y(n_30)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_11),
.A2(n_36),
.B1(n_243),
.B2(n_245),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_11),
.A2(n_36),
.B1(n_126),
.B2(n_431),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_11),
.A2(n_36),
.B1(n_526),
.B2(n_529),
.Y(n_525)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_12),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_13),
.B(n_93),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_13),
.A2(n_92),
.B(n_243),
.Y(n_276)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_13),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_13),
.B(n_78),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_13),
.A2(n_104),
.B1(n_483),
.B2(n_485),
.Y(n_482)
);

OAI32xp33_ASAP7_75t_L g498 ( 
.A1(n_13),
.A2(n_499),
.A3(n_501),
.B1(n_504),
.B2(n_509),
.Y(n_498)
);

AOI22xp33_ASAP7_75t_SL g517 ( 
.A1(n_13),
.A2(n_314),
.B1(n_518),
.B2(n_520),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_14),
.A2(n_146),
.B1(n_149),
.B2(n_153),
.Y(n_145)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_14),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_14),
.A2(n_153),
.B1(n_295),
.B2(n_300),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_14),
.A2(n_153),
.B1(n_425),
.B2(n_427),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_14),
.A2(n_153),
.B1(n_461),
.B2(n_484),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_15),
.A2(n_177),
.B1(n_180),
.B2(n_182),
.Y(n_176)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_15),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_15),
.A2(n_182),
.B1(n_378),
.B2(n_381),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_L g599 ( 
.A1(n_15),
.A2(n_182),
.B1(n_351),
.B2(n_600),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g199 ( 
.A(n_16),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_16),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_16),
.Y(n_220)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_16),
.Y(n_229)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_16),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_16),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_16),
.Y(n_508)
);

INVxp33_ASAP7_75t_L g610 ( 
.A(n_17),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_19),
.Y(n_94)
);

BUFx8_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_19),
.Y(n_148)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_19),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_584),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_557),
.B(n_583),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_395),
.B(n_552),
.Y(n_24)
);

NAND3xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_317),
.C(n_359),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_259),
.B(n_287),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_27),
.B(n_259),
.C(n_554),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_162),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_28),
.B(n_163),
.C(n_221),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_80),
.C(n_132),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_29),
.A2(n_132),
.B1(n_133),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_29),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_41),
.B1(n_69),
.B2(n_78),
.Y(n_29)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_30),
.Y(n_274)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_34),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_35),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx2_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_40),
.Y(n_141)
);

INVx3_ASAP7_75t_SL g248 ( 
.A(n_41),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_41),
.A2(n_78),
.B1(n_367),
.B2(n_368),
.Y(n_366)
);

OA21x2_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_51),
.B(n_57),
.Y(n_41)
);

INVxp33_ASAP7_75t_L g509 ( 
.A(n_42),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_48),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_50),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_61),
.B1(n_63),
.B2(n_66),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_61),
.Y(n_195)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_61),
.Y(n_212)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_64),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_65),
.Y(n_217)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_65),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_65),
.Y(n_423)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_65),
.Y(n_453)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_69),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_70),
.Y(n_500)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_71),
.Y(n_519)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AO22x2_ASAP7_75t_L g140 ( 
.A1(n_76),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_140)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_76),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_77),
.Y(n_254)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_77),
.Y(n_299)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_77),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_77),
.Y(n_577)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22x1_ASAP7_75t_SL g246 ( 
.A1(n_79),
.A2(n_247),
.B1(n_248),
.B2(n_249),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_79),
.A2(n_248),
.B1(n_267),
.B2(n_274),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_79),
.A2(n_248),
.B1(n_267),
.B2(n_294),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_79),
.A2(n_248),
.B1(n_249),
.B2(n_350),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_79),
.A2(n_248),
.B1(n_294),
.B2(n_517),
.Y(n_516)
);

OAI22x1_ASAP7_75t_L g572 ( 
.A1(n_79),
.A2(n_248),
.B1(n_369),
.B2(n_573),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_79),
.A2(n_248),
.B1(n_573),
.B2(n_599),
.Y(n_598)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_80),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_103),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_81),
.B(n_103),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_91),
.B1(n_95),
.B2(n_99),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_88),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_90),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_SL g161 ( 
.A(n_93),
.Y(n_161)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_94),
.Y(n_245)
);

AO21x2_ASAP7_75t_L g134 ( 
.A1(n_95),
.A2(n_135),
.B(n_140),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_96),
.Y(n_139)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_110),
.B1(n_120),
.B2(n_121),
.Y(n_103)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_104),
.A2(n_121),
.B1(n_167),
.B2(n_236),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_104),
.A2(n_176),
.B(n_335),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_104),
.A2(n_430),
.B1(n_435),
.B2(n_437),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_104),
.A2(n_459),
.B1(n_483),
.B2(n_489),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.Y(n_104)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_105),
.A2(n_165),
.B1(n_458),
.B2(n_467),
.Y(n_457)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_107),
.A2(n_188),
.B1(n_189),
.B2(n_191),
.Y(n_187)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_107),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_108),
.Y(n_170)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_108),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_111),
.A2(n_165),
.B1(n_306),
.B2(n_312),
.Y(n_305)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_112),
.Y(n_442)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_112),
.Y(n_484)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_114),
.Y(n_190)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI32xp33_ASAP7_75t_L g401 ( 
.A1(n_117),
.A2(n_402),
.A3(n_405),
.B1(n_409),
.B2(n_411),
.Y(n_401)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_119),
.Y(n_168)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_119),
.Y(n_179)
);

INVx5_ASAP7_75t_L g434 ( 
.A(n_119),
.Y(n_434)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_125),
.Y(n_417)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_125),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_130),
.Y(n_311)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_145),
.B1(n_154),
.B2(n_155),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g241 ( 
.A1(n_134),
.A2(n_154),
.B1(n_155),
.B2(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_134),
.A2(n_145),
.B1(n_154),
.B2(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_134),
.A2(n_154),
.B1(n_242),
.B2(n_344),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_134),
.A2(n_154),
.B1(n_344),
.B2(n_391),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_134),
.A2(n_154),
.B1(n_391),
.B2(n_568),
.Y(n_567)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_134),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_140),
.A2(n_591),
.B1(n_592),
.B2(n_593),
.Y(n_590)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_141),
.Y(n_601)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_148),
.Y(n_244)
);

INVx3_ASAP7_75t_SL g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx5_ASAP7_75t_L g346 ( 
.A(n_151),
.Y(n_346)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_151),
.Y(n_348)
);

INVx8_ASAP7_75t_L g596 ( 
.A(n_151),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_154),
.B(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_221),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_183),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_164),
.A2(n_184),
.B(n_200),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_172),
.B2(n_175),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_165),
.A2(n_306),
.B1(n_438),
.B2(n_511),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_168),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx6_ASAP7_75t_L g489 ( 
.A(n_173),
.Y(n_489)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_174),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_179),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_200),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_192),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_185),
.A2(n_201),
.B1(n_213),
.B2(n_225),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_185),
.A2(n_201),
.B1(n_376),
.B2(n_377),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_185),
.A2(n_201),
.B1(n_420),
.B2(n_424),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_185),
.A2(n_201),
.B1(n_424),
.B2(n_447),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_185),
.A2(n_201),
.B1(n_447),
.B2(n_525),
.Y(n_524)
);

OA21x2_ASAP7_75t_L g579 ( 
.A1(n_185),
.A2(n_201),
.B(n_377),
.Y(n_579)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_186),
.A2(n_278),
.B1(n_279),
.B2(n_286),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_186),
.A2(n_193),
.B1(n_278),
.B2(n_325),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_186),
.B(n_314),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_186),
.A2(n_278),
.B1(n_279),
.B2(n_542),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_202),
.Y(n_201)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_188),
.Y(n_191)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_199),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_213),
.Y(n_200)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_201),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_207),
.B1(n_210),
.B2(n_212),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_205),
.Y(n_503)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_211),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_219),
.Y(n_427)
);

BUFx12f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx4_ASAP7_75t_L g383 ( 
.A(n_220),
.Y(n_383)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_220),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_220),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_240),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_222),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_235),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_223),
.A2(n_224),
.B1(n_235),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_225),
.Y(n_286)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_229),
.Y(n_332)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_234),
.Y(n_530)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_236),
.Y(n_312)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_236),
.Y(n_511)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_239),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_246),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_241),
.Y(n_320)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_245),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_246),
.B(n_320),
.C(n_321),
.Y(n_319)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_254),
.Y(n_303)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_263),
.C(n_265),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_260),
.B(n_316),
.Y(n_315)
);

XNOR2x1_ASAP7_75t_L g316 ( 
.A(n_263),
.B(n_265),
.Y(n_316)
);

MAJx2_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_275),
.C(n_277),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_277),
.Y(n_290)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_272),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_275),
.B(n_290),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_315),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_288),
.B(n_315),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_291),
.C(n_292),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_289),
.B(n_549),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_291),
.B(n_292),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_304),
.C(n_313),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_293),
.B(n_536),
.Y(n_535)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx5_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx6_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx6_ASAP7_75t_L g371 ( 
.A(n_299),
.Y(n_371)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_302),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_304),
.A2(n_305),
.B1(n_313),
.B2(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_311),
.Y(n_466)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_313),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_314),
.B(n_410),
.Y(n_409)
);

OAI21xp33_ASAP7_75t_SL g420 ( 
.A1(n_314),
.A2(n_409),
.B(n_421),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_314),
.B(n_477),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_314),
.B(n_505),
.Y(n_504)
);

A2O1A1O1Ixp25_ASAP7_75t_L g552 ( 
.A1(n_317),
.A2(n_359),
.B(n_553),
.C(n_555),
.D(n_556),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_318),
.B(n_358),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_318),
.B(n_358),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_322),
.Y(n_318)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_319),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_340),
.B1(n_356),
.B2(n_357),
.Y(n_322)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_323),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_323),
.B(n_357),
.C(n_394),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_324),
.A2(n_333),
.B1(n_334),
.B2(n_339),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_324),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_324),
.B(n_334),
.Y(n_386)
);

INVxp33_ASAP7_75t_SL g376 ( 
.A(n_325),
.Y(n_376)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_326),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_328),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_332),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_333),
.A2(n_334),
.B1(n_389),
.B2(n_390),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g563 ( 
.A1(n_333),
.A2(n_390),
.B(n_392),
.Y(n_563)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_340),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_341),
.B(n_362),
.C(n_363),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_349),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_343),
.Y(n_363)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_345),
.Y(n_570)
);

INVx6_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_349),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_350),
.Y(n_367)
);

INVx8_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_360),
.B(n_393),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_360),
.B(n_393),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_364),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_361),
.B(n_560),
.C(n_561),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_385),
.Y(n_364)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_365),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_366),
.A2(n_375),
.B(n_384),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_366),
.B(n_375),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_384),
.A2(n_565),
.B1(n_581),
.B2(n_582),
.Y(n_564)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_384),
.Y(n_581)
);

INVxp67_ASAP7_75t_L g560 ( 
.A(n_385),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_386),
.A2(n_387),
.B1(n_388),
.B2(n_392),
.Y(n_385)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_386),
.Y(n_392)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

AOI21x1_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_547),
.B(n_551),
.Y(n_395)
);

OAI21x1_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_532),
.B(n_546),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_398),
.A2(n_494),
.B(n_531),
.Y(n_397)
);

OAI21x1_ASAP7_75t_L g398 ( 
.A1(n_399),
.A2(n_455),
.B(n_493),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_428),
.Y(n_399)
);

OR2x2_ASAP7_75t_L g493 ( 
.A(n_400),
.B(n_428),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_418),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_401),
.A2(n_418),
.B1(n_419),
.B2(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_401),
.Y(n_469)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_414),
.Y(n_411)
);

INVx6_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_443),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_429),
.B(n_445),
.C(n_454),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_430),
.Y(n_467)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_444),
.A2(n_445),
.B1(n_446),
.B2(n_454),
.Y(n_443)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_444),
.Y(n_454)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_456),
.A2(n_470),
.B(n_492),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_468),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_457),
.B(n_468),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_471),
.A2(n_487),
.B(n_491),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_482),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_476),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_480),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_490),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_488),
.B(n_490),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_496),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_495),
.B(n_496),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_514),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_497),
.B(n_515),
.C(n_524),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_498),
.A2(n_510),
.B1(n_512),
.B2(n_513),
.Y(n_497)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_498),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_498),
.B(n_513),
.Y(n_540)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_510),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_515),
.A2(n_516),
.B1(n_523),
.B2(n_524),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx2_ASAP7_75t_SL g521 ( 
.A(n_522),
.Y(n_521)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g542 ( 
.A(n_525),
.Y(n_542)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

NOR2xp67_ASAP7_75t_L g532 ( 
.A(n_533),
.B(n_545),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_533),
.B(n_545),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_534),
.A2(n_535),
.B1(n_538),
.B2(n_539),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_534),
.B(n_541),
.C(n_543),
.Y(n_550)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_540),
.A2(n_541),
.B1(n_543),
.B2(n_544),
.Y(n_539)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_540),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_541),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_548),
.B(n_550),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_548),
.B(n_550),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_559),
.B(n_562),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_559),
.B(n_562),
.Y(n_583)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_563),
.B(n_564),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_563),
.B(n_581),
.C(n_606),
.Y(n_605)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_565),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_565),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_566),
.A2(n_567),
.B1(n_571),
.B2(n_580),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_566),
.B(n_572),
.C(n_579),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_566),
.A2(n_567),
.B1(n_589),
.B2(n_604),
.Y(n_588)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g591 ( 
.A(n_568),
.Y(n_591)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_571),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_572),
.B(n_579),
.Y(n_571)
);

INVx1_ASAP7_75t_SL g574 ( 
.A(n_575),
.Y(n_574)
);

INVx6_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

INVx6_ASAP7_75t_L g576 ( 
.A(n_577),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_579),
.A2(n_598),
.B1(n_602),
.B2(n_603),
.Y(n_597)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_579),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_SL g584 ( 
.A(n_585),
.B(n_607),
.Y(n_584)
);

NOR2x1_ASAP7_75t_L g585 ( 
.A(n_586),
.B(n_605),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_586),
.B(n_605),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_587),
.B(n_588),
.Y(n_586)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_589),
.Y(n_604)
);

XNOR2x1_ASAP7_75t_L g589 ( 
.A(n_590),
.B(n_597),
.Y(n_589)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_595),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_598),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_601),
.Y(n_600)
);

INVxp33_ASAP7_75t_L g607 ( 
.A(n_608),
.Y(n_607)
);


endmodule