module fake_jpeg_11376_n_106 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_106);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_106;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_32),
.A2(n_16),
.B(n_29),
.C(n_28),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_44),
.B(n_37),
.Y(n_60)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_0),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_52),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_50)
);

NOR2x1_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_36),
.Y(n_53)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_1),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_53),
.B(n_63),
.Y(n_68)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_60),
.B(n_62),
.Y(n_69)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_41),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_32),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_34),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_65),
.Y(n_78)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

MAJx2_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_33),
.C(n_45),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_3),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_74),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_63),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_72),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_58),
.B(n_42),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_71),
.B(n_4),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_43),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_41),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_75),
.A2(n_6),
.B(n_7),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_3),
.Y(n_76)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_86),
.C(n_87),
.Y(n_94)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_67),
.B(n_5),
.Y(n_81)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_83),
.B(n_85),
.Y(n_95)
);

AO21x1_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_6),
.B(n_8),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_9),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_84),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_12),
.B(n_13),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_66),
.B(n_17),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_18),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_74),
.B1(n_22),
.B2(n_23),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_93),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_80),
.A2(n_20),
.B1(n_24),
.B2(n_30),
.Y(n_93)
);

HAxp5_ASAP7_75t_SL g97 ( 
.A(n_95),
.B(n_88),
.CON(n_97),
.SN(n_97)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_97),
.B(n_99),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_86),
.C(n_88),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_94),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_101),
.B(n_97),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_90),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

MAJx2_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_96),
.C(n_89),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_91),
.B(n_93),
.Y(n_106)
);


endmodule