module fake_jpeg_13180_n_410 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_410);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_410;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_38),
.B(n_69),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_41),
.Y(n_84)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_44),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

CKINVDCx6p67_ASAP7_75t_R g93 ( 
.A(n_52),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx5_ASAP7_75t_SL g87 ( 
.A(n_54),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_56),
.Y(n_82)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

CKINVDCx9p33_ASAP7_75t_R g81 ( 
.A(n_57),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_59),
.Y(n_94)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_61),
.A2(n_33),
.B1(n_31),
.B2(n_30),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_65),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_64),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_67),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_28),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_21),
.B(n_0),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_71),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_34),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_36),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_78),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_36),
.Y(n_78)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_52),
.B(n_1),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_79),
.B(n_102),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_62),
.A2(n_15),
.B1(n_16),
.B2(n_32),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_83),
.A2(n_19),
.B1(n_22),
.B2(n_25),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_30),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_86),
.B(n_92),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_39),
.A2(n_47),
.B1(n_45),
.B2(n_44),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_90),
.A2(n_99),
.B1(n_31),
.B2(n_33),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_21),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_42),
.A2(n_15),
.B1(n_16),
.B2(n_32),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_96),
.A2(n_97),
.B1(n_46),
.B2(n_25),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_57),
.A2(n_15),
.B1(n_16),
.B2(n_32),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_64),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_103),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_63),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_34),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_69),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_3),
.Y(n_142)
);

NAND2x1_ASAP7_75t_SL g115 ( 
.A(n_87),
.B(n_22),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_115),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_101),
.B(n_67),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_116),
.B(n_125),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_92),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_130),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_74),
.A2(n_19),
.B(n_28),
.C(n_25),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_121),
.A2(n_137),
.B(n_93),
.C(n_103),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_123),
.A2(n_124),
.B1(n_127),
.B2(n_133),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_78),
.A2(n_58),
.B1(n_56),
.B2(n_55),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_28),
.Y(n_125)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_126),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_81),
.A2(n_40),
.B1(n_53),
.B2(n_19),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_128),
.A2(n_147),
.B1(n_91),
.B2(n_88),
.Y(n_168)
);

BUFx6f_ASAP7_75t_SL g129 ( 
.A(n_81),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_129),
.Y(n_178)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_SL g194 ( 
.A1(n_132),
.A2(n_90),
.B(n_93),
.C(n_95),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_86),
.A2(n_65),
.B1(n_22),
.B2(n_27),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_77),
.B(n_1),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_134),
.B(n_144),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_105),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_135),
.B(n_141),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_94),
.A2(n_27),
.B1(n_2),
.B2(n_3),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_136),
.A2(n_140),
.B1(n_150),
.B2(n_151),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_79),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_L g140 ( 
.A1(n_76),
.A2(n_27),
.B1(n_4),
.B2(n_5),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_105),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_152),
.Y(n_160)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_87),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_84),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_145),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_113),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_146),
.B(n_148),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_84),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_79),
.B(n_6),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_94),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_113),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_79),
.B(n_11),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_73),
.B(n_12),
.Y(n_154)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_154),
.A2(n_156),
.A3(n_112),
.B1(n_109),
.B2(n_100),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_91),
.B(n_12),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_13),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_85),
.B(n_13),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_95),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_157),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_162),
.B(n_137),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_163),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_146),
.A2(n_106),
.B1(n_88),
.B2(n_84),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_167),
.A2(n_155),
.B(n_93),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_168),
.B(n_82),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_117),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_182),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_122),
.A2(n_100),
.B1(n_76),
.B2(n_75),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_174),
.A2(n_123),
.B1(n_133),
.B2(n_136),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_177),
.Y(n_235)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_120),
.Y(n_179)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_181),
.Y(n_232)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_131),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_117),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_185),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_130),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_125),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_191),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_189),
.B(n_110),
.Y(n_237)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_139),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_131),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_193),
.Y(n_210)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_143),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_194),
.A2(n_196),
.B1(n_109),
.B2(n_143),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_139),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_115),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_155),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_161),
.B(n_118),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_198),
.B(n_221),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_L g199 ( 
.A1(n_171),
.A2(n_135),
.B1(n_141),
.B2(n_125),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_199),
.A2(n_216),
.B1(n_219),
.B2(n_224),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_183),
.B(n_153),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_202),
.B(n_204),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_184),
.B(n_153),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_188),
.A2(n_124),
.B1(n_144),
.B2(n_129),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_205),
.A2(n_206),
.B1(n_222),
.B2(n_229),
.Y(n_242)
);

INVxp33_ASAP7_75t_SL g207 ( 
.A(n_186),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_207),
.B(n_218),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_209),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_212),
.B(n_223),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_213),
.A2(n_217),
.B(n_231),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_215),
.A2(n_226),
.B1(n_194),
.B2(n_180),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_171),
.A2(n_122),
.B1(n_116),
.B2(n_152),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_195),
.A2(n_138),
.B(n_148),
.C(n_142),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_172),
.A2(n_154),
.B1(n_156),
.B2(n_138),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_164),
.B(n_138),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_227),
.Y(n_251)
);

BUFx24_ASAP7_75t_SL g221 ( 
.A(n_186),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_187),
.A2(n_175),
.B1(n_174),
.B2(n_195),
.Y(n_222)
);

OA22x2_ASAP7_75t_L g223 ( 
.A1(n_162),
.A2(n_121),
.B1(n_157),
.B2(n_115),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_172),
.A2(n_134),
.B1(n_121),
.B2(n_111),
.Y(n_224)
);

AOI21xp33_ASAP7_75t_L g225 ( 
.A1(n_190),
.A2(n_142),
.B(n_150),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_225),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_175),
.A2(n_137),
.B1(n_75),
.B2(n_104),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_151),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_160),
.B(n_80),
.C(n_98),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_220),
.C(n_219),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_160),
.A2(n_104),
.B1(n_111),
.B2(n_119),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_177),
.Y(n_230)
);

INVxp33_ASAP7_75t_L g249 ( 
.A(n_230),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_190),
.A2(n_160),
.B(n_167),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_169),
.B(n_119),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_234),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_169),
.B(n_93),
.Y(n_234)
);

NOR2x1_ASAP7_75t_L g236 ( 
.A(n_177),
.B(n_112),
.Y(n_236)
);

AO22x1_ASAP7_75t_L g270 ( 
.A1(n_236),
.A2(n_178),
.B1(n_158),
.B2(n_82),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_237),
.B(n_173),
.Y(n_272)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_238),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_239),
.B(n_265),
.C(n_271),
.Y(n_276)
);

AND2x6_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_194),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_241),
.B(n_253),
.Y(n_286)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_200),
.Y(n_243)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_243),
.Y(n_293)
);

XOR2x1_ASAP7_75t_SL g283 ( 
.A(n_244),
.B(n_270),
.Y(n_283)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_245),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_227),
.A2(n_194),
.B1(n_179),
.B2(n_111),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_247),
.A2(n_242),
.B1(n_215),
.B2(n_226),
.Y(n_274)
);

CKINVDCx10_ASAP7_75t_R g248 ( 
.A(n_234),
.Y(n_248)
);

INVxp67_ASAP7_75t_SL g290 ( 
.A(n_248),
.Y(n_290)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_250),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_206),
.A2(n_166),
.B1(n_192),
.B2(n_182),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_252),
.A2(n_255),
.B1(n_272),
.B2(n_229),
.Y(n_284)
);

AND2x6_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_80),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_210),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_254),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_198),
.A2(n_166),
.B1(n_173),
.B2(n_180),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_210),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_267),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_201),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_258),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_201),
.Y(n_258)
);

CKINVDCx12_ASAP7_75t_R g262 ( 
.A(n_228),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_262),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_203),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_263),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_202),
.B(n_158),
.C(n_181),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_233),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_204),
.B(n_191),
.C(n_110),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_239),
.B(n_203),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_273),
.B(n_291),
.C(n_292),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_274),
.A2(n_285),
.B1(n_297),
.B2(n_244),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_212),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_277),
.Y(n_319)
);

AOI22x1_ASAP7_75t_L g281 ( 
.A1(n_272),
.A2(n_264),
.B1(n_247),
.B2(n_251),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_281),
.A2(n_300),
.B(n_270),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_248),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_282),
.B(n_289),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_284),
.A2(n_295),
.B1(n_289),
.B2(n_294),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_251),
.A2(n_224),
.B1(n_237),
.B2(n_216),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_254),
.B(n_222),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_223),
.C(n_208),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_223),
.C(n_208),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_261),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_294),
.B(n_261),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_266),
.A2(n_217),
.B1(n_213),
.B2(n_231),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_240),
.B(n_235),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_301),
.C(n_271),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_264),
.A2(n_215),
.B1(n_211),
.B2(n_200),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_259),
.A2(n_236),
.B(n_218),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_240),
.B(n_211),
.C(n_232),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_288),
.Y(n_302)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_302),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_273),
.B(n_246),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_303),
.B(n_309),
.C(n_322),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_279),
.Y(n_305)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_305),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_277),
.A2(n_246),
.B(n_253),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_306),
.A2(n_300),
.B(n_292),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_260),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_307),
.B(n_275),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_276),
.B(n_266),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_280),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_310),
.B(n_325),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_311),
.A2(n_274),
.B1(n_285),
.B2(n_278),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g337 ( 
.A1(n_312),
.A2(n_321),
.B1(n_324),
.B2(n_249),
.Y(n_337)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_288),
.Y(n_313)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_313),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_295),
.A2(n_267),
.B1(n_259),
.B2(n_241),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_314),
.A2(n_286),
.B1(n_283),
.B2(n_281),
.Y(n_340)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_315),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_280),
.B(n_256),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_316),
.B(n_320),
.Y(n_334)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_298),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_317),
.Y(n_329)
);

MAJx2_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_304),
.C(n_325),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_297),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_298),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_276),
.B(n_269),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_323),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_301),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_296),
.B(n_265),
.C(n_249),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_278),
.B(n_245),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_316),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_327),
.B(n_347),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_330),
.B(n_332),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_335),
.B(n_336),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_312),
.A2(n_277),
.B1(n_291),
.B2(n_283),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_337),
.B(n_339),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_340),
.B(n_341),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_322),
.B(n_299),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_303),
.B(n_281),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_343),
.B(n_311),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_320),
.A2(n_290),
.B1(n_293),
.B2(n_299),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_344),
.B(n_326),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_304),
.B(n_270),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_349),
.B(n_351),
.Y(n_367)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_338),
.Y(n_350)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_350),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_346),
.B(n_332),
.Y(n_351)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_338),
.Y(n_353)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_353),
.Y(n_375)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_329),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_354),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_346),
.B(n_309),
.C(n_324),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_355),
.B(n_356),
.C(n_359),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_347),
.B(n_306),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_327),
.B(n_318),
.C(n_319),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_360),
.B(n_330),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_336),
.B(n_314),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_361),
.B(n_362),
.C(n_328),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_331),
.B(n_319),
.C(n_308),
.Y(n_362)
);

FAx1_ASAP7_75t_SL g364 ( 
.A(n_348),
.B(n_343),
.CI(n_334),
.CON(n_364),
.SN(n_364)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_364),
.B(n_238),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_357),
.A2(n_334),
.B1(n_345),
.B2(n_333),
.Y(n_365)
);

OR2x2_ASAP7_75t_L g386 ( 
.A(n_365),
.B(n_370),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_352),
.A2(n_345),
.B1(n_344),
.B2(n_340),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_371),
.B(n_372),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_361),
.A2(n_349),
.B1(n_356),
.B2(n_362),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_358),
.A2(n_315),
.B(n_305),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_373),
.B(n_236),
.Y(n_383)
);

AND2x2_ASAP7_75t_SL g381 ( 
.A(n_374),
.B(n_243),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_359),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_376),
.B(n_342),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_368),
.A2(n_355),
.B(n_351),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_377),
.B(n_379),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_368),
.A2(n_363),
.B(n_328),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_374),
.B(n_363),
.C(n_293),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_380),
.B(n_381),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_382),
.B(n_383),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_384),
.B(n_364),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_372),
.A2(n_159),
.B(n_165),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_385),
.B(n_365),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_367),
.B(n_196),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_387),
.A2(n_370),
.B1(n_373),
.B2(n_366),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_389),
.B(n_391),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_390),
.B(n_393),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_378),
.B(n_381),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_386),
.A2(n_367),
.B1(n_369),
.B2(n_375),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_392),
.Y(n_402)
);

AOI322xp5_ASAP7_75t_L g395 ( 
.A1(n_378),
.A2(n_375),
.A3(n_369),
.B1(n_364),
.B2(n_165),
.C1(n_159),
.C2(n_104),
.Y(n_395)
);

AOI31xp67_ASAP7_75t_L g397 ( 
.A1(n_395),
.A2(n_383),
.A3(n_82),
.B(n_178),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_397),
.B(n_399),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_396),
.B(n_13),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_388),
.B(n_107),
.C(n_13),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_400),
.B(n_14),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_403),
.B(n_398),
.C(n_394),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_401),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_404),
.A2(n_402),
.B(n_392),
.Y(n_407)
);

AOI322xp5_ASAP7_75t_L g408 ( 
.A1(n_406),
.A2(n_407),
.A3(n_402),
.B1(n_405),
.B2(n_393),
.C1(n_107),
.C2(n_14),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_408),
.B(n_14),
.C(n_107),
.Y(n_409)
);

BUFx24_ASAP7_75t_SL g410 ( 
.A(n_409),
.Y(n_410)
);


endmodule