module fake_netlist_6_3377_n_1842 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1842);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1842;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1736;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1828;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_142),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_14),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_76),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_109),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_111),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_128),
.Y(n_181)
);

BUFx2_ASAP7_75t_SL g182 ( 
.A(n_147),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_74),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_39),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_163),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_152),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_91),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_138),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_25),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_86),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_31),
.Y(n_195)
);

INVxp33_ASAP7_75t_R g196 ( 
.A(n_16),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_2),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_13),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_71),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_28),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_47),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_28),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_37),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_23),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_101),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_10),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_29),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_156),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_57),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_169),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_53),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_47),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_56),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g214 ( 
.A(n_174),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_95),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_31),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_127),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_40),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_75),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_102),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_155),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_38),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_117),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_110),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_20),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_107),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_133),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_15),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_72),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_33),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_19),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_40),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_29),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_33),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_77),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_136),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_49),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_63),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_46),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_10),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_41),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_158),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_83),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_73),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_65),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_25),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_145),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_94),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_144),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_113),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_1),
.Y(n_251)
);

BUFx2_ASAP7_75t_SL g252 ( 
.A(n_131),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_80),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_119),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_17),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_22),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_167),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_13),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_151),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_116),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_140),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_123),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_172),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_78),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_148),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_159),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_50),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_165),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_66),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_146),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_8),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_36),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_0),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_43),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_61),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_139),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_68),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_106),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_50),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_143),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_108),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_170),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_32),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_56),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_103),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_17),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_34),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_57),
.Y(n_288)
);

BUFx5_ASAP7_75t_L g289 ( 
.A(n_99),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_104),
.Y(n_290)
);

BUFx5_ASAP7_75t_L g291 ( 
.A(n_46),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_45),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_98),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_3),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_121),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_154),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_129),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_160),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_114),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_100),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_135),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_69),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_14),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_15),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_18),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_7),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_27),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_82),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_93),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_23),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_173),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_92),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_89),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_62),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_4),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_171),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_84),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_5),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_41),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_70),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_30),
.Y(n_321)
);

CKINVDCx6p67_ASAP7_75t_R g322 ( 
.A(n_45),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_34),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_61),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_43),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_4),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_30),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_124),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_53),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_49),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_122),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_63),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_37),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_59),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_54),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_97),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_64),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_134),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_51),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_79),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_141),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_120),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_112),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_132),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_38),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_36),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_125),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_215),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_291),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_291),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_291),
.Y(n_351)
);

BUFx6f_ASAP7_75t_SL g352 ( 
.A(n_214),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_189),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_217),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_291),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_224),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_205),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_291),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_226),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_229),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_235),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_250),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_236),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_291),
.Y(n_364)
);

NOR2xp67_ASAP7_75t_L g365 ( 
.A(n_288),
.B(n_0),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_291),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_257),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_291),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_244),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_329),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_245),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_177),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_249),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_329),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_329),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_329),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_220),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_329),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_212),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_273),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_273),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_253),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_187),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_346),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_346),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_340),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_347),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_335),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_260),
.Y(n_389)
);

NOR2xp67_ASAP7_75t_L g390 ( 
.A(n_319),
.B(n_1),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_300),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_263),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_213),
.Y(n_393)
);

NOR2xp67_ASAP7_75t_L g394 ( 
.A(n_319),
.B(n_2),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_264),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_276),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_278),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_335),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_220),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_185),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_187),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_280),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_306),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_193),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_201),
.Y(n_405)
);

AND2x6_ASAP7_75t_L g406 ( 
.A(n_261),
.B(n_168),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_281),
.Y(n_407)
);

NOR2xp67_ASAP7_75t_L g408 ( 
.A(n_326),
.B(n_3),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_206),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_246),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_L g411 ( 
.A(n_326),
.B(n_5),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_282),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_211),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_218),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_222),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_179),
.B(n_247),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_295),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_296),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_230),
.Y(n_419)
);

INVxp67_ASAP7_75t_SL g420 ( 
.A(n_312),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_203),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_297),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_299),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_261),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_301),
.Y(n_425)
);

INVxp33_ASAP7_75t_SL g426 ( 
.A(n_195),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_241),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_214),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_255),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_256),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_308),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_271),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_272),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_309),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_311),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_370),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_349),
.B(n_259),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_349),
.B(n_259),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_416),
.B(n_420),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_406),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_350),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_350),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_377),
.B(n_293),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_426),
.B(n_293),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_351),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_351),
.B(n_277),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g447 ( 
.A(n_370),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_377),
.B(n_399),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_383),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_399),
.B(n_277),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_374),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_374),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_388),
.B(n_398),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_383),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_388),
.B(n_331),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_355),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_375),
.B(n_175),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_375),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_355),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_401),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_358),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_401),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_398),
.B(n_358),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_406),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_376),
.B(n_331),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_376),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_364),
.Y(n_467)
);

NOR2x1_ASAP7_75t_L g468 ( 
.A(n_424),
.B(n_336),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_353),
.B(n_267),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_378),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_364),
.B(n_336),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_366),
.B(n_176),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_378),
.B(n_175),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_406),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_366),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_368),
.B(n_178),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_368),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_424),
.B(n_180),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_379),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_424),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_406),
.Y(n_481)
);

INVxp33_ASAP7_75t_L g482 ( 
.A(n_403),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_400),
.B(n_180),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_357),
.A2(n_279),
.B1(n_209),
.B2(n_207),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_380),
.Y(n_485)
);

BUFx8_ASAP7_75t_L g486 ( 
.A(n_352),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_406),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_406),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_390),
.B(n_322),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_372),
.B(n_221),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_380),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_406),
.B(n_184),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_381),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_381),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_384),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_394),
.B(n_186),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_384),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_385),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_410),
.B(n_214),
.Y(n_499)
);

AND2x2_ASAP7_75t_SL g500 ( 
.A(n_428),
.B(n_190),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_412),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_385),
.Y(n_502)
);

OA21x2_ASAP7_75t_L g503 ( 
.A1(n_400),
.A2(n_303),
.B(n_287),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_404),
.Y(n_504)
);

OA21x2_ASAP7_75t_L g505 ( 
.A1(n_404),
.A2(n_330),
.B(n_227),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_405),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_405),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_409),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_409),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_408),
.B(n_219),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_411),
.B(n_242),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_413),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_365),
.B(n_322),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_441),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_444),
.B(n_348),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_441),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_441),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_448),
.Y(n_518)
);

AND3x2_ASAP7_75t_L g519 ( 
.A(n_489),
.B(n_248),
.C(n_243),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_496),
.A2(n_182),
.B1(n_252),
.B2(n_429),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_464),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_441),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_442),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_444),
.B(n_354),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_442),
.Y(n_525)
);

NAND2xp33_ASAP7_75t_L g526 ( 
.A(n_464),
.B(n_474),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_475),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_450),
.B(n_413),
.Y(n_528)
);

INVx4_ASAP7_75t_L g529 ( 
.A(n_464),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_442),
.Y(n_530)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_479),
.B(n_421),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_442),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_475),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_475),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_439),
.B(n_356),
.Y(n_535)
);

INVx5_ASAP7_75t_L g536 ( 
.A(n_464),
.Y(n_536)
);

NOR2x1p5_ASAP7_75t_L g537 ( 
.A(n_483),
.B(n_195),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_445),
.Y(n_538)
);

OR2x6_ASAP7_75t_L g539 ( 
.A(n_448),
.B(n_254),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_448),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_489),
.B(n_359),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_464),
.Y(n_542)
);

INVx2_ASAP7_75t_SL g543 ( 
.A(n_448),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_449),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_445),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_445),
.Y(n_546)
);

AND2x6_ASAP7_75t_L g547 ( 
.A(n_464),
.B(n_262),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_479),
.B(n_360),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_477),
.Y(n_549)
);

INVx4_ASAP7_75t_L g550 ( 
.A(n_464),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_443),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_477),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_445),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_477),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_463),
.Y(n_555)
);

INVxp67_ASAP7_75t_SL g556 ( 
.A(n_449),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_450),
.B(n_443),
.Y(n_557)
);

BUFx8_ASAP7_75t_SL g558 ( 
.A(n_501),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_463),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_456),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_456),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_449),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_463),
.B(n_361),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_449),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_464),
.Y(n_565)
);

INVx5_ASAP7_75t_L g566 ( 
.A(n_464),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_439),
.B(n_363),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_456),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_456),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_463),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_459),
.Y(n_571)
);

INVx1_ASAP7_75t_SL g572 ( 
.A(n_469),
.Y(n_572)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_469),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_489),
.B(n_369),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_490),
.B(n_371),
.Y(n_575)
);

OR2x6_ASAP7_75t_L g576 ( 
.A(n_450),
.B(n_265),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_478),
.Y(n_577)
);

BUFx4f_ASAP7_75t_L g578 ( 
.A(n_505),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_443),
.Y(n_579)
);

OAI22xp33_ASAP7_75t_L g580 ( 
.A1(n_513),
.A2(n_202),
.B1(n_307),
.B2(n_332),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_443),
.B(n_373),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_459),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_459),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_450),
.B(n_414),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_472),
.B(n_476),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_449),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_464),
.Y(n_587)
);

BUFx8_ASAP7_75t_SL g588 ( 
.A(n_501),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_459),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_490),
.B(n_382),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_474),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_483),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_461),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_461),
.Y(n_594)
);

NAND3xp33_ASAP7_75t_L g595 ( 
.A(n_505),
.B(n_415),
.C(n_414),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_461),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_449),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_472),
.B(n_389),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_461),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_478),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_467),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_455),
.B(n_453),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_467),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_467),
.Y(n_604)
);

OR2x2_ASAP7_75t_L g605 ( 
.A(n_457),
.B(n_473),
.Y(n_605)
);

OA22x2_ASAP7_75t_L g606 ( 
.A1(n_455),
.A2(n_415),
.B1(n_433),
.B2(n_432),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_513),
.B(n_392),
.Y(n_607)
);

AO22x1_ASAP7_75t_L g608 ( 
.A1(n_496),
.A2(n_321),
.B1(n_197),
.B2(n_198),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_492),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_467),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_513),
.B(n_395),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_436),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_503),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_503),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_449),
.Y(n_615)
);

INVxp67_ASAP7_75t_SL g616 ( 
.A(n_449),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_455),
.B(n_419),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_486),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_500),
.B(n_396),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_482),
.B(n_397),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_496),
.A2(n_419),
.B1(n_433),
.B2(n_432),
.Y(n_621)
);

OAI22xp33_ASAP7_75t_L g622 ( 
.A1(n_482),
.A2(n_237),
.B1(n_216),
.B2(n_225),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_499),
.B(n_402),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_496),
.A2(n_427),
.B1(n_430),
.B2(n_352),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_492),
.Y(n_625)
);

AND2x2_ASAP7_75t_SL g626 ( 
.A(n_500),
.B(n_266),
.Y(n_626)
);

OR2x6_ASAP7_75t_L g627 ( 
.A(n_499),
.B(n_285),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_457),
.B(n_473),
.Y(n_628)
);

OAI22xp33_ASAP7_75t_SL g629 ( 
.A1(n_492),
.A2(n_313),
.B1(n_316),
.B2(n_302),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_474),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_474),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_436),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_SL g633 ( 
.A1(n_500),
.A2(n_352),
.B1(n_393),
.B2(n_362),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_503),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_472),
.B(n_407),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_449),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_436),
.Y(n_637)
);

OR2x6_ASAP7_75t_L g638 ( 
.A(n_453),
.B(n_290),
.Y(n_638)
);

NAND3xp33_ASAP7_75t_L g639 ( 
.A(n_505),
.B(n_430),
.C(n_427),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_474),
.Y(n_640)
);

NOR3xp33_ASAP7_75t_L g641 ( 
.A(n_484),
.B(n_223),
.C(n_344),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_451),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_500),
.B(n_417),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_503),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_496),
.B(n_418),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_451),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_451),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_503),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_472),
.B(n_422),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_452),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_476),
.B(n_425),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_486),
.B(n_431),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_496),
.B(n_434),
.Y(n_653)
);

BUFx10_ASAP7_75t_L g654 ( 
.A(n_492),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_503),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_486),
.B(n_435),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_484),
.A2(n_204),
.B1(n_345),
.B2(n_339),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_503),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_452),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_476),
.B(n_342),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_505),
.Y(n_661)
);

BUFx2_ASAP7_75t_L g662 ( 
.A(n_505),
.Y(n_662)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_453),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_452),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_486),
.B(n_391),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_555),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_592),
.B(n_423),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_585),
.A2(n_487),
.B(n_481),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_514),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_579),
.B(n_476),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_579),
.B(n_474),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_609),
.B(n_474),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_592),
.B(n_496),
.Y(n_673)
);

NAND3xp33_ASAP7_75t_L g674 ( 
.A(n_535),
.B(n_511),
.C(n_510),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_605),
.B(n_510),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_605),
.B(n_510),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_628),
.B(n_510),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_514),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_555),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_521),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_628),
.B(n_510),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_600),
.B(n_510),
.Y(n_682)
);

A2O1A1Ixp33_ASAP7_75t_L g683 ( 
.A1(n_559),
.A2(n_481),
.B(n_487),
.C(n_492),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_516),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_516),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_531),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_SL g687 ( 
.A1(n_626),
.A2(n_484),
.B1(n_386),
.B2(n_387),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_600),
.B(n_577),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_609),
.B(n_474),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_567),
.B(n_510),
.Y(n_690)
);

HB1xp67_ASAP7_75t_L g691 ( 
.A(n_551),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_517),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_625),
.B(n_474),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_559),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_570),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_575),
.B(n_511),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_521),
.Y(n_697)
);

OAI22xp33_ASAP7_75t_L g698 ( 
.A1(n_657),
.A2(n_437),
.B1(n_438),
.B2(n_200),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_570),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_518),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_517),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_518),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_590),
.B(n_511),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_540),
.B(n_455),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_557),
.B(n_511),
.Y(n_705)
);

INVxp67_ASAP7_75t_L g706 ( 
.A(n_531),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_557),
.B(n_511),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_602),
.B(n_511),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_620),
.B(n_367),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_540),
.Y(n_710)
);

O2A1O1Ixp33_ASAP7_75t_L g711 ( 
.A1(n_663),
.A2(n_438),
.B(n_437),
.C(n_446),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_602),
.B(n_511),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_SL g713 ( 
.A(n_618),
.B(n_486),
.Y(n_713)
);

OAI21xp5_ASAP7_75t_L g714 ( 
.A1(n_578),
.A2(n_487),
.B(n_481),
.Y(n_714)
);

NAND3xp33_ASAP7_75t_L g715 ( 
.A(n_524),
.B(n_486),
.C(n_231),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_543),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_522),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_625),
.B(n_474),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_626),
.A2(n_492),
.B1(n_471),
.B2(n_481),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_543),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_522),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_598),
.B(n_471),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_617),
.Y(n_723)
);

NOR2x1_ASAP7_75t_L g724 ( 
.A(n_623),
.B(n_437),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_563),
.B(n_438),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_617),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_638),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_523),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_635),
.B(n_649),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_626),
.A2(n_492),
.B1(n_471),
.B2(n_481),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_662),
.A2(n_505),
.B1(n_471),
.B2(n_488),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_528),
.B(n_504),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_523),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_548),
.B(n_469),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_662),
.A2(n_505),
.B1(n_488),
.B2(n_440),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_651),
.B(n_507),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_645),
.B(n_507),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_584),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_584),
.Y(n_739)
);

INVx8_ASAP7_75t_L g740 ( 
.A(n_539),
.Y(n_740)
);

NOR3xp33_ASAP7_75t_L g741 ( 
.A(n_619),
.B(n_512),
.C(n_504),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_548),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_527),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_653),
.B(n_660),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_527),
.B(n_507),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_525),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_613),
.A2(n_488),
.B1(n_440),
.B2(n_487),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_515),
.B(n_181),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_533),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_533),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_638),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_581),
.B(n_181),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_578),
.B(n_488),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_574),
.B(n_183),
.Y(n_754)
);

NAND2xp33_ASAP7_75t_L g755 ( 
.A(n_521),
.B(n_488),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_534),
.Y(n_756)
);

A2O1A1Ixp33_ASAP7_75t_L g757 ( 
.A1(n_578),
.A2(n_487),
.B(n_481),
.C(n_440),
.Y(n_757)
);

BUFx5_ASAP7_75t_L g758 ( 
.A(n_661),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_549),
.B(n_507),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_549),
.B(n_552),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_607),
.B(n_183),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_613),
.A2(n_488),
.B1(n_440),
.B2(n_487),
.Y(n_762)
);

AND2x6_ASAP7_75t_L g763 ( 
.A(n_614),
.B(n_488),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_552),
.B(n_507),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_614),
.A2(n_488),
.B1(n_446),
.B2(n_512),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_624),
.B(n_488),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_554),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_554),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_643),
.B(n_188),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_556),
.B(n_446),
.Y(n_770)
);

INVx8_ASAP7_75t_L g771 ( 
.A(n_539),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_612),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_616),
.B(n_447),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_521),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_634),
.B(n_447),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_634),
.B(n_447),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_644),
.B(n_447),
.Y(n_777)
);

INVx1_ASAP7_75t_SL g778 ( 
.A(n_558),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_644),
.B(n_449),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_521),
.B(n_565),
.Y(n_780)
);

INVxp67_ASAP7_75t_SL g781 ( 
.A(n_565),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_612),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_632),
.Y(n_783)
);

INVxp67_ASAP7_75t_L g784 ( 
.A(n_537),
.Y(n_784)
);

OR2x6_ASAP7_75t_L g785 ( 
.A(n_665),
.B(n_196),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_632),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_565),
.B(n_488),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_537),
.B(n_504),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_648),
.B(n_462),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_565),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_519),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_648),
.B(n_462),
.Y(n_792)
);

NOR3xp33_ASAP7_75t_L g793 ( 
.A(n_580),
.B(n_512),
.C(n_238),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_541),
.B(n_191),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_637),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_637),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_565),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_611),
.B(n_192),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_587),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_655),
.B(n_462),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_655),
.B(n_462),
.Y(n_801)
);

NOR2xp67_ASAP7_75t_SL g802 ( 
.A(n_587),
.B(n_591),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_525),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_530),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_627),
.B(n_192),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_587),
.B(n_187),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_530),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_658),
.B(n_661),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_587),
.B(n_187),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_658),
.B(n_462),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_532),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_627),
.A2(n_343),
.B1(n_341),
.B2(n_337),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_520),
.B(n_462),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_532),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_642),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_544),
.B(n_462),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_627),
.B(n_194),
.Y(n_817)
);

AND2x6_ASAP7_75t_SL g818 ( 
.A(n_539),
.B(n_298),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_622),
.B(n_194),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_587),
.B(n_187),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_544),
.B(n_462),
.Y(n_821)
);

NOR2xp67_ASAP7_75t_L g822 ( 
.A(n_595),
.B(n_494),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_591),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_544),
.B(n_462),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_562),
.B(n_462),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_591),
.B(n_187),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_538),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_562),
.B(n_454),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_642),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_638),
.B(n_199),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_562),
.B(n_454),
.Y(n_831)
);

A2O1A1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_725),
.A2(n_595),
.B(n_639),
.C(n_641),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_725),
.B(n_638),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_770),
.A2(n_542),
.B(n_529),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_729),
.B(n_657),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_744),
.B(n_638),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_716),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_755),
.A2(n_542),
.B(n_529),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_680),
.Y(n_839)
);

NAND2x1p5_ASAP7_75t_L g840 ( 
.A(n_704),
.B(n_591),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_716),
.Y(n_841)
);

AO21x1_ASAP7_75t_L g842 ( 
.A1(n_690),
.A2(n_629),
.B(n_652),
.Y(n_842)
);

A2O1A1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_690),
.A2(n_639),
.B(n_526),
.C(n_656),
.Y(n_843)
);

INVxp67_ASAP7_75t_L g844 ( 
.A(n_686),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_735),
.A2(n_576),
.B1(n_539),
.B2(n_633),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_724),
.B(n_591),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_696),
.B(n_576),
.Y(n_847)
);

A2O1A1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_696),
.A2(n_621),
.B(n_328),
.C(n_338),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_758),
.B(n_630),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_781),
.A2(n_542),
.B(n_529),
.Y(n_850)
);

OAI21xp5_ASAP7_75t_L g851 ( 
.A1(n_808),
.A2(n_542),
.B(n_529),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_703),
.B(n_576),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_680),
.A2(n_631),
.B(n_550),
.Y(n_853)
);

INVxp67_ASAP7_75t_L g854 ( 
.A(n_673),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_704),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_680),
.A2(n_774),
.B(n_697),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_L g857 ( 
.A1(n_735),
.A2(n_576),
.B1(n_539),
.B2(n_631),
.Y(n_857)
);

O2A1O1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_698),
.A2(n_629),
.B(n_576),
.C(n_659),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_758),
.B(n_630),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_666),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_703),
.B(n_630),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_722),
.B(n_673),
.Y(n_862)
);

INVxp67_ASAP7_75t_L g863 ( 
.A(n_691),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_758),
.B(n_630),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_742),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_758),
.B(n_630),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_754),
.B(n_640),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_688),
.B(n_608),
.Y(n_868)
);

AO21x1_ASAP7_75t_L g869 ( 
.A1(n_761),
.A2(n_647),
.B(n_646),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_680),
.A2(n_631),
.B(n_550),
.Y(n_870)
);

A2O1A1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_761),
.A2(n_664),
.B(n_650),
.C(n_647),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_697),
.A2(n_631),
.B(n_550),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_675),
.B(n_640),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_757),
.A2(n_731),
.B(n_668),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_698),
.A2(n_547),
.B1(n_606),
.B2(n_664),
.Y(n_875)
);

AOI21x1_ASAP7_75t_L g876 ( 
.A1(n_753),
.A2(n_582),
.B(n_571),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_SL g877 ( 
.A(n_778),
.B(n_588),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_700),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_702),
.Y(n_879)
);

INVxp67_ASAP7_75t_L g880 ( 
.A(n_691),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_697),
.A2(n_550),
.B(n_640),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_676),
.B(n_640),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_758),
.B(n_640),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_706),
.B(n_608),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_L g885 ( 
.A1(n_747),
.A2(n_564),
.B1(n_636),
.B2(n_615),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_697),
.A2(n_566),
.B(n_536),
.Y(n_886)
);

A2O1A1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_769),
.A2(n_586),
.B(n_636),
.C(n_615),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_677),
.B(n_564),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_679),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_710),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_747),
.A2(n_564),
.B1(n_597),
.B2(n_593),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_681),
.B(n_748),
.Y(n_892)
);

OAI21xp33_ASAP7_75t_L g893 ( 
.A1(n_819),
.A2(n_198),
.B(n_197),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_694),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_682),
.B(n_597),
.Y(n_895)
);

OR2x2_ASAP7_75t_SL g896 ( 
.A(n_734),
.B(n_687),
.Y(n_896)
);

O2A1O1Ixp5_ASAP7_75t_L g897 ( 
.A1(n_737),
.A2(n_546),
.B(n_610),
.C(n_538),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_667),
.B(n_573),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_667),
.B(n_572),
.Y(n_899)
);

AOI21xp33_ASAP7_75t_L g900 ( 
.A1(n_794),
.A2(n_572),
.B(n_606),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_720),
.B(n_583),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_774),
.A2(n_566),
.B(n_536),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_732),
.B(n_695),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_752),
.B(n_654),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_723),
.B(n_606),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_699),
.B(n_583),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_774),
.A2(n_566),
.B(n_536),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_774),
.A2(n_566),
.B(n_536),
.Y(n_908)
);

OAI21xp5_ASAP7_75t_L g909 ( 
.A1(n_731),
.A2(n_596),
.B(n_593),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_758),
.B(n_654),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_752),
.B(n_654),
.Y(n_911)
);

CKINVDCx10_ASAP7_75t_R g912 ( 
.A(n_785),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_819),
.B(n_654),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_790),
.A2(n_566),
.B(n_536),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_790),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_794),
.A2(n_596),
.B(n_599),
.C(n_603),
.Y(n_916)
);

AOI21xp33_ASAP7_75t_L g917 ( 
.A1(n_798),
.A2(n_232),
.B(n_228),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_743),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_790),
.A2(n_536),
.B(n_566),
.Y(n_919)
);

OAI21xp33_ASAP7_75t_L g920 ( 
.A1(n_798),
.A2(n_321),
.B(n_209),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_736),
.B(n_599),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_790),
.A2(n_610),
.B(n_604),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_670),
.B(n_603),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_799),
.A2(n_604),
.B(n_601),
.Y(n_924)
);

INVx4_ASAP7_75t_L g925 ( 
.A(n_799),
.Y(n_925)
);

O2A1O1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_711),
.A2(n_601),
.B(n_594),
.C(n_589),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_726),
.B(n_208),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_799),
.A2(n_594),
.B(n_589),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_765),
.B(n_545),
.Y(n_929)
);

O2A1O1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_705),
.A2(n_569),
.B(n_568),
.C(n_561),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_799),
.A2(n_569),
.B(n_568),
.Y(n_931)
);

AND2x2_ASAP7_75t_SL g932 ( 
.A(n_805),
.B(n_465),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_779),
.A2(n_561),
.B(n_560),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_762),
.A2(n_337),
.B1(n_268),
.B2(n_269),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_683),
.A2(n_553),
.B(n_545),
.Y(n_935)
);

NOR3xp33_ASAP7_75t_L g936 ( 
.A(n_784),
.B(n_269),
.C(n_268),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_762),
.A2(n_270),
.B1(n_210),
.B2(n_317),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_765),
.B(n_547),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_789),
.A2(n_460),
.B(n_454),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_674),
.A2(n_547),
.B1(n_465),
.B2(n_270),
.Y(n_940)
);

AOI22xp5_ASAP7_75t_L g941 ( 
.A1(n_708),
.A2(n_547),
.B1(n_465),
.B2(n_317),
.Y(n_941)
);

AOI21x1_ASAP7_75t_L g942 ( 
.A1(n_802),
.A2(n_466),
.B(n_470),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_712),
.B(n_547),
.Y(n_943)
);

NOR3xp33_ASAP7_75t_L g944 ( 
.A(n_817),
.B(n_210),
.C(n_320),
.Y(n_944)
);

O2A1O1Ixp5_ASAP7_75t_L g945 ( 
.A1(n_760),
.A2(n_465),
.B(n_470),
.C(n_466),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_749),
.B(n_547),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_788),
.A2(n_547),
.B1(n_465),
.B2(n_343),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_792),
.A2(n_460),
.B(n_454),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_750),
.B(n_756),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_738),
.B(n_233),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_739),
.B(n_320),
.Y(n_951)
);

OR2x6_ASAP7_75t_L g952 ( 
.A(n_740),
.B(n_506),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_797),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_800),
.A2(n_460),
.B(n_454),
.Y(n_954)
);

AOI21x1_ASAP7_75t_L g955 ( 
.A1(n_787),
.A2(n_458),
.B(n_470),
.Y(n_955)
);

NOR3xp33_ASAP7_75t_L g956 ( 
.A(n_817),
.B(n_341),
.C(n_234),
.Y(n_956)
);

INVx11_ASAP7_75t_L g957 ( 
.A(n_763),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_801),
.A2(n_454),
.B(n_460),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_810),
.A2(n_714),
.B(n_780),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_767),
.B(n_465),
.Y(n_960)
);

BUFx10_ASAP7_75t_L g961 ( 
.A(n_830),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_768),
.B(n_465),
.Y(n_962)
);

OAI22x1_ASAP7_75t_L g963 ( 
.A1(n_812),
.A2(n_200),
.B1(n_345),
.B2(n_339),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_780),
.A2(n_460),
.B(n_480),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_707),
.B(n_506),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_787),
.A2(n_460),
.B(n_480),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_741),
.A2(n_468),
.B1(n_508),
.B2(n_506),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_822),
.B(n_506),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_830),
.B(n_508),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_672),
.A2(n_480),
.B(n_468),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_672),
.A2(n_480),
.B(n_468),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_709),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_SL g973 ( 
.A(n_713),
.B(n_204),
.Y(n_973)
);

AO21x1_ASAP7_75t_L g974 ( 
.A1(n_766),
.A2(n_466),
.B(n_458),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_689),
.A2(n_509),
.B(n_508),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_L g976 ( 
.A1(n_719),
.A2(n_509),
.B1(n_187),
.B2(n_289),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_671),
.B(n_485),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_671),
.B(n_485),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_693),
.A2(n_485),
.B(n_498),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_772),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_782),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_783),
.B(n_485),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_727),
.B(n_239),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_718),
.A2(n_773),
.B(n_775),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_727),
.B(n_751),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_786),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_793),
.B(n_207),
.Y(n_987)
);

O2A1O1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_813),
.A2(n_502),
.B(n_497),
.C(n_495),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_795),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_718),
.A2(n_498),
.B(n_493),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_785),
.B(n_315),
.Y(n_991)
);

BUFx8_ASAP7_75t_L g992 ( 
.A(n_791),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_751),
.B(n_240),
.Y(n_993)
);

INVx1_ASAP7_75t_SL g994 ( 
.A(n_785),
.Y(n_994)
);

NOR3xp33_ASAP7_75t_L g995 ( 
.A(n_715),
.B(n_314),
.C(n_258),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_796),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_815),
.B(n_491),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_829),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_669),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_763),
.B(n_491),
.Y(n_1000)
);

OAI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_730),
.A2(n_502),
.B(n_497),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_763),
.B(n_491),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_763),
.B(n_491),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_678),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_763),
.B(n_493),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_776),
.B(n_251),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_777),
.A2(n_498),
.B(n_493),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_745),
.B(n_493),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_797),
.B(n_502),
.Y(n_1009)
);

AOI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_740),
.A2(n_187),
.B1(n_289),
.B2(n_495),
.Y(n_1010)
);

NAND2xp33_ASAP7_75t_L g1011 ( 
.A(n_740),
.B(n_289),
.Y(n_1011)
);

INVxp67_ASAP7_75t_L g1012 ( 
.A(n_759),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_860),
.Y(n_1013)
);

INVx3_ASAP7_75t_SL g1014 ( 
.A(n_865),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_838),
.A2(n_823),
.B(n_816),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_862),
.B(n_823),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_892),
.B(n_764),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_980),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_851),
.A2(n_824),
.B(n_821),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_SL g1020 ( 
.A1(n_904),
.A2(n_827),
.B(n_684),
.C(n_692),
.Y(n_1020)
);

BUFx3_ASAP7_75t_L g1021 ( 
.A(n_992),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_R g1022 ( 
.A(n_973),
.B(n_771),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_861),
.A2(n_825),
.B(n_771),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_855),
.B(n_806),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_876),
.A2(n_831),
.B(n_828),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_889),
.Y(n_1026)
);

A2O1A1Ixp33_ASAP7_75t_SL g1027 ( 
.A1(n_904),
.A2(n_701),
.B(n_728),
.C(n_733),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_867),
.A2(n_771),
.B(n_820),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_894),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_981),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_835),
.B(n_685),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_835),
.A2(n_807),
.B1(n_746),
.B2(n_717),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_854),
.B(n_721),
.Y(n_1033)
);

OAI21xp33_ASAP7_75t_L g1034 ( 
.A1(n_893),
.A2(n_325),
.B(n_318),
.Y(n_1034)
);

O2A1O1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_917),
.A2(n_826),
.B(n_820),
.C(n_806),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_913),
.A2(n_803),
.B1(n_814),
.B2(n_811),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_918),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_853),
.A2(n_826),
.B(n_809),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_913),
.B(n_804),
.Y(n_1039)
);

NOR2xp67_ASAP7_75t_SL g1040 ( 
.A(n_839),
.B(n_809),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_956),
.A2(n_868),
.B1(n_932),
.B2(n_898),
.Y(n_1041)
);

NAND3xp33_ASAP7_75t_SL g1042 ( 
.A(n_956),
.B(n_323),
.C(n_324),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_833),
.B(n_305),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_903),
.B(n_304),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_870),
.A2(n_498),
.B(n_818),
.Y(n_1045)
);

BUFx2_ASAP7_75t_L g1046 ( 
.A(n_844),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_868),
.B(n_294),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_932),
.A2(n_289),
.B1(n_274),
.B2(n_292),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_836),
.A2(n_310),
.B(n_283),
.C(n_284),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_898),
.B(n_275),
.Y(n_1050)
);

NAND2xp33_ASAP7_75t_R g1051 ( 
.A(n_899),
.B(n_334),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_992),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_839),
.Y(n_1053)
);

INVx4_ASAP7_75t_L g1054 ( 
.A(n_839),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_863),
.B(n_880),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_986),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_989),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_961),
.B(n_286),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_854),
.B(n_289),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_844),
.Y(n_1060)
);

INVx4_ASAP7_75t_L g1061 ( 
.A(n_839),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_1012),
.B(n_289),
.Y(n_1062)
);

NOR2xp67_ASAP7_75t_L g1063 ( 
.A(n_878),
.B(n_130),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_863),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_872),
.A2(n_137),
.B(n_81),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_996),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_875),
.A2(n_334),
.B1(n_333),
.B2(n_327),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_972),
.B(n_333),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_998),
.Y(n_1069)
);

O2A1O1Ixp5_ASAP7_75t_L g1070 ( 
.A1(n_869),
.A2(n_289),
.B(n_67),
.C(n_115),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_880),
.B(n_884),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_1009),
.Y(n_1072)
);

NOR3xp33_ASAP7_75t_L g1073 ( 
.A(n_920),
.B(n_327),
.C(n_325),
.Y(n_1073)
);

NOR2xp67_ASAP7_75t_SL g1074 ( 
.A(n_915),
.B(n_324),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_949),
.Y(n_1075)
);

INVx3_ASAP7_75t_L g1076 ( 
.A(n_840),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_873),
.A2(n_105),
.B(n_161),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_882),
.A2(n_96),
.B(n_157),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_912),
.Y(n_1079)
);

CKINVDCx16_ASAP7_75t_R g1080 ( 
.A(n_877),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_R g1081 ( 
.A(n_961),
.B(n_153),
.Y(n_1081)
);

CKINVDCx8_ASAP7_75t_R g1082 ( 
.A(n_884),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_879),
.B(n_150),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_875),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_915),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_R g1086 ( 
.A(n_837),
.B(n_118),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_834),
.A2(n_90),
.B(n_88),
.Y(n_1087)
);

INVx4_ASAP7_75t_L g1088 ( 
.A(n_915),
.Y(n_1088)
);

O2A1O1Ixp5_ASAP7_75t_L g1089 ( 
.A1(n_842),
.A2(n_289),
.B(n_87),
.C(n_85),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_950),
.B(n_9),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1012),
.B(n_11),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_896),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_901),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_900),
.B(n_11),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_841),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_944),
.B(n_12),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1009),
.Y(n_1097)
);

INVx1_ASAP7_75t_SL g1098 ( 
.A(n_905),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_840),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_994),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_890),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_952),
.B(n_12),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_952),
.B(n_16),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_850),
.A2(n_62),
.B(n_19),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_944),
.B(n_18),
.Y(n_1105)
);

BUFx2_ASAP7_75t_L g1106 ( 
.A(n_991),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_999),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_959),
.A2(n_857),
.B(n_910),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_858),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_832),
.B(n_21),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1004),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_923),
.B(n_24),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_843),
.A2(n_24),
.B(n_26),
.C(n_27),
.Y(n_1113)
);

AOI21x1_ASAP7_75t_L g1114 ( 
.A1(n_911),
.A2(n_26),
.B(n_32),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_915),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_847),
.A2(n_852),
.B1(n_845),
.B2(n_929),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_927),
.A2(n_35),
.B(n_39),
.C(n_42),
.Y(n_1117)
);

O2A1O1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_951),
.A2(n_35),
.B(n_42),
.C(n_44),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_952),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_1006),
.B(n_44),
.Y(n_1120)
);

CKINVDCx6p67_ASAP7_75t_R g1121 ( 
.A(n_987),
.Y(n_1121)
);

INVxp67_ASAP7_75t_L g1122 ( 
.A(n_983),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_925),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_1006),
.A2(n_48),
.B(n_51),
.C(n_52),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_881),
.A2(n_48),
.B(n_52),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_965),
.A2(n_55),
.B(n_58),
.Y(n_1126)
);

BUFx3_ASAP7_75t_L g1127 ( 
.A(n_985),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_936),
.B(n_55),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_983),
.B(n_58),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_938),
.A2(n_59),
.B1(n_60),
.B2(n_848),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_909),
.A2(n_60),
.B1(n_874),
.B2(n_957),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_921),
.B(n_888),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_SL g1133 ( 
.A1(n_963),
.A2(n_993),
.B1(n_937),
.B2(n_934),
.Y(n_1133)
);

BUFx12f_ASAP7_75t_L g1134 ( 
.A(n_925),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_849),
.A2(n_883),
.B(n_859),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_982),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_997),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_993),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_984),
.B(n_895),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_936),
.B(n_995),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_906),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1001),
.A2(n_916),
.B1(n_871),
.B2(n_891),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_968),
.B(n_953),
.Y(n_1143)
);

OAI21xp33_ASAP7_75t_L g1144 ( 
.A1(n_976),
.A2(n_995),
.B(n_947),
.Y(n_1144)
);

BUFx4f_ASAP7_75t_SL g1145 ( 
.A(n_969),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_864),
.A2(n_866),
.B(n_943),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_887),
.A2(n_962),
.B(n_960),
.C(n_1011),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_846),
.B(n_953),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_977),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_955),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_885),
.A2(n_856),
.B(n_1000),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1002),
.A2(n_1003),
.B(n_1005),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1008),
.B(n_978),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_926),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_933),
.B(n_939),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_R g1156 ( 
.A(n_942),
.B(n_946),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_930),
.Y(n_1157)
);

INVx6_ASAP7_75t_L g1158 ( 
.A(n_1010),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_974),
.Y(n_1159)
);

NAND2x1p5_ASAP7_75t_L g1160 ( 
.A(n_967),
.B(n_940),
.Y(n_1160)
);

AO32x1_ASAP7_75t_L g1161 ( 
.A1(n_945),
.A2(n_897),
.A3(n_988),
.B1(n_935),
.B2(n_1007),
.Y(n_1161)
);

OR2x4_ASAP7_75t_L g1162 ( 
.A(n_941),
.B(n_975),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_979),
.A2(n_990),
.B(n_971),
.C(n_970),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_966),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_964),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_948),
.A2(n_958),
.B(n_954),
.C(n_922),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_924),
.B(n_931),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_1122),
.B(n_928),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1041),
.A2(n_886),
.B(n_902),
.C(n_907),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_1131),
.A2(n_908),
.B(n_914),
.C(n_919),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1015),
.A2(n_1025),
.B(n_1151),
.Y(n_1171)
);

BUFx2_ASAP7_75t_L g1172 ( 
.A(n_1014),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1139),
.A2(n_1108),
.B(n_1132),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_1053),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1075),
.A2(n_1093),
.B1(n_1158),
.B2(n_1141),
.Y(n_1175)
);

OR2x2_ASAP7_75t_L g1176 ( 
.A(n_1098),
.B(n_1138),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1131),
.A2(n_1050),
.B(n_1144),
.C(n_1090),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1163),
.A2(n_1146),
.B(n_1167),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1139),
.A2(n_1132),
.B(n_1019),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1013),
.Y(n_1180)
);

NAND3xp33_ASAP7_75t_L g1181 ( 
.A(n_1120),
.B(n_1105),
.C(n_1096),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1026),
.Y(n_1182)
);

CKINVDCx11_ASAP7_75t_R g1183 ( 
.A(n_1080),
.Y(n_1183)
);

AO21x1_ASAP7_75t_L g1184 ( 
.A1(n_1110),
.A2(n_1142),
.B(n_1130),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1116),
.A2(n_1152),
.B(n_1035),
.Y(n_1185)
);

A2O1A1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1140),
.A2(n_1129),
.B(n_1110),
.C(n_1147),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_1046),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1049),
.A2(n_1043),
.B(n_1092),
.C(n_1089),
.Y(n_1188)
);

AOI221xp5_ASAP7_75t_L g1189 ( 
.A1(n_1133),
.A2(n_1042),
.B1(n_1130),
.B2(n_1034),
.C(n_1067),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1167),
.A2(n_1038),
.B(n_1135),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1154),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1029),
.Y(n_1192)
);

BUFx10_ASAP7_75t_L g1193 ( 
.A(n_1079),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1142),
.A2(n_1116),
.B(n_1017),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1017),
.A2(n_1023),
.B(n_1028),
.Y(n_1195)
);

INVx1_ASAP7_75t_SL g1196 ( 
.A(n_1060),
.Y(n_1196)
);

AO31x2_ASAP7_75t_L g1197 ( 
.A1(n_1166),
.A2(n_1157),
.A3(n_1113),
.B(n_1109),
.Y(n_1197)
);

O2A1O1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1128),
.A2(n_1124),
.B(n_1047),
.C(n_1094),
.Y(n_1198)
);

OR2x6_ASAP7_75t_L g1199 ( 
.A(n_1134),
.B(n_1102),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_1053),
.Y(n_1200)
);

INVx6_ASAP7_75t_L g1201 ( 
.A(n_1100),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1037),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1057),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_1123),
.Y(n_1204)
);

INVxp67_ASAP7_75t_L g1205 ( 
.A(n_1064),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1071),
.B(n_1149),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1016),
.A2(n_1153),
.B(n_1039),
.Y(n_1207)
);

AO31x2_ASAP7_75t_L g1208 ( 
.A1(n_1036),
.A2(n_1059),
.A3(n_1032),
.B(n_1062),
.Y(n_1208)
);

AO21x1_ASAP7_75t_L g1209 ( 
.A1(n_1160),
.A2(n_1084),
.B(n_1104),
.Y(n_1209)
);

CKINVDCx11_ASAP7_75t_R g1210 ( 
.A(n_1121),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1091),
.B(n_1136),
.Y(n_1211)
);

AND2x4_ASAP7_75t_L g1212 ( 
.A(n_1119),
.B(n_1072),
.Y(n_1212)
);

NOR2x1_ASAP7_75t_R g1213 ( 
.A(n_1021),
.B(n_1052),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1158),
.A2(n_1160),
.B1(n_1145),
.B2(n_1127),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1106),
.B(n_1068),
.Y(n_1215)
);

CKINVDCx16_ASAP7_75t_R g1216 ( 
.A(n_1022),
.Y(n_1216)
);

O2A1O1Ixp5_ASAP7_75t_L g1217 ( 
.A1(n_1070),
.A2(n_1031),
.B(n_1045),
.C(n_1112),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_1082),
.Y(n_1218)
);

AO31x2_ASAP7_75t_L g1219 ( 
.A1(n_1032),
.A2(n_1084),
.A3(n_1148),
.B(n_1125),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1091),
.B(n_1137),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1153),
.A2(n_1161),
.B(n_1143),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1055),
.B(n_1073),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1069),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1033),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1048),
.A2(n_1117),
.B(n_1118),
.C(n_1126),
.Y(n_1225)
);

INVx4_ASAP7_75t_L g1226 ( 
.A(n_1123),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1161),
.A2(n_1143),
.B(n_1020),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1044),
.A2(n_1083),
.B(n_1024),
.C(n_1087),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1097),
.A2(n_1101),
.B1(n_1056),
.B2(n_1018),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1161),
.A2(n_1027),
.B(n_1162),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1095),
.Y(n_1231)
);

OAI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1033),
.A2(n_1159),
.B(n_1024),
.Y(n_1232)
);

AO31x2_ASAP7_75t_L g1233 ( 
.A1(n_1164),
.A2(n_1065),
.A3(n_1078),
.B(n_1077),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1165),
.A2(n_1159),
.B(n_1114),
.Y(n_1234)
);

OR2x6_ASAP7_75t_L g1235 ( 
.A(n_1102),
.B(n_1103),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1030),
.B(n_1066),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1076),
.A2(n_1099),
.B(n_1115),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1111),
.B(n_1107),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1067),
.B(n_1083),
.Y(n_1239)
);

AOI221xp5_ASAP7_75t_L g1240 ( 
.A1(n_1058),
.A2(n_1074),
.B1(n_1103),
.B2(n_1051),
.C(n_1086),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_1081),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1119),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_1119),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1076),
.B(n_1099),
.Y(n_1244)
);

AO31x2_ASAP7_75t_L g1245 ( 
.A1(n_1054),
.A2(n_1088),
.A3(n_1061),
.B(n_1156),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1123),
.A2(n_1115),
.B1(n_1053),
.B2(n_1085),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1040),
.B(n_1063),
.Y(n_1247)
);

O2A1O1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1150),
.A2(n_567),
.B(n_535),
.C(n_835),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_1085),
.B(n_1150),
.Y(n_1249)
);

A2O1A1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1150),
.A2(n_1085),
.B(n_835),
.C(n_913),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1041),
.A2(n_835),
.B(n_913),
.C(n_690),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1015),
.A2(n_1025),
.B(n_1151),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_1014),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1075),
.B(n_835),
.Y(n_1254)
);

NOR2xp67_ASAP7_75t_L g1255 ( 
.A(n_1122),
.B(n_686),
.Y(n_1255)
);

OAI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1131),
.A2(n_833),
.B(n_904),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1122),
.B(n_353),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1013),
.Y(n_1258)
);

AOI221x1_ASAP7_75t_L g1259 ( 
.A1(n_1131),
.A2(n_1109),
.B1(n_1130),
.B2(n_1113),
.C(n_956),
.Y(n_1259)
);

AO21x2_ASAP7_75t_L g1260 ( 
.A1(n_1108),
.A2(n_869),
.B(n_1139),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1139),
.A2(n_861),
.B(n_867),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1131),
.A2(n_833),
.B(n_904),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1015),
.A2(n_1025),
.B(n_1151),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1075),
.B(n_835),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1139),
.A2(n_861),
.B(n_867),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1015),
.A2(n_1025),
.B(n_1151),
.Y(n_1266)
);

BUFx4f_ASAP7_75t_L g1267 ( 
.A(n_1014),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1139),
.A2(n_861),
.B(n_867),
.Y(n_1268)
);

OAI22x1_ASAP7_75t_L g1269 ( 
.A1(n_1041),
.A2(n_835),
.B1(n_657),
.B2(n_1092),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1131),
.A2(n_833),
.B(n_904),
.Y(n_1270)
);

BUFx8_ASAP7_75t_L g1271 ( 
.A(n_1106),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1041),
.A2(n_835),
.B1(n_913),
.B2(n_761),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1013),
.Y(n_1273)
);

OR2x2_ASAP7_75t_L g1274 ( 
.A(n_1098),
.B(n_899),
.Y(n_1274)
);

INVx1_ASAP7_75t_SL g1275 ( 
.A(n_1014),
.Y(n_1275)
);

AO31x2_ASAP7_75t_L g1276 ( 
.A1(n_1131),
.A2(n_869),
.A3(n_1142),
.B(n_1116),
.Y(n_1276)
);

OR2x2_ASAP7_75t_L g1277 ( 
.A(n_1098),
.B(n_899),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1139),
.A2(n_861),
.B(n_867),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1075),
.B(n_835),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1122),
.B(n_353),
.Y(n_1280)
);

AOI31xp67_ASAP7_75t_L g1281 ( 
.A1(n_1039),
.A2(n_1139),
.A3(n_1041),
.B(n_1155),
.Y(n_1281)
);

BUFx2_ASAP7_75t_SL g1282 ( 
.A(n_1021),
.Y(n_1282)
);

AO32x2_ASAP7_75t_L g1283 ( 
.A1(n_1131),
.A2(n_1116),
.A3(n_1130),
.B1(n_1133),
.B2(n_1084),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_SL g1284 ( 
.A1(n_1110),
.A2(n_1114),
.B(n_1104),
.Y(n_1284)
);

BUFx4_ASAP7_75t_SL g1285 ( 
.A(n_1021),
.Y(n_1285)
);

OAI22x1_ASAP7_75t_L g1286 ( 
.A1(n_1041),
.A2(n_835),
.B1(n_657),
.B2(n_1092),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1013),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1075),
.B(n_835),
.Y(n_1288)
);

NOR2xp67_ASAP7_75t_SL g1289 ( 
.A(n_1080),
.B(n_618),
.Y(n_1289)
);

AO31x2_ASAP7_75t_L g1290 ( 
.A1(n_1131),
.A2(n_869),
.A3(n_1142),
.B(n_1116),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1131),
.A2(n_833),
.B(n_904),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1139),
.A2(n_861),
.B(n_867),
.Y(n_1292)
);

INVx2_ASAP7_75t_SL g1293 ( 
.A(n_1014),
.Y(n_1293)
);

AO21x2_ASAP7_75t_L g1294 ( 
.A1(n_1108),
.A2(n_869),
.B(n_1139),
.Y(n_1294)
);

AO32x2_ASAP7_75t_L g1295 ( 
.A1(n_1131),
.A2(n_1116),
.A3(n_1130),
.B1(n_1133),
.B2(n_1084),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_SL g1296 ( 
.A1(n_1131),
.A2(n_904),
.B(n_857),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1013),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1122),
.B(n_353),
.Y(n_1298)
);

AO22x1_ASAP7_75t_L g1299 ( 
.A1(n_1050),
.A2(n_835),
.B1(n_501),
.B2(n_567),
.Y(n_1299)
);

AO31x2_ASAP7_75t_L g1300 ( 
.A1(n_1131),
.A2(n_869),
.A3(n_1142),
.B(n_1116),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1075),
.B(n_835),
.Y(n_1301)
);

INVxp67_ASAP7_75t_L g1302 ( 
.A(n_1064),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1131),
.A2(n_833),
.B(n_904),
.Y(n_1303)
);

AO31x2_ASAP7_75t_L g1304 ( 
.A1(n_1131),
.A2(n_869),
.A3(n_1142),
.B(n_1116),
.Y(n_1304)
);

O2A1O1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1050),
.A2(n_567),
.B(n_535),
.C(n_835),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1154),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1041),
.A2(n_835),
.B1(n_913),
.B2(n_761),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1139),
.A2(n_861),
.B(n_867),
.Y(n_1308)
);

AO32x2_ASAP7_75t_L g1309 ( 
.A1(n_1131),
.A2(n_1116),
.A3(n_1130),
.B1(n_1133),
.B2(n_1084),
.Y(n_1309)
);

OR2x2_ASAP7_75t_L g1310 ( 
.A(n_1098),
.B(n_899),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1139),
.A2(n_861),
.B(n_867),
.Y(n_1311)
);

AOI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1050),
.A2(n_898),
.B1(n_667),
.B2(n_835),
.Y(n_1312)
);

AO32x2_ASAP7_75t_L g1313 ( 
.A1(n_1131),
.A2(n_1116),
.A3(n_1130),
.B1(n_1133),
.B2(n_1084),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1139),
.A2(n_861),
.B(n_867),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1075),
.B(n_835),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1013),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1122),
.B(n_667),
.Y(n_1317)
);

O2A1O1Ixp5_ASAP7_75t_SL g1318 ( 
.A1(n_1131),
.A2(n_1094),
.B(n_1130),
.C(n_1120),
.Y(n_1318)
);

O2A1O1Ixp33_ASAP7_75t_L g1319 ( 
.A1(n_1050),
.A2(n_567),
.B(n_535),
.C(n_835),
.Y(n_1319)
);

AO31x2_ASAP7_75t_L g1320 ( 
.A1(n_1131),
.A2(n_869),
.A3(n_1142),
.B(n_1116),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1154),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1015),
.A2(n_1025),
.B(n_1151),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1013),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_SL g1324 ( 
.A1(n_1272),
.A2(n_1307),
.B1(n_1222),
.B2(n_1181),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1192),
.Y(n_1325)
);

INVx3_ASAP7_75t_SL g1326 ( 
.A(n_1201),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_SL g1327 ( 
.A1(n_1256),
.A2(n_1291),
.B1(n_1270),
.B2(n_1262),
.Y(n_1327)
);

INVx1_ASAP7_75t_SL g1328 ( 
.A(n_1196),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1312),
.A2(n_1189),
.B1(n_1269),
.B2(n_1286),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1303),
.A2(n_1299),
.B1(n_1214),
.B2(n_1239),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1305),
.A2(n_1319),
.B1(n_1177),
.B2(n_1251),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_SL g1332 ( 
.A1(n_1254),
.A2(n_1264),
.B1(n_1315),
.B2(n_1279),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1184),
.A2(n_1209),
.B1(n_1288),
.B2(n_1301),
.Y(n_1333)
);

INVx6_ASAP7_75t_L g1334 ( 
.A(n_1201),
.Y(n_1334)
);

CKINVDCx6p67_ASAP7_75t_R g1335 ( 
.A(n_1253),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_SL g1336 ( 
.A1(n_1257),
.A2(n_1298),
.B1(n_1280),
.B2(n_1175),
.Y(n_1336)
);

INVx6_ASAP7_75t_L g1337 ( 
.A(n_1226),
.Y(n_1337)
);

BUFx12f_ASAP7_75t_L g1338 ( 
.A(n_1183),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_SL g1339 ( 
.A1(n_1240),
.A2(n_1259),
.B(n_1248),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1180),
.Y(n_1340)
);

BUFx4f_ASAP7_75t_SL g1341 ( 
.A(n_1193),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1182),
.Y(n_1342)
);

CKINVDCx11_ASAP7_75t_R g1343 ( 
.A(n_1193),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1194),
.A2(n_1317),
.B1(n_1211),
.B2(n_1220),
.Y(n_1344)
);

INVx2_ASAP7_75t_SL g1345 ( 
.A(n_1267),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1203),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1206),
.B(n_1274),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1185),
.A2(n_1277),
.B1(n_1310),
.B2(n_1224),
.Y(n_1348)
);

CKINVDCx20_ASAP7_75t_R g1349 ( 
.A(n_1210),
.Y(n_1349)
);

CKINVDCx11_ASAP7_75t_R g1350 ( 
.A(n_1275),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1224),
.A2(n_1321),
.B1(n_1306),
.B2(n_1191),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_SL g1352 ( 
.A1(n_1216),
.A2(n_1241),
.B1(n_1271),
.B2(n_1267),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1176),
.B(n_1186),
.Y(n_1353)
);

BUFx12f_ASAP7_75t_L g1354 ( 
.A(n_1172),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_SL g1355 ( 
.A1(n_1271),
.A2(n_1235),
.B1(n_1313),
.B2(n_1309),
.Y(n_1355)
);

CKINVDCx11_ASAP7_75t_R g1356 ( 
.A(n_1187),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1191),
.A2(n_1321),
.B1(n_1306),
.B2(n_1168),
.Y(n_1357)
);

INVx6_ASAP7_75t_L g1358 ( 
.A(n_1226),
.Y(n_1358)
);

OAI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1235),
.A2(n_1215),
.B1(n_1231),
.B2(n_1316),
.Y(n_1359)
);

INVx2_ASAP7_75t_SL g1360 ( 
.A(n_1293),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1258),
.Y(n_1361)
);

INVx4_ASAP7_75t_L g1362 ( 
.A(n_1174),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1273),
.Y(n_1363)
);

INVx6_ASAP7_75t_L g1364 ( 
.A(n_1174),
.Y(n_1364)
);

OAI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1287),
.A2(n_1323),
.B1(n_1297),
.B2(n_1202),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1223),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1232),
.A2(n_1283),
.B1(n_1295),
.B2(n_1309),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1205),
.Y(n_1368)
);

INVx8_ASAP7_75t_L g1369 ( 
.A(n_1174),
.Y(n_1369)
);

CKINVDCx11_ASAP7_75t_R g1370 ( 
.A(n_1199),
.Y(n_1370)
);

BUFx12f_ASAP7_75t_L g1371 ( 
.A(n_1243),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1283),
.A2(n_1313),
.B1(n_1309),
.B2(n_1295),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1281),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1238),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1236),
.Y(n_1375)
);

INVx6_ASAP7_75t_L g1376 ( 
.A(n_1200),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1296),
.A2(n_1250),
.B1(n_1255),
.B2(n_1302),
.Y(n_1377)
);

BUFx8_ASAP7_75t_SL g1378 ( 
.A(n_1218),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1198),
.B(n_1179),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1229),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_1200),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1283),
.A2(n_1313),
.B1(n_1295),
.B2(n_1284),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_1285),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1244),
.Y(n_1384)
);

NAND2x1p5_ASAP7_75t_L g1385 ( 
.A(n_1237),
.B(n_1204),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1178),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1173),
.A2(n_1207),
.B1(n_1199),
.B2(n_1294),
.Y(n_1387)
);

BUFx4_ASAP7_75t_R g1388 ( 
.A(n_1289),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1260),
.A2(n_1294),
.B1(n_1311),
.B2(n_1308),
.Y(n_1389)
);

NAND2x1p5_ASAP7_75t_L g1390 ( 
.A(n_1249),
.B(n_1212),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1188),
.B(n_1212),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_1242),
.Y(n_1392)
);

INVx4_ASAP7_75t_L g1393 ( 
.A(n_1260),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1246),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_1282),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_1213),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1318),
.B(n_1265),
.Y(n_1397)
);

AOI22x1_ASAP7_75t_SL g1398 ( 
.A1(n_1228),
.A2(n_1247),
.B1(n_1225),
.B2(n_1245),
.Y(n_1398)
);

CKINVDCx20_ASAP7_75t_R g1399 ( 
.A(n_1230),
.Y(n_1399)
);

OAI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1261),
.A2(n_1268),
.B1(n_1292),
.B2(n_1314),
.Y(n_1400)
);

INVx1_ASAP7_75t_SL g1401 ( 
.A(n_1195),
.Y(n_1401)
);

CKINVDCx6p67_ASAP7_75t_R g1402 ( 
.A(n_1245),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1278),
.A2(n_1221),
.B1(n_1227),
.B2(n_1190),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1234),
.Y(n_1404)
);

AOI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1169),
.A2(n_1170),
.B1(n_1171),
.B2(n_1263),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_SL g1406 ( 
.A1(n_1276),
.A2(n_1320),
.B1(n_1304),
.B2(n_1300),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1219),
.B(n_1197),
.Y(n_1407)
);

BUFx2_ASAP7_75t_SL g1408 ( 
.A(n_1217),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1197),
.Y(n_1409)
);

OA22x2_ASAP7_75t_L g1410 ( 
.A1(n_1252),
.A2(n_1322),
.B1(n_1266),
.B2(n_1290),
.Y(n_1410)
);

BUFx2_ASAP7_75t_SL g1411 ( 
.A(n_1219),
.Y(n_1411)
);

CKINVDCx16_ASAP7_75t_R g1412 ( 
.A(n_1219),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1208),
.Y(n_1413)
);

INVx1_ASAP7_75t_SL g1414 ( 
.A(n_1208),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1276),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1276),
.Y(n_1416)
);

BUFx3_ASAP7_75t_L g1417 ( 
.A(n_1233),
.Y(n_1417)
);

BUFx10_ASAP7_75t_L g1418 ( 
.A(n_1233),
.Y(n_1418)
);

OAI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1290),
.A2(n_1300),
.B1(n_1304),
.B2(n_1320),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1300),
.A2(n_835),
.B1(n_1307),
.B2(n_1272),
.Y(n_1420)
);

INVx3_ASAP7_75t_L g1421 ( 
.A(n_1320),
.Y(n_1421)
);

CKINVDCx11_ASAP7_75t_R g1422 ( 
.A(n_1193),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1272),
.A2(n_835),
.B1(n_1307),
.B2(n_1312),
.Y(n_1423)
);

BUFx12f_ASAP7_75t_L g1424 ( 
.A(n_1183),
.Y(n_1424)
);

BUFx3_ASAP7_75t_L g1425 ( 
.A(n_1267),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1187),
.Y(n_1426)
);

AOI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1312),
.A2(n_898),
.B1(n_501),
.B2(n_1299),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1267),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1272),
.A2(n_835),
.B1(n_1307),
.B2(n_1312),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1312),
.A2(n_1305),
.B1(n_1319),
.B2(n_1307),
.Y(n_1430)
);

CKINVDCx20_ASAP7_75t_R g1431 ( 
.A(n_1183),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1192),
.Y(n_1432)
);

BUFx3_ASAP7_75t_L g1433 ( 
.A(n_1267),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_1267),
.Y(n_1434)
);

INVx6_ASAP7_75t_L g1435 ( 
.A(n_1201),
.Y(n_1435)
);

INVx1_ASAP7_75t_SL g1436 ( 
.A(n_1196),
.Y(n_1436)
);

BUFx4_ASAP7_75t_R g1437 ( 
.A(n_1193),
.Y(n_1437)
);

INVxp67_ASAP7_75t_L g1438 ( 
.A(n_1187),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_SL g1439 ( 
.A1(n_1272),
.A2(n_500),
.B1(n_1307),
.B2(n_623),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_SL g1440 ( 
.A1(n_1272),
.A2(n_500),
.B1(n_1307),
.B2(n_623),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1272),
.A2(n_835),
.B1(n_1307),
.B2(n_1312),
.Y(n_1441)
);

INVx6_ASAP7_75t_L g1442 ( 
.A(n_1201),
.Y(n_1442)
);

INVx6_ASAP7_75t_L g1443 ( 
.A(n_1201),
.Y(n_1443)
);

INVx2_ASAP7_75t_SL g1444 ( 
.A(n_1267),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_SL g1445 ( 
.A1(n_1272),
.A2(n_500),
.B1(n_1307),
.B2(n_623),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_SL g1446 ( 
.A1(n_1272),
.A2(n_500),
.B1(n_1307),
.B2(n_623),
.Y(n_1446)
);

OAI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1312),
.A2(n_1131),
.B1(n_1307),
.B2(n_1272),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1192),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1272),
.A2(n_835),
.B1(n_1307),
.B2(n_1312),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1272),
.A2(n_835),
.B1(n_1307),
.B2(n_1312),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_SL g1451 ( 
.A1(n_1344),
.A2(n_1391),
.B(n_1377),
.Y(n_1451)
);

INVx1_ASAP7_75t_SL g1452 ( 
.A(n_1328),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1332),
.B(n_1347),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1407),
.B(n_1404),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1409),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_1334),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1412),
.B(n_1415),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1432),
.Y(n_1458)
);

INVx2_ASAP7_75t_SL g1459 ( 
.A(n_1448),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1325),
.Y(n_1460)
);

AO31x2_ASAP7_75t_L g1461 ( 
.A1(n_1331),
.A2(n_1373),
.A3(n_1393),
.B(n_1430),
.Y(n_1461)
);

INVx6_ASAP7_75t_L g1462 ( 
.A(n_1334),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1366),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1367),
.B(n_1382),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1327),
.A2(n_1446),
.B1(n_1439),
.B2(n_1445),
.Y(n_1465)
);

INVx2_ASAP7_75t_SL g1466 ( 
.A(n_1366),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_SL g1467 ( 
.A(n_1383),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1344),
.B(n_1348),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1400),
.A2(n_1379),
.B(n_1401),
.Y(n_1469)
);

CKINVDCx11_ASAP7_75t_R g1470 ( 
.A(n_1349),
.Y(n_1470)
);

INVx3_ASAP7_75t_L g1471 ( 
.A(n_1404),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1413),
.Y(n_1472)
);

AO21x2_ASAP7_75t_L g1473 ( 
.A1(n_1400),
.A2(n_1405),
.B(n_1397),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1414),
.B(n_1416),
.Y(n_1474)
);

INVxp67_ASAP7_75t_L g1475 ( 
.A(n_1368),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1348),
.B(n_1353),
.Y(n_1476)
);

BUFx2_ASAP7_75t_L g1477 ( 
.A(n_1399),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1440),
.A2(n_1429),
.B(n_1450),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1342),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1342),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1367),
.B(n_1382),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1421),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1421),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1411),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1417),
.B(n_1387),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1372),
.B(n_1355),
.Y(n_1486)
);

AOI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1410),
.A2(n_1386),
.B(n_1373),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1410),
.A2(n_1389),
.B(n_1386),
.Y(n_1488)
);

INVx2_ASAP7_75t_SL g1489 ( 
.A(n_1337),
.Y(n_1489)
);

BUFx3_ASAP7_75t_L g1490 ( 
.A(n_1334),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1372),
.B(n_1420),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1363),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1420),
.B(n_1329),
.Y(n_1493)
);

INVxp67_ASAP7_75t_SL g1494 ( 
.A(n_1365),
.Y(n_1494)
);

CKINVDCx6p67_ASAP7_75t_R g1495 ( 
.A(n_1326),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1340),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1329),
.B(n_1406),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1351),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1426),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1351),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1419),
.Y(n_1501)
);

AOI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1380),
.A2(n_1394),
.B(n_1346),
.Y(n_1502)
);

AOI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1361),
.A2(n_1384),
.B(n_1374),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1419),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1375),
.B(n_1336),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1418),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1333),
.B(n_1324),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1392),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1385),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1365),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1408),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1402),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1398),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1357),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1333),
.B(n_1357),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1387),
.Y(n_1516)
);

NAND4xp25_ASAP7_75t_L g1517 ( 
.A(n_1427),
.B(n_1423),
.C(n_1450),
.D(n_1449),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_1435),
.Y(n_1518)
);

OR2x6_ASAP7_75t_L g1519 ( 
.A(n_1339),
.B(n_1390),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1389),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1403),
.A2(n_1390),
.B(n_1441),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1438),
.Y(n_1522)
);

AO21x2_ASAP7_75t_L g1523 ( 
.A1(n_1447),
.A2(n_1359),
.B(n_1403),
.Y(n_1523)
);

AOI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1330),
.A2(n_1447),
.B(n_1449),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1423),
.B(n_1441),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1381),
.Y(n_1526)
);

BUFx4f_ASAP7_75t_SL g1527 ( 
.A(n_1338),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_L g1528 ( 
.A1(n_1429),
.A2(n_1359),
.B(n_1388),
.Y(n_1528)
);

BUFx4f_ASAP7_75t_SL g1529 ( 
.A(n_1424),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1436),
.Y(n_1530)
);

NOR2xp67_ASAP7_75t_L g1531 ( 
.A(n_1362),
.B(n_1444),
.Y(n_1531)
);

AO21x2_ASAP7_75t_L g1532 ( 
.A1(n_1469),
.A2(n_1388),
.B(n_1437),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1457),
.B(n_1472),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1517),
.A2(n_1370),
.B1(n_1356),
.B2(n_1350),
.Y(n_1534)
);

INVxp67_ASAP7_75t_L g1535 ( 
.A(n_1463),
.Y(n_1535)
);

O2A1O1Ixp33_ASAP7_75t_L g1536 ( 
.A1(n_1478),
.A2(n_1360),
.B(n_1345),
.C(n_1326),
.Y(n_1536)
);

OAI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1524),
.A2(n_1352),
.B(n_1431),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1465),
.A2(n_1395),
.B1(n_1341),
.B2(n_1425),
.Y(n_1538)
);

AOI21xp33_ASAP7_75t_L g1539 ( 
.A1(n_1451),
.A2(n_1354),
.B(n_1434),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1453),
.B(n_1428),
.Y(n_1540)
);

AOI221xp5_ASAP7_75t_L g1541 ( 
.A1(n_1507),
.A2(n_1434),
.B1(n_1433),
.B2(n_1428),
.C(n_1425),
.Y(n_1541)
);

NAND2xp33_ASAP7_75t_SL g1542 ( 
.A(n_1513),
.B(n_1507),
.Y(n_1542)
);

O2A1O1Ixp33_ASAP7_75t_L g1543 ( 
.A1(n_1451),
.A2(n_1341),
.B(n_1422),
.C(n_1343),
.Y(n_1543)
);

O2A1O1Ixp33_ASAP7_75t_SL g1544 ( 
.A1(n_1513),
.A2(n_1468),
.B(n_1476),
.C(n_1505),
.Y(n_1544)
);

CKINVDCx6p67_ASAP7_75t_R g1545 ( 
.A(n_1470),
.Y(n_1545)
);

AOI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1525),
.A2(n_1335),
.B1(n_1371),
.B2(n_1443),
.Y(n_1546)
);

OAI211xp5_ASAP7_75t_L g1547 ( 
.A1(n_1524),
.A2(n_1396),
.B(n_1362),
.C(n_1369),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1457),
.B(n_1369),
.Y(n_1548)
);

A2O1A1Ixp33_ASAP7_75t_L g1549 ( 
.A1(n_1528),
.A2(n_1369),
.B(n_1337),
.C(n_1358),
.Y(n_1549)
);

AO21x1_ASAP7_75t_L g1550 ( 
.A1(n_1497),
.A2(n_1364),
.B(n_1376),
.Y(n_1550)
);

OAI21x1_ASAP7_75t_L g1551 ( 
.A1(n_1487),
.A2(n_1488),
.B(n_1502),
.Y(n_1551)
);

OAI21x1_ASAP7_75t_SL g1552 ( 
.A1(n_1503),
.A2(n_1358),
.B(n_1378),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1460),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1493),
.B(n_1435),
.Y(n_1554)
);

OA21x2_ASAP7_75t_L g1555 ( 
.A1(n_1488),
.A2(n_1376),
.B(n_1435),
.Y(n_1555)
);

OAI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1477),
.A2(n_1442),
.B1(n_1443),
.B2(n_1519),
.Y(n_1556)
);

OA21x2_ASAP7_75t_L g1557 ( 
.A1(n_1521),
.A2(n_1520),
.B(n_1504),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1473),
.A2(n_1442),
.B(n_1443),
.Y(n_1558)
);

A2O1A1Ixp33_ASAP7_75t_L g1559 ( 
.A1(n_1528),
.A2(n_1442),
.B(n_1493),
.C(n_1497),
.Y(n_1559)
);

OA21x2_ASAP7_75t_L g1560 ( 
.A1(n_1521),
.A2(n_1520),
.B(n_1504),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1499),
.B(n_1508),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1519),
.A2(n_1495),
.B1(n_1475),
.B2(n_1494),
.Y(n_1562)
);

O2A1O1Ixp33_ASAP7_75t_L g1563 ( 
.A1(n_1522),
.A2(n_1519),
.B(n_1530),
.C(n_1511),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1495),
.A2(n_1452),
.B1(n_1462),
.B2(n_1515),
.Y(n_1564)
);

OA21x2_ASAP7_75t_L g1565 ( 
.A1(n_1501),
.A2(n_1516),
.B(n_1484),
.Y(n_1565)
);

AOI211xp5_ASAP7_75t_L g1566 ( 
.A1(n_1514),
.A2(n_1512),
.B(n_1510),
.C(n_1474),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1496),
.B(n_1458),
.Y(n_1567)
);

AOI221xp5_ASAP7_75t_L g1568 ( 
.A1(n_1514),
.A2(n_1491),
.B1(n_1498),
.B2(n_1500),
.C(n_1501),
.Y(n_1568)
);

NOR2x1_ASAP7_75t_SL g1569 ( 
.A(n_1523),
.B(n_1506),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1454),
.B(n_1471),
.Y(n_1570)
);

AO32x2_ASAP7_75t_L g1571 ( 
.A1(n_1459),
.A2(n_1466),
.A3(n_1489),
.B1(n_1481),
.B2(n_1464),
.Y(n_1571)
);

NAND3xp33_ASAP7_75t_L g1572 ( 
.A(n_1498),
.B(n_1500),
.C(n_1484),
.Y(n_1572)
);

A2O1A1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1485),
.A2(n_1491),
.B(n_1486),
.C(n_1523),
.Y(n_1573)
);

NOR2x1_ASAP7_75t_SL g1574 ( 
.A(n_1523),
.B(n_1506),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1486),
.B(n_1526),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1526),
.B(n_1481),
.Y(n_1576)
);

A2O1A1Ixp33_ASAP7_75t_L g1577 ( 
.A1(n_1485),
.A2(n_1464),
.B(n_1459),
.C(n_1531),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1571),
.B(n_1557),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1553),
.Y(n_1579)
);

OAI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1573),
.A2(n_1485),
.B1(n_1462),
.B2(n_1518),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1571),
.B(n_1473),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1571),
.B(n_1485),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1565),
.B(n_1557),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1571),
.B(n_1482),
.Y(n_1584)
);

CKINVDCx20_ASAP7_75t_R g1585 ( 
.A(n_1545),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1565),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1560),
.B(n_1483),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1560),
.B(n_1455),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_1552),
.Y(n_1589)
);

INVx4_ASAP7_75t_L g1590 ( 
.A(n_1532),
.Y(n_1590)
);

BUFx2_ASAP7_75t_L g1591 ( 
.A(n_1555),
.Y(n_1591)
);

NOR2x1_ASAP7_75t_SL g1592 ( 
.A(n_1532),
.B(n_1509),
.Y(n_1592)
);

INVxp67_ASAP7_75t_SL g1593 ( 
.A(n_1572),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_L g1594 ( 
.A(n_1544),
.B(n_1456),
.Y(n_1594)
);

BUFx3_ASAP7_75t_L g1595 ( 
.A(n_1555),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1570),
.B(n_1471),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1567),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1533),
.B(n_1535),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1535),
.Y(n_1599)
);

OAI221xp5_ASAP7_75t_SL g1600 ( 
.A1(n_1534),
.A2(n_1490),
.B1(n_1489),
.B2(n_1479),
.C(n_1480),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1538),
.A2(n_1529),
.B1(n_1527),
.B2(n_1492),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1573),
.B(n_1461),
.Y(n_1602)
);

OR2x2_ASAP7_75t_SL g1603 ( 
.A(n_1555),
.B(n_1548),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1576),
.B(n_1455),
.Y(n_1604)
);

INVx5_ASAP7_75t_SL g1605 ( 
.A(n_1596),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1593),
.B(n_1597),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1582),
.B(n_1578),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1579),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1588),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1579),
.Y(n_1610)
);

NOR3xp33_ASAP7_75t_SL g1611 ( 
.A(n_1594),
.B(n_1547),
.C(n_1537),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1582),
.B(n_1569),
.Y(n_1612)
);

INVx4_ASAP7_75t_L g1613 ( 
.A(n_1589),
.Y(n_1613)
);

NAND2xp33_ASAP7_75t_R g1614 ( 
.A(n_1594),
.B(n_1540),
.Y(n_1614)
);

AOI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1593),
.A2(n_1542),
.B(n_1544),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1582),
.B(n_1574),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1578),
.B(n_1551),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1586),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1597),
.B(n_1568),
.Y(n_1619)
);

AOI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1580),
.A2(n_1542),
.B1(n_1540),
.B2(n_1541),
.Y(n_1620)
);

NOR2xp33_ASAP7_75t_L g1621 ( 
.A(n_1598),
.B(n_1554),
.Y(n_1621)
);

OAI31xp33_ASAP7_75t_L g1622 ( 
.A1(n_1580),
.A2(n_1559),
.A3(n_1536),
.B(n_1534),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_SL g1623 ( 
.A1(n_1592),
.A2(n_1543),
.B(n_1563),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1602),
.A2(n_1566),
.B1(n_1559),
.B2(n_1577),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1578),
.B(n_1561),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1581),
.B(n_1584),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1583),
.B(n_1575),
.Y(n_1627)
);

INVx2_ASAP7_75t_SL g1628 ( 
.A(n_1595),
.Y(n_1628)
);

INVxp67_ASAP7_75t_L g1629 ( 
.A(n_1586),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1584),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1584),
.Y(n_1631)
);

BUFx2_ASAP7_75t_L g1632 ( 
.A(n_1603),
.Y(n_1632)
);

NAND2x1_ASAP7_75t_L g1633 ( 
.A(n_1632),
.B(n_1623),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1607),
.B(n_1591),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1606),
.B(n_1599),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1618),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1618),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1627),
.B(n_1602),
.Y(n_1638)
);

AOI21xp33_ASAP7_75t_SL g1639 ( 
.A1(n_1622),
.A2(n_1539),
.B(n_1546),
.Y(n_1639)
);

INVx1_ASAP7_75t_SL g1640 ( 
.A(n_1606),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1609),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1608),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1626),
.B(n_1630),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1629),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1627),
.B(n_1602),
.Y(n_1645)
);

INVx2_ASAP7_75t_SL g1646 ( 
.A(n_1628),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_R g1647 ( 
.A(n_1614),
.B(n_1585),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1628),
.B(n_1595),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1630),
.B(n_1583),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1626),
.B(n_1595),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1626),
.B(n_1590),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1631),
.B(n_1590),
.Y(n_1652)
);

BUFx2_ASAP7_75t_L g1653 ( 
.A(n_1613),
.Y(n_1653)
);

AOI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1622),
.A2(n_1590),
.B1(n_1556),
.B2(n_1562),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1628),
.B(n_1587),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1608),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1627),
.B(n_1625),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1631),
.B(n_1590),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1610),
.Y(n_1659)
);

OAI221xp5_ASAP7_75t_L g1660 ( 
.A1(n_1615),
.A2(n_1590),
.B1(n_1601),
.B2(n_1600),
.C(n_1549),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1632),
.B(n_1587),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1619),
.B(n_1599),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1612),
.B(n_1604),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1662),
.B(n_1619),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1637),
.Y(n_1665)
);

NAND2xp33_ASAP7_75t_R g1666 ( 
.A(n_1647),
.B(n_1611),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1637),
.Y(n_1667)
);

OAI211xp5_ASAP7_75t_SL g1668 ( 
.A1(n_1654),
.A2(n_1611),
.B(n_1615),
.C(n_1620),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1644),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1649),
.Y(n_1670)
);

INVx1_ASAP7_75t_SL g1671 ( 
.A(n_1633),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1644),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1636),
.Y(n_1673)
);

INVx2_ASAP7_75t_SL g1674 ( 
.A(n_1646),
.Y(n_1674)
);

NOR2xp67_ASAP7_75t_L g1675 ( 
.A(n_1646),
.B(n_1613),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1636),
.Y(n_1676)
);

INVxp67_ASAP7_75t_L g1677 ( 
.A(n_1662),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1663),
.B(n_1605),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1640),
.B(n_1621),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1640),
.B(n_1625),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1663),
.B(n_1605),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1642),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1635),
.Y(n_1683)
);

INVx2_ASAP7_75t_SL g1684 ( 
.A(n_1646),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1663),
.B(n_1605),
.Y(n_1685)
);

AND2x4_ASAP7_75t_L g1686 ( 
.A(n_1653),
.B(n_1613),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1643),
.B(n_1605),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1635),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1642),
.Y(n_1689)
);

AOI21xp33_ASAP7_75t_L g1690 ( 
.A1(n_1633),
.A2(n_1624),
.B(n_1620),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1643),
.B(n_1605),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1638),
.B(n_1625),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1656),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1649),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1656),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1653),
.B(n_1613),
.Y(n_1696)
);

HB1xp67_ASAP7_75t_L g1697 ( 
.A(n_1643),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1649),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1639),
.B(n_1621),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1638),
.B(n_1645),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1659),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1650),
.B(n_1605),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1660),
.A2(n_1624),
.B1(n_1550),
.B2(n_1613),
.Y(n_1703)
);

NOR2x1_ASAP7_75t_SL g1704 ( 
.A(n_1657),
.B(n_1612),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1645),
.B(n_1617),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1659),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1704),
.B(n_1650),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1669),
.B(n_1657),
.Y(n_1708)
);

AO21x2_ASAP7_75t_L g1709 ( 
.A1(n_1690),
.A2(n_1639),
.B(n_1661),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1682),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1674),
.Y(n_1711)
);

INVx1_ASAP7_75t_SL g1712 ( 
.A(n_1671),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_L g1713 ( 
.A(n_1699),
.B(n_1585),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1664),
.B(n_1661),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1682),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1693),
.Y(n_1716)
);

NOR2xp67_ASAP7_75t_L g1717 ( 
.A(n_1703),
.B(n_1660),
.Y(n_1717)
);

HB1xp67_ASAP7_75t_L g1718 ( 
.A(n_1697),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1677),
.B(n_1661),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1693),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1672),
.B(n_1612),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1667),
.B(n_1617),
.Y(n_1722)
);

NOR2x1_ASAP7_75t_SL g1723 ( 
.A(n_1674),
.B(n_1652),
.Y(n_1723)
);

NOR2x1_ASAP7_75t_L g1724 ( 
.A(n_1668),
.B(n_1648),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1684),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1679),
.B(n_1616),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1700),
.B(n_1617),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1683),
.B(n_1616),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1688),
.B(n_1616),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1686),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1704),
.B(n_1650),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1700),
.B(n_1641),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1673),
.B(n_1651),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1665),
.B(n_1641),
.Y(n_1734)
);

INVx2_ASAP7_75t_SL g1735 ( 
.A(n_1684),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1702),
.B(n_1634),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1706),
.Y(n_1737)
);

BUFx2_ASAP7_75t_L g1738 ( 
.A(n_1686),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1673),
.B(n_1651),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1670),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1676),
.B(n_1651),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1702),
.B(n_1634),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1717),
.B(n_1665),
.Y(n_1743)
);

NOR2x1_ASAP7_75t_L g1744 ( 
.A(n_1709),
.B(n_1675),
.Y(n_1744)
);

OAI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1717),
.A2(n_1724),
.B1(n_1712),
.B2(n_1713),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1723),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_SL g1747 ( 
.A(n_1724),
.B(n_1686),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1723),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1718),
.Y(n_1749)
);

OAI32xp33_ASAP7_75t_L g1750 ( 
.A1(n_1712),
.A2(n_1666),
.A3(n_1680),
.B1(n_1692),
.B2(n_1705),
.Y(n_1750)
);

OA21x2_ASAP7_75t_L g1751 ( 
.A1(n_1711),
.A2(n_1676),
.B(n_1670),
.Y(n_1751)
);

INVxp33_ASAP7_75t_L g1752 ( 
.A(n_1708),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1710),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1710),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1709),
.A2(n_1687),
.B1(n_1691),
.B2(n_1696),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1709),
.B(n_1467),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1730),
.B(n_1696),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1730),
.B(n_1696),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1715),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1738),
.B(n_1687),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1715),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1716),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1738),
.B(n_1691),
.Y(n_1763)
);

AOI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1719),
.A2(n_1680),
.B(n_1592),
.Y(n_1764)
);

INVx1_ASAP7_75t_SL g1765 ( 
.A(n_1708),
.Y(n_1765)
);

CKINVDCx20_ASAP7_75t_R g1766 ( 
.A(n_1714),
.Y(n_1766)
);

AOI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1707),
.A2(n_1685),
.B1(n_1678),
.B2(n_1681),
.Y(n_1767)
);

CKINVDCx16_ASAP7_75t_R g1768 ( 
.A(n_1736),
.Y(n_1768)
);

INVxp33_ASAP7_75t_L g1769 ( 
.A(n_1756),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1765),
.B(n_1736),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1753),
.Y(n_1771)
);

INVx3_ASAP7_75t_L g1772 ( 
.A(n_1751),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1754),
.Y(n_1773)
);

OAI211xp5_ASAP7_75t_L g1774 ( 
.A1(n_1747),
.A2(n_1707),
.B(n_1731),
.C(n_1735),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1749),
.B(n_1742),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1768),
.B(n_1742),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1759),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1761),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1743),
.B(n_1711),
.Y(n_1779)
);

INVx1_ASAP7_75t_SL g1780 ( 
.A(n_1747),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1752),
.B(n_1735),
.Y(n_1781)
);

OAI321xp33_ASAP7_75t_L g1782 ( 
.A1(n_1745),
.A2(n_1731),
.A3(n_1740),
.B1(n_1725),
.B2(n_1741),
.C(n_1733),
.Y(n_1782)
);

INVx2_ASAP7_75t_SL g1783 ( 
.A(n_1746),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1752),
.B(n_1725),
.Y(n_1784)
);

AND2x4_ASAP7_75t_SL g1785 ( 
.A(n_1746),
.B(n_1740),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1756),
.A2(n_1721),
.B1(n_1726),
.B2(n_1740),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1762),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1767),
.B(n_1678),
.Y(n_1788)
);

INVx3_ASAP7_75t_L g1789 ( 
.A(n_1772),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1780),
.B(n_1748),
.Y(n_1790)
);

INVx1_ASAP7_75t_SL g1791 ( 
.A(n_1776),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1772),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1784),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1781),
.B(n_1766),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1772),
.Y(n_1795)
);

NOR2x1_ASAP7_75t_L g1796 ( 
.A(n_1774),
.B(n_1744),
.Y(n_1796)
);

NAND2xp33_ASAP7_75t_SL g1797 ( 
.A(n_1769),
.B(n_1755),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1785),
.Y(n_1798)
);

NAND3xp33_ASAP7_75t_SL g1799 ( 
.A(n_1769),
.B(n_1766),
.C(n_1748),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1785),
.Y(n_1800)
);

BUFx6f_ASAP7_75t_L g1801 ( 
.A(n_1789),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1789),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1790),
.B(n_1781),
.Y(n_1803)
);

OAI211xp5_ASAP7_75t_SL g1804 ( 
.A1(n_1794),
.A2(n_1779),
.B(n_1775),
.C(n_1770),
.Y(n_1804)
);

NOR2xp33_ASAP7_75t_L g1805 ( 
.A(n_1791),
.B(n_1799),
.Y(n_1805)
);

AOI21x1_ASAP7_75t_L g1806 ( 
.A1(n_1795),
.A2(n_1783),
.B(n_1751),
.Y(n_1806)
);

OAI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1796),
.A2(n_1786),
.B1(n_1763),
.B2(n_1760),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1789),
.Y(n_1808)
);

NAND3xp33_ASAP7_75t_L g1809 ( 
.A(n_1797),
.B(n_1783),
.C(n_1773),
.Y(n_1809)
);

NOR3xp33_ASAP7_75t_L g1810 ( 
.A(n_1797),
.B(n_1782),
.C(n_1750),
.Y(n_1810)
);

OAI321xp33_ASAP7_75t_L g1811 ( 
.A1(n_1807),
.A2(n_1793),
.A3(n_1798),
.B1(n_1800),
.B2(n_1790),
.C(n_1788),
.Y(n_1811)
);

OAI221xp5_ASAP7_75t_L g1812 ( 
.A1(n_1810),
.A2(n_1788),
.B1(n_1757),
.B2(n_1758),
.C(n_1764),
.Y(n_1812)
);

NOR2x1_ASAP7_75t_L g1813 ( 
.A(n_1809),
.B(n_1792),
.Y(n_1813)
);

OAI21xp5_ASAP7_75t_SL g1814 ( 
.A1(n_1805),
.A2(n_1777),
.B(n_1771),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1803),
.B(n_1792),
.Y(n_1815)
);

AOI221xp5_ASAP7_75t_L g1816 ( 
.A1(n_1811),
.A2(n_1812),
.B1(n_1814),
.B2(n_1804),
.C(n_1815),
.Y(n_1816)
);

AOI221xp5_ASAP7_75t_L g1817 ( 
.A1(n_1813),
.A2(n_1778),
.B1(n_1787),
.B2(n_1808),
.C(n_1801),
.Y(n_1817)
);

NOR3xp33_ASAP7_75t_L g1818 ( 
.A(n_1811),
.B(n_1802),
.C(n_1806),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1813),
.B(n_1801),
.Y(n_1819)
);

AOI221xp5_ASAP7_75t_L g1820 ( 
.A1(n_1811),
.A2(n_1801),
.B1(n_1716),
.B2(n_1737),
.C(n_1720),
.Y(n_1820)
);

NOR2xp67_ASAP7_75t_L g1821 ( 
.A(n_1811),
.B(n_1720),
.Y(n_1821)
);

AND2x4_ASAP7_75t_L g1822 ( 
.A(n_1819),
.B(n_1681),
.Y(n_1822)
);

INVxp67_ASAP7_75t_L g1823 ( 
.A(n_1821),
.Y(n_1823)
);

XNOR2x1_ASAP7_75t_L g1824 ( 
.A(n_1816),
.B(n_1685),
.Y(n_1824)
);

NOR2x1_ASAP7_75t_L g1825 ( 
.A(n_1818),
.B(n_1751),
.Y(n_1825)
);

AO22x2_ASAP7_75t_L g1826 ( 
.A1(n_1817),
.A2(n_1737),
.B1(n_1734),
.B2(n_1694),
.Y(n_1826)
);

A2O1A1Ixp33_ASAP7_75t_SL g1827 ( 
.A1(n_1823),
.A2(n_1820),
.B(n_1698),
.C(n_1694),
.Y(n_1827)
);

AOI22x1_ASAP7_75t_L g1828 ( 
.A1(n_1826),
.A2(n_1734),
.B1(n_1698),
.B2(n_1732),
.Y(n_1828)
);

OAI22xp33_ASAP7_75t_SL g1829 ( 
.A1(n_1825),
.A2(n_1732),
.B1(n_1722),
.B2(n_1739),
.Y(n_1829)
);

AOI22xp33_ASAP7_75t_SL g1830 ( 
.A1(n_1828),
.A2(n_1822),
.B1(n_1824),
.B2(n_1722),
.Y(n_1830)
);

AOI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1830),
.A2(n_1829),
.B1(n_1827),
.B2(n_1729),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1831),
.B(n_1728),
.Y(n_1832)
);

OR3x1_ASAP7_75t_L g1833 ( 
.A(n_1831),
.B(n_1706),
.C(n_1695),
.Y(n_1833)
);

HB1xp67_ASAP7_75t_L g1834 ( 
.A(n_1833),
.Y(n_1834)
);

AOI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1832),
.A2(n_1727),
.B1(n_1648),
.B2(n_1658),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1834),
.B(n_1689),
.Y(n_1836)
);

AOI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1835),
.A2(n_1727),
.B1(n_1648),
.B2(n_1652),
.Y(n_1837)
);

OAI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1836),
.A2(n_1705),
.B(n_1701),
.Y(n_1838)
);

OAI31xp33_ASAP7_75t_L g1839 ( 
.A1(n_1838),
.A2(n_1837),
.A3(n_1658),
.B(n_1652),
.Y(n_1839)
);

XNOR2xp5_ASAP7_75t_L g1840 ( 
.A(n_1839),
.B(n_1531),
.Y(n_1840)
);

AOI221xp5_ASAP7_75t_L g1841 ( 
.A1(n_1840),
.A2(n_1658),
.B1(n_1648),
.B2(n_1629),
.C(n_1655),
.Y(n_1841)
);

AOI211xp5_ASAP7_75t_L g1842 ( 
.A1(n_1841),
.A2(n_1564),
.B(n_1692),
.C(n_1558),
.Y(n_1842)
);


endmodule