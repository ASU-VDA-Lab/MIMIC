module fake_jpeg_6324_n_326 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_34),
.B(n_38),
.Y(n_52)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_40),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_18),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_44),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

NAND2xp33_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_28),
.Y(n_46)
);

OR2x2_ASAP7_75t_SL g85 ( 
.A(n_46),
.B(n_69),
.Y(n_85)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_28),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_51),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_44),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_53),
.Y(n_71)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_58),
.Y(n_78)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_20),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_60),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_38),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_62),
.Y(n_87)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_64),
.Y(n_92)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_36),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_77),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_56),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_84),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_43),
.B1(n_35),
.B2(n_41),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_74),
.A2(n_82),
.B1(n_88),
.B2(n_25),
.Y(n_104)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_45),
.B(n_20),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_80),
.B(n_30),
.Y(n_107)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_89),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_43),
.B1(n_35),
.B2(n_36),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_35),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_34),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_93),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_49),
.A2(n_32),
.B1(n_43),
.B2(n_35),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_34),
.Y(n_93)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_102),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_93),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_83),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_43),
.B1(n_41),
.B2(n_32),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_100),
.A2(n_101),
.B1(n_120),
.B2(n_25),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_L g101 ( 
.A1(n_74),
.A2(n_66),
.B1(n_41),
.B2(n_42),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_104),
.A2(n_118),
.B1(n_79),
.B2(n_87),
.Y(n_136)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_109),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_107),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_80),
.B(n_31),
.Y(n_115)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_19),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_73),
.A2(n_57),
.B1(n_58),
.B2(n_25),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_85),
.A2(n_25),
.B1(n_66),
.B2(n_42),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_92),
.Y(n_121)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_85),
.C(n_73),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_127),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_140),
.Y(n_158)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_118),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_135),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_82),
.C(n_87),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_128),
.A2(n_133),
.B1(n_143),
.B2(n_144),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_96),
.A2(n_83),
.B1(n_71),
.B2(n_79),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_103),
.A2(n_23),
.B(n_19),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_136),
.A2(n_138),
.B1(n_108),
.B2(n_112),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_SL g138 ( 
.A1(n_103),
.A2(n_101),
.B(n_120),
.C(n_100),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_97),
.A2(n_94),
.B(n_26),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_22),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_94),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_106),
.B1(n_104),
.B2(n_114),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_89),
.B1(n_81),
.B2(n_70),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_109),
.A2(n_19),
.B1(n_23),
.B2(n_30),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_147),
.A2(n_30),
.B1(n_23),
.B2(n_31),
.Y(n_176)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_148),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_146),
.B(n_95),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_149),
.B(n_156),
.Y(n_186)
);

INVx3_ASAP7_75t_SL g150 ( 
.A(n_124),
.Y(n_150)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_105),
.Y(n_151)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

OAI22x1_ASAP7_75t_L g154 ( 
.A1(n_138),
.A2(n_76),
.B1(n_22),
.B2(n_67),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_154),
.A2(n_171),
.B1(n_175),
.B2(n_176),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_155),
.A2(n_166),
.B1(n_128),
.B2(n_139),
.Y(n_180)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

OA21x2_ASAP7_75t_L g159 ( 
.A1(n_129),
.A2(n_42),
.B(n_17),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_160),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_144),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_163),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_140),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_162),
.Y(n_183)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_22),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_138),
.A2(n_62),
.B1(n_64),
.B2(n_42),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_98),
.Y(n_167)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_125),
.Y(n_168)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_125),
.Y(n_169)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_142),
.Y(n_170)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_133),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_122),
.B(n_110),
.Y(n_173)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_173),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_142),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_174),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_130),
.B(n_31),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_171),
.A2(n_135),
.B(n_136),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_185),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_157),
.Y(n_213)
);

OAI22x1_ASAP7_75t_SL g181 ( 
.A1(n_154),
.A2(n_138),
.B1(n_127),
.B2(n_145),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_181),
.A2(n_191),
.B1(n_156),
.B2(n_159),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_163),
.A2(n_138),
.B1(n_141),
.B2(n_126),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_182),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_150),
.A2(n_126),
.B(n_141),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_145),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_165),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_166),
.A2(n_130),
.B1(n_119),
.B2(n_132),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_173),
.C(n_172),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_195),
.C(n_202),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_197),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_132),
.C(n_67),
.Y(n_195)
);

CKINVDCx12_ASAP7_75t_R g196 ( 
.A(n_153),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_153),
.B(n_67),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_67),
.C(n_65),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_181),
.A2(n_158),
.B(n_157),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_204),
.B(n_220),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_203),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_206),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_186),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_152),
.Y(n_207)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_191),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_211),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_209),
.A2(n_213),
.B1(n_221),
.B2(n_188),
.Y(n_238)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_225),
.Y(n_243)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_202),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_170),
.Y(n_214)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_214),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_183),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_224),
.Y(n_241)
);

XOR2x1_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_152),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_218),
.B(n_227),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_161),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_170),
.C(n_168),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_228),
.C(n_201),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_198),
.B(n_159),
.Y(n_223)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_179),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_194),
.B(n_29),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_197),
.B(n_22),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_137),
.C(n_98),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_240),
.C(n_217),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_222),
.C(n_227),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_204),
.C(n_220),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_219),
.A2(n_177),
.B1(n_180),
.B2(n_190),
.Y(n_234)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_238),
.A2(n_239),
.B1(n_235),
.B2(n_241),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_218),
.A2(n_200),
.B1(n_188),
.B2(n_178),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_216),
.B(n_193),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_207),
.A2(n_184),
.B1(n_199),
.B2(n_189),
.Y(n_242)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_187),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_246),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_137),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_111),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_239),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_75),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_249),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_33),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_33),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_33),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_251),
.B(n_253),
.C(n_259),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_263),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_231),
.B(n_229),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_255),
.B(n_262),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_226),
.C(n_209),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_257),
.C(n_266),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_226),
.C(n_209),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_55),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_17),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_237),
.A2(n_18),
.B1(n_26),
.B2(n_29),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_265),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_238),
.A2(n_29),
.B1(n_26),
.B2(n_18),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_55),
.C(n_33),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_21),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_21),
.C(n_17),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_21),
.Y(n_281)
);

AO221x1_ASAP7_75t_L g269 ( 
.A1(n_261),
.A2(n_232),
.B1(n_248),
.B2(n_243),
.C(n_240),
.Y(n_269)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_269),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_260),
.Y(n_270)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_252),
.A2(n_230),
.B1(n_9),
.B2(n_10),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_6),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_267),
.B(n_230),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_275),
.A2(n_278),
.B(n_281),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_266),
.A2(n_24),
.B1(n_21),
.B2(n_17),
.Y(n_276)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_276),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_259),
.B(n_8),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_283),
.C(n_279),
.Y(n_288)
);

A2O1A1O1Ixp25_ASAP7_75t_L g282 ( 
.A1(n_251),
.A2(n_7),
.B(n_14),
.C(n_12),
.D(n_11),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_257),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_256),
.A2(n_15),
.B(n_12),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_285),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_258),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_258),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_289),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_288),
.A2(n_282),
.B1(n_1),
.B2(n_2),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_15),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_6),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_0),
.Y(n_294)
);

AOI21xp33_ASAP7_75t_L g305 ( 
.A1(n_294),
.A2(n_296),
.B(n_2),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_0),
.C(n_1),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_295),
.B(n_277),
.C(n_280),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_0),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_298),
.C(n_299),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_290),
.A2(n_15),
.B1(n_12),
.B2(n_10),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_0),
.C(n_1),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_301),
.C(n_306),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_292),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_305),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_3),
.C(n_4),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_291),
.Y(n_307)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_307),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_297),
.A2(n_288),
.B(n_293),
.Y(n_308)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_308),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_302),
.A2(n_289),
.B(n_8),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_3),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_5),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_314),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_5),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_310),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_319),
.B(n_320),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_317),
.B(n_307),
.C(n_311),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_315),
.B(n_312),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_322),
.Y(n_323)
);

AOI21x1_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_313),
.B(n_316),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_3),
.Y(n_325)
);

AO21x2_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_4),
.B(n_5),
.Y(n_326)
);


endmodule