module fake_jpeg_26157_n_236 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_236);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_236;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_33),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_25),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_39),
.A2(n_23),
.B1(n_15),
.B2(n_21),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_40),
.A2(n_44),
.B(n_46),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_51),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_23),
.B1(n_15),
.B2(n_20),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_23),
.B1(n_20),
.B2(n_19),
.Y(n_46)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_32),
.C(n_35),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_64),
.C(n_73),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_51),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_59),
.Y(n_94)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_51),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_62),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_63),
.B(n_66),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_32),
.C(n_35),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_40),
.A2(n_36),
.B1(n_31),
.B2(n_19),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_53),
.B1(n_43),
.B2(n_31),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_51),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_49),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_68),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_37),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_71),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_37),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_35),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_74),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_35),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_17),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_44),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_75),
.B(n_77),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_35),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_32),
.Y(n_91)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_63),
.A2(n_43),
.B1(n_18),
.B2(n_25),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_84),
.A2(n_93),
.B1(n_100),
.B2(n_73),
.Y(n_119)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_7),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_86),
.B(n_74),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_61),
.B(n_32),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_91),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_96),
.B1(n_101),
.B2(n_60),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_75),
.A2(n_43),
.B1(n_18),
.B2(n_28),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_69),
.A2(n_38),
.B1(n_34),
.B2(n_32),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_66),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_69),
.A2(n_28),
.B1(n_16),
.B2(n_26),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_55),
.B(n_70),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_102),
.A2(n_72),
.B(n_76),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_55),
.B(n_38),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_54),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_106),
.B(n_107),
.Y(n_147)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_111),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_71),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_112),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_104),
.B(n_86),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_58),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_87),
.A2(n_64),
.B1(n_77),
.B2(n_57),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_115),
.B1(n_118),
.B2(n_123),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_90),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_114),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_90),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_116),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_103),
.B(n_24),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_121),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_92),
.A2(n_57),
.B1(n_60),
.B2(n_79),
.Y(n_118)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_97),
.A2(n_60),
.B1(n_67),
.B2(n_80),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_120),
.A2(n_122),
.B1(n_82),
.B2(n_88),
.Y(n_130)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_67),
.B1(n_78),
.B2(n_68),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_96),
.A2(n_78),
.B1(n_59),
.B2(n_58),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_125),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_59),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_81),
.B(n_103),
.Y(n_126)
);

OAI32xp33_ASAP7_75t_L g139 ( 
.A1(n_126),
.A2(n_86),
.A3(n_98),
.B1(n_82),
.B2(n_88),
.Y(n_139)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_102),
.B(n_98),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_22),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_130),
.A2(n_146),
.B1(n_123),
.B2(n_118),
.Y(n_162)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_135),
.B(n_136),
.Y(n_164)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_138),
.A2(n_139),
.B1(n_143),
.B2(n_152),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_99),
.C(n_83),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_148),
.C(n_150),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_99),
.B1(n_83),
.B2(n_85),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_110),
.A2(n_16),
.B(n_22),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_144),
.A2(n_153),
.B(n_117),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_111),
.A2(n_83),
.B1(n_85),
.B2(n_26),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_105),
.B(n_116),
.C(n_114),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_113),
.A2(n_85),
.B1(n_24),
.B2(n_29),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_0),
.B(n_1),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_154),
.A2(n_161),
.B1(n_162),
.B2(n_152),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_126),
.Y(n_155)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_129),
.C(n_150),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_157),
.B(n_138),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_131),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_160),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_135),
.A2(n_124),
.B1(n_121),
.B2(n_108),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_127),
.B(n_119),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_165),
.A2(n_168),
.B1(n_169),
.B2(n_151),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_27),
.B1(n_6),
.B2(n_7),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_166),
.A2(n_167),
.B1(n_153),
.B2(n_149),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_27),
.B1(n_5),
.B2(n_9),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g168 ( 
.A1(n_145),
.A2(n_0),
.B(n_1),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_L g169 ( 
.A1(n_145),
.A2(n_0),
.B(n_2),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_171),
.Y(n_175)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_173),
.Y(n_180)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

XNOR2x2_ASAP7_75t_SL g174 ( 
.A(n_164),
.B(n_148),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_174),
.A2(n_186),
.B1(n_188),
.B2(n_168),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_159),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_184),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_178),
.A2(n_187),
.B1(n_133),
.B2(n_162),
.Y(n_190)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_183),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_165),
.Y(n_198)
);

NOR3xp33_ASAP7_75t_SL g183 ( 
.A(n_154),
.B(n_144),
.C(n_139),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_136),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_185),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_158),
.A2(n_133),
.B1(n_137),
.B2(n_141),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_178),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_157),
.C(n_156),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_192),
.C(n_199),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_156),
.C(n_129),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_141),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_196),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_167),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_188),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_198),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_143),
.C(n_166),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_169),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_191),
.C(n_198),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_200),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_210),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_203),
.B(n_9),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_181),
.Y(n_204)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_175),
.Y(n_206)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_209),
.B(n_3),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_183),
.C(n_176),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_5),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_5),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_202),
.A2(n_193),
.B(n_199),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_214),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_216),
.B(n_217),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_213),
.A2(n_208),
.B1(n_211),
.B2(n_205),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_223),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_207),
.C(n_10),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_220),
.B(n_222),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_215),
.A2(n_218),
.B1(n_2),
.B2(n_0),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_213),
.A2(n_3),
.B(n_4),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_3),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_219),
.Y(n_226)
);

AOI31xp33_ASAP7_75t_L g229 ( 
.A1(n_226),
.A2(n_228),
.A3(n_222),
.B(n_4),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_4),
.C(n_10),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_229),
.A2(n_230),
.B(n_231),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_10),
.C(n_11),
.Y(n_231)
);

A2O1A1O1Ixp25_ASAP7_75t_L g232 ( 
.A1(n_229),
.A2(n_2),
.B(n_11),
.C(n_12),
.D(n_226),
.Y(n_232)
);

BUFx24_ASAP7_75t_SL g234 ( 
.A(n_232),
.Y(n_234)
);

BUFx24_ASAP7_75t_SL g235 ( 
.A(n_234),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_233),
.Y(n_236)
);


endmodule