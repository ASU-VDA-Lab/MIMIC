module real_jpeg_16224_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_4),
.B1(n_15),
.B2(n_17),
.Y(n_14)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_2),
.A2(n_73),
.B1(n_76),
.B2(n_77),
.Y(n_72)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_2),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_2),
.A2(n_76),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

OAI22x1_ASAP7_75t_SL g343 ( 
.A1(n_2),
.A2(n_76),
.B1(n_344),
.B2(n_348),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g366 ( 
.A1(n_2),
.A2(n_76),
.B1(n_218),
.B2(n_367),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_3),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_3),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_3),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_5),
.A2(n_142),
.B1(n_146),
.B2(n_147),
.Y(n_141)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_5),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_5),
.A2(n_146),
.B1(n_228),
.B2(n_231),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g450 ( 
.A1(n_5),
.A2(n_146),
.B1(n_451),
.B2(n_454),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_6),
.B(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_6),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_6),
.A2(n_61),
.B1(n_124),
.B2(n_126),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_6),
.A2(n_61),
.B1(n_102),
.B2(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_6),
.B(n_361),
.Y(n_360)
);

OAI32xp33_ASAP7_75t_L g384 ( 
.A1(n_6),
.A2(n_385),
.A3(n_387),
.B1(n_389),
.B2(n_391),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_6),
.B(n_249),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_6),
.B(n_235),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_7),
.Y(n_159)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_7),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g199 ( 
.A(n_7),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g249 ( 
.A(n_7),
.Y(n_249)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_8),
.Y(n_116)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_8),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_8),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_8),
.Y(n_230)
);

BUFx5_ASAP7_75t_L g350 ( 
.A(n_8),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_8),
.Y(n_394)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_9),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_10),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_10),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_10),
.A2(n_85),
.B1(n_133),
.B2(n_137),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_10),
.B(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_10),
.A2(n_85),
.B1(n_270),
.B2(n_273),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_12),
.Y(n_105)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_12),
.Y(n_109)
);

BUFx4f_ASAP7_75t_L g145 ( 
.A(n_12),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g220 ( 
.A(n_12),
.Y(n_220)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_13),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_13),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_13),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_13),
.Y(n_87)
);

BUFx8_ASAP7_75t_L g94 ( 
.A(n_13),
.Y(n_94)
);

BUFx12f_ASAP7_75t_SL g15 ( 
.A(n_16),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_437),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_279),
.B(n_436),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_239),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_20),
.B(n_239),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_174),
.C(n_214),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_22),
.B(n_214),
.Y(n_285)
);

XNOR2x1_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_95),
.Y(n_22)
);

XOR2x1_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_62),
.Y(n_23)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_24),
.Y(n_241)
);

AOI21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_38),
.B(n_54),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2x1p5_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_26),
.B(n_55),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_26),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_26),
.B(n_204),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_26),
.Y(n_361)
);

AO22x2_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_30),
.B1(n_33),
.B2(n_35),
.Y(n_26)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_32),
.Y(n_136)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_33),
.Y(n_125)
);

INVxp67_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_34),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_34),
.Y(n_326)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_37),
.Y(n_331)
);

NOR2x1p5_ASAP7_75t_SL g276 ( 
.A(n_38),
.B(n_54),
.Y(n_276)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_39),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_39),
.B(n_269),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_45),
.B1(n_46),
.B2(n_50),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_41),
.B(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_66),
.B1(n_67),
.B2(n_69),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_43),
.Y(n_272)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_44),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g457 ( 
.A(n_44),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_48),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_53),
.Y(n_194)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_53),
.Y(n_275)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_60),
.Y(n_55)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_57),
.Y(n_205)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI32xp33_ASAP7_75t_L g324 ( 
.A1(n_60),
.A2(n_178),
.A3(n_325),
.B1(n_327),
.B2(n_332),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_61),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_61),
.B(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_61),
.A2(n_187),
.B(n_265),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_61),
.B(n_262),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_61),
.B(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_62),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_81),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_63),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_72),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_64),
.B(n_82),
.Y(n_212)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_64),
.Y(n_262)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_65),
.B(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_66),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_67),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_89)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_72),
.B(n_88),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_72),
.Y(n_260)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_74),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_77),
.Y(n_265)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_88),
.Y(n_81)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_85),
.B(n_163),
.Y(n_162)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_88),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_88),
.B(n_264),
.Y(n_296)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_91),
.Y(n_186)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_94),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_95),
.B(n_241),
.C(n_242),
.Y(n_240)
);

NAND2x1p5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_140),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_96),
.B(n_140),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_130),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_97),
.B(n_380),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_123),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_98),
.B(n_132),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_98),
.Y(n_254)
);

OA21x2_ASAP7_75t_L g294 ( 
.A1(n_98),
.A2(n_123),
.B(n_131),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_98),
.B(n_343),
.Y(n_342)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_112),
.Y(n_98)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_102),
.B1(n_106),
.B2(n_110),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g112 ( 
.A1(n_100),
.A2(n_113),
.B1(n_117),
.B2(n_121),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_107),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_111),
.Y(n_396)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_122),
.Y(n_347)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_123),
.Y(n_341)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_130),
.A2(n_253),
.B(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_130),
.B(n_342),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_131),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_131),
.B(n_343),
.Y(n_380)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_136),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_152),
.B(n_160),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_141),
.A2(n_196),
.B(n_200),
.Y(n_195)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_145),
.Y(n_415)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_152),
.B(n_165),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_152),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_152),
.B(n_217),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_152),
.B(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_154),
.Y(n_164)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_161),
.B(n_313),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_161),
.B(n_365),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_165),
.B(n_169),
.Y(n_161)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_170),
.Y(n_364)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_172),
.Y(n_224)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_174),
.B(n_285),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_202),
.C(n_210),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_175),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_195),
.Y(n_175)
);

XOR2x2_ASAP7_75t_SL g306 ( 
.A(n_176),
.B(n_195),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_182),
.B1(n_187),
.B2(n_189),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_181),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_199),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_200),
.B(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_201),
.A2(n_216),
.B(n_221),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_202),
.A2(n_210),
.B1(n_211),
.B2(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_202),
.Y(n_290)
);

AND2x2_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_209),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_203),
.B(n_268),
.Y(n_309)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_225),
.Y(n_214)
);

AOI21x1_ASAP7_75t_L g257 ( 
.A1(n_215),
.A2(n_226),
.B(n_237),
.Y(n_257)
);

OA21x2_ASAP7_75t_L g245 ( 
.A1(n_216),
.A2(n_246),
.B(n_250),
.Y(n_245)
);

AO21x1_ASAP7_75t_L g363 ( 
.A1(n_216),
.A2(n_364),
.B(n_365),
.Y(n_363)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx5_ASAP7_75t_L g369 ( 
.A(n_220),
.Y(n_369)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_220),
.Y(n_388)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp67_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_237),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_235),
.Y(n_226)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_227),
.Y(n_253)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_236),
.B(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_238),
.B(n_379),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_238),
.B(n_340),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_243),
.Y(n_239)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_240),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_256),
.B1(n_277),
.B2(n_278),
.Y(n_243)
);

INVxp67_ASAP7_75t_SL g278 ( 
.A(n_244),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_244),
.B(n_440),
.C(n_441),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_251),
.B1(n_252),
.B2(n_255),
.Y(n_244)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_245),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_245),
.B(n_324),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_245),
.A2(n_255),
.B1(n_324),
.B2(n_372),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_245),
.A2(n_255),
.B1(n_464),
.B2(n_465),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_245),
.B(n_252),
.Y(n_466)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_256),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_257),
.B(n_444),
.C(n_445),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_266),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_259),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_259)
);

AOI21x1_ASAP7_75t_L g464 ( 
.A1(n_261),
.A2(n_262),
.B(n_263),
.Y(n_464)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_266),
.Y(n_444)
);

NOR2x1_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_276),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_276),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_277),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_316),
.B(n_432),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_301),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_283),
.B(n_435),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g433 ( 
.A(n_284),
.B(n_286),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_291),
.C(n_300),
.Y(n_286)
);

INVxp67_ASAP7_75t_SL g287 ( 
.A(n_288),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_288),
.B(n_315),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_300),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_295),
.C(n_297),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_294),
.B1(n_297),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_294),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_295),
.B(n_304),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_297),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_298),
.B(n_376),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_299),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_314),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_302),
.B(n_314),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_306),
.C(n_307),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_303),
.B(n_352),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_306),
.Y(n_353)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.C(n_311),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_321),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_310),
.A2(n_311),
.B1(n_312),
.B2(n_322),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_310),
.Y(n_322)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_313),
.B(n_405),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_354),
.B(n_431),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_351),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_319),
.B(n_351),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_323),
.C(n_337),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_320),
.B(n_427),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_323),
.A2(n_337),
.B1(n_338),
.B2(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_323),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_324),
.Y(n_372)
);

INVx6_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_326),
.Y(n_336)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_336),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_342),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_350),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_425),
.B(n_430),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_356),
.A2(n_381),
.B(n_424),
.Y(n_355)
);

NOR2xp67_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_370),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_357),
.B(n_370),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_360),
.C(n_362),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_358),
.A2(n_359),
.B1(n_360),
.B2(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_360),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_361),
.A2(n_449),
.B(n_458),
.Y(n_448)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_363),
.B(n_399),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_366),
.B(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_371),
.B(n_373),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_371),
.B(n_375),
.C(n_377),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_374),
.A2(n_375),
.B1(n_377),
.B2(n_378),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

AOI21x1_ASAP7_75t_L g381 ( 
.A1(n_382),
.A2(n_401),
.B(n_423),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_398),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_SL g423 ( 
.A(n_383),
.B(n_398),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_397),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_384),
.B(n_397),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_395),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_402),
.A2(n_409),
.B(n_422),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_408),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_403),
.B(n_408),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_410),
.A2(n_418),
.B(n_421),
.Y(n_409)
);

NOR2xp67_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_417),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_416),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_419),
.B(n_420),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_419),
.B(n_420),
.Y(n_421)
);

NAND2xp33_ASAP7_75t_SL g425 ( 
.A(n_426),
.B(n_429),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_426),
.B(n_429),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_SL g432 ( 
.A(n_433),
.B(n_434),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_470),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_442),
.Y(n_438)
);

NOR2x1p5_ASAP7_75t_L g470 ( 
.A(n_439),
.B(n_442),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_446),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_447),
.A2(n_461),
.B1(n_468),
.B2(n_469),
.Y(n_446)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_447),
.Y(n_469)
);

OA21x2_ASAP7_75t_L g447 ( 
.A1(n_448),
.A2(n_459),
.B(n_460),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_448),
.B(n_459),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_461),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_462),
.A2(n_463),
.B1(n_466),
.B2(n_467),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_464),
.Y(n_465)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_466),
.Y(n_467)
);


endmodule