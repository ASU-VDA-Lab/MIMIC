module fake_jpeg_29330_n_452 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_452);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_452;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_8),
.B(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_13),
.B(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_47),
.Y(n_126)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_49),
.B(n_81),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_16),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_55),
.B(n_63),
.Y(n_134)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_58),
.B(n_59),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_60),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_16),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_64),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_65),
.Y(n_135)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_71),
.Y(n_146)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_35),
.B(n_16),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_73),
.B(n_80),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_32),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_74),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_75),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_77),
.Y(n_145)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_29),
.Y(n_78)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

CKINVDCx12_ASAP7_75t_R g79 ( 
.A(n_34),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_23),
.Y(n_81)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

INVx6_ASAP7_75t_SL g84 ( 
.A(n_40),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_86),
.Y(n_96)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_17),
.B(n_15),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_92),
.Y(n_106)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_17),
.B(n_14),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_18),
.Y(n_93)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_84),
.A2(n_45),
.B1(n_23),
.B2(n_24),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_99),
.A2(n_112),
.B1(n_136),
.B2(n_25),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_78),
.A2(n_45),
.B1(n_23),
.B2(n_24),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_55),
.B(n_32),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_114),
.B(n_140),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_74),
.A2(n_32),
.B1(n_46),
.B2(n_26),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_115),
.A2(n_138),
.B1(n_144),
.B2(n_72),
.Y(n_177)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_51),
.Y(n_117)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_119),
.Y(n_192)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_48),
.A2(n_19),
.B1(n_41),
.B2(n_37),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_124),
.A2(n_21),
.B1(n_33),
.B2(n_22),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_47),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_131),
.B(n_125),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_86),
.A2(n_24),
.B1(n_34),
.B2(n_25),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_52),
.Y(n_137)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_L g138 ( 
.A1(n_50),
.A2(n_19),
.B1(n_41),
.B2(n_37),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_46),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_53),
.A2(n_26),
.B1(n_21),
.B2(n_33),
.Y(n_144)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_150),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_151),
.A2(n_177),
.B1(n_187),
.B2(n_126),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_27),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_152),
.B(n_158),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_106),
.B(n_59),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_153),
.B(n_159),
.Y(n_219)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_154),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_142),
.A2(n_71),
.B1(n_61),
.B2(n_64),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_156),
.A2(n_147),
.B1(n_146),
.B2(n_135),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_94),
.B(n_22),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_68),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_160),
.B(n_162),
.Y(n_235)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_105),
.Y(n_161)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_161),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_101),
.B(n_91),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_104),
.Y(n_163)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_163),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_14),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_164),
.B(n_181),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_96),
.Y(n_165)
);

BUFx2_ASAP7_75t_SL g207 ( 
.A(n_165),
.Y(n_207)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_112),
.A2(n_56),
.B(n_27),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_167),
.B(n_170),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_123),
.Y(n_168)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_168),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_116),
.B(n_76),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_169),
.B(n_172),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_62),
.C(n_65),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_129),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_171),
.B(n_175),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_111),
.B(n_75),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_123),
.Y(n_173)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_113),
.A2(n_120),
.B(n_141),
.C(n_139),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_174),
.A2(n_158),
.B(n_165),
.C(n_176),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_148),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_108),
.B(n_138),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_176),
.B(n_186),
.Y(n_238)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_103),
.Y(n_178)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_178),
.Y(n_208)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_122),
.Y(n_179)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_179),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_100),
.Y(n_180)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_180),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_122),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_124),
.B(n_83),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_182),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_99),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_183),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_136),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_109),
.B(n_47),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_133),
.B(n_0),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_95),
.B(n_80),
.Y(n_188)
);

FAx1_ASAP7_75t_SL g218 ( 
.A(n_188),
.B(n_190),
.CI(n_194),
.CON(n_218),
.SN(n_218)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_110),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_189),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_95),
.B(n_80),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_133),
.B(n_86),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_191),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_143),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_193),
.Y(n_233)
);

AND2x2_ASAP7_75t_SL g194 ( 
.A(n_110),
.B(n_0),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_97),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_195),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_107),
.B(n_77),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_196),
.B(n_60),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_102),
.B(n_77),
.Y(n_197)
);

FAx1_ASAP7_75t_SL g220 ( 
.A(n_197),
.B(n_199),
.CI(n_97),
.CON(n_220),
.SN(n_220)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_198),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_102),
.B(n_67),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_98),
.Y(n_200)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_98),
.Y(n_201)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_203),
.A2(n_216),
.B1(n_230),
.B2(n_240),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_152),
.A2(n_97),
.B(n_126),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_214),
.A2(n_149),
.B(n_178),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_220),
.B(n_179),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_222),
.B(n_4),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_167),
.A2(n_130),
.B1(n_60),
.B2(n_67),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_223),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_154),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_228),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_177),
.A2(n_147),
.B1(n_146),
.B2(n_135),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_193),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_180),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_172),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_182),
.A2(n_132),
.B1(n_127),
.B2(n_82),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_169),
.Y(n_241)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_241),
.Y(n_246)
);

AOI32xp33_ASAP7_75t_L g244 ( 
.A1(n_185),
.A2(n_130),
.A3(n_132),
.B1(n_127),
.B2(n_3),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_189),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_170),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_245),
.A2(n_151),
.B1(n_194),
.B2(n_156),
.Y(n_250)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_215),
.Y(n_247)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_247),
.Y(n_295)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_248),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_250),
.B(n_261),
.Y(n_286)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_251),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_213),
.A2(n_241),
.B1(n_225),
.B2(n_217),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_252),
.A2(n_263),
.B1(n_267),
.B2(n_270),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_196),
.C(n_186),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_253),
.B(n_255),
.Y(n_313)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_232),
.Y(n_254)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_254),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_199),
.C(n_197),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_226),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_256),
.B(n_258),
.Y(n_290)
);

XNOR2x1_ASAP7_75t_L g316 ( 
.A(n_257),
.B(n_259),
.Y(n_316)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_205),
.Y(n_258)
);

MAJx2_ASAP7_75t_L g259 ( 
.A(n_210),
.B(n_164),
.C(n_174),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_260),
.B(n_264),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_238),
.A2(n_190),
.B1(n_188),
.B2(n_192),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_217),
.A2(n_194),
.B1(n_155),
.B2(n_161),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_235),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_242),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_265),
.B(n_272),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_238),
.A2(n_149),
.B1(n_150),
.B2(n_168),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_276),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_202),
.A2(n_173),
.B1(n_163),
.B2(n_201),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_268),
.A2(n_271),
.B(n_274),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_202),
.A2(n_222),
.B1(n_211),
.B2(n_203),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_239),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_210),
.B(n_157),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_237),
.A2(n_157),
.B1(n_200),
.B2(n_166),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_275),
.B(n_281),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_237),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_277),
.B(n_278),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_219),
.B(n_4),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_214),
.A2(n_5),
.B(n_6),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_279),
.A2(n_284),
.B(n_263),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_224),
.Y(n_280)
);

INVxp33_ASAP7_75t_SL g301 ( 
.A(n_280),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_224),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_208),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_282),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_218),
.B(n_220),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_284),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_218),
.B(n_6),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_218),
.B(n_12),
.C(n_9),
.Y(n_285)
);

MAJx2_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_239),
.C(n_231),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_271),
.A2(n_283),
.B(n_279),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_293),
.B(n_304),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_296),
.B(n_299),
.Y(n_328)
);

AOI31xp33_ASAP7_75t_L g297 ( 
.A1(n_259),
.A2(n_207),
.A3(n_211),
.B(n_252),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_297),
.B(n_298),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_268),
.A2(n_220),
.B(n_212),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_273),
.B(n_204),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_262),
.A2(n_212),
.B(n_228),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_300),
.B(n_314),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_246),
.A2(n_206),
.B1(n_205),
.B2(n_208),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_302),
.A2(n_317),
.B1(n_319),
.B2(n_269),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_260),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_305),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_262),
.A2(n_231),
.B1(n_243),
.B2(n_233),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_307),
.A2(n_269),
.B1(n_227),
.B2(n_258),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_254),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_311),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_253),
.A2(n_243),
.B(n_206),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_312),
.B(n_320),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_246),
.B(n_234),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_249),
.A2(n_270),
.B1(n_250),
.B2(n_255),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_249),
.A2(n_229),
.B1(n_209),
.B2(n_221),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_285),
.A2(n_233),
.B(n_227),
.Y(n_320)
);

BUFx24_ASAP7_75t_SL g323 ( 
.A(n_308),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_323),
.B(n_332),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_264),
.Y(n_324)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_324),
.Y(n_355)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_314),
.Y(n_325)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_325),
.Y(n_366)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_301),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_326),
.B(n_341),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_327),
.A2(n_330),
.B1(n_310),
.B2(n_288),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_261),
.Y(n_329)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_329),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_286),
.A2(n_266),
.B1(n_257),
.B2(n_281),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_331),
.A2(n_346),
.B1(n_349),
.B2(n_310),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_295),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_317),
.A2(n_276),
.B1(n_272),
.B2(n_256),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_333),
.A2(n_287),
.B1(n_286),
.B2(n_305),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_315),
.B(n_248),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_335),
.B(n_336),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_291),
.B(n_247),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_313),
.B(n_251),
.C(n_232),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_337),
.B(n_342),
.C(n_343),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_291),
.B(n_209),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_339),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_318),
.Y(n_340)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_340),
.Y(n_352)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_295),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_313),
.B(n_229),
.C(n_221),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_316),
.B(n_8),
.C(n_9),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_303),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_344),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_316),
.B(n_8),
.C(n_10),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_345),
.B(n_304),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_290),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_290),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_351),
.A2(n_353),
.B1(n_363),
.B2(n_374),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_331),
.A2(n_293),
.B1(n_287),
.B2(n_294),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_338),
.B(n_316),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_356),
.B(n_365),
.Y(n_387)
);

INVx3_ASAP7_75t_SL g357 ( 
.A(n_326),
.Y(n_357)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_357),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_358),
.B(n_359),
.Y(n_380)
);

OA22x2_ASAP7_75t_L g359 ( 
.A1(n_325),
.A2(n_298),
.B1(n_288),
.B2(n_319),
.Y(n_359)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_362),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_321),
.A2(n_306),
.B1(n_296),
.B2(n_289),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_334),
.A2(n_347),
.B(n_328),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_364),
.B(n_372),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_338),
.B(n_289),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_330),
.A2(n_310),
.B1(n_292),
.B2(n_300),
.Y(n_369)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_369),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_348),
.B(n_312),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_371),
.B(n_343),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_321),
.A2(n_310),
.B1(n_292),
.B2(n_302),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_373),
.B(n_320),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_333),
.A2(n_328),
.B1(n_334),
.B2(n_342),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_361),
.B(n_337),
.C(n_348),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_375),
.B(n_378),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_370),
.Y(n_376)
);

NAND3xp33_ASAP7_75t_L g395 ( 
.A(n_376),
.B(n_379),
.C(n_386),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_361),
.B(n_299),
.C(n_304),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_350),
.B(n_306),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_383),
.B(n_384),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_371),
.B(n_356),
.C(n_373),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_365),
.B(n_345),
.Y(n_385)
);

XNOR2x1_ASAP7_75t_L g410 ( 
.A(n_385),
.B(n_388),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_370),
.Y(n_386)
);

XNOR2x1_ASAP7_75t_L g390 ( 
.A(n_374),
.B(n_297),
.Y(n_390)
);

A2O1A1O1Ixp25_ASAP7_75t_L g399 ( 
.A1(n_390),
.A2(n_360),
.B(n_359),
.C(n_372),
.D(n_358),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_353),
.B(n_349),
.C(n_346),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_391),
.A2(n_354),
.B(n_326),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_355),
.B(n_322),
.Y(n_393)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_393),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_364),
.B(n_344),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_394),
.B(n_369),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_396),
.B(n_397),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_381),
.A2(n_389),
.B1(n_380),
.B2(n_392),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_394),
.A2(n_351),
.B1(n_368),
.B2(n_366),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_398),
.B(n_403),
.Y(n_417)
);

OAI21xp33_ASAP7_75t_L g413 ( 
.A1(n_399),
.A2(n_359),
.B(n_387),
.Y(n_413)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_393),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_402),
.B(n_404),
.Y(n_415)
);

AO221x1_ASAP7_75t_L g403 ( 
.A1(n_377),
.A2(n_352),
.B1(n_341),
.B2(n_318),
.C(n_303),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_391),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_405),
.B(n_406),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_382),
.A2(n_367),
.B1(n_322),
.B2(n_354),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_390),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_408),
.Y(n_422)
);

AO221x1_ASAP7_75t_L g408 ( 
.A1(n_383),
.A2(n_352),
.B1(n_309),
.B2(n_357),
.C(n_340),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_375),
.A2(n_359),
.B1(n_340),
.B2(n_309),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_409),
.B(n_387),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_395),
.A2(n_378),
.B(n_384),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_412),
.B(n_401),
.Y(n_427)
);

XNOR2x1_ASAP7_75t_L g424 ( 
.A(n_413),
.B(n_396),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_400),
.B(n_311),
.Y(n_414)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_414),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_411),
.A2(n_385),
.B(n_388),
.Y(n_416)
);

CKINVDCx14_ASAP7_75t_R g426 ( 
.A(n_416),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_418),
.B(n_396),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_SL g420 ( 
.A1(n_399),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_420),
.B(n_398),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_411),
.B(n_11),
.C(n_12),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_423),
.B(n_414),
.Y(n_428)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_424),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_427),
.B(n_428),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_419),
.B(n_401),
.C(n_409),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_429),
.B(n_430),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_415),
.B(n_397),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_431),
.B(n_421),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_432),
.B(n_433),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_417),
.B(n_12),
.Y(n_433)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_437),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_429),
.B(n_422),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_438),
.B(n_440),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_426),
.B(n_418),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_435),
.A2(n_425),
.B(n_420),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_443),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_436),
.A2(n_432),
.B(n_424),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_444),
.B(n_434),
.C(n_431),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_445),
.Y(n_448)
);

AOI21xp33_ASAP7_75t_L g446 ( 
.A1(n_441),
.A2(n_442),
.B(n_439),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_448),
.B(n_447),
.C(n_446),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_449),
.B(n_437),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_450),
.B(n_413),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_451),
.B(n_410),
.C(n_436),
.Y(n_452)
);


endmodule