module real_jpeg_14275_n_7 (n_5, n_4, n_0, n_1, n_2, n_6, n_3, n_7);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_3;

output n_7;

wire n_17;
wire n_8;
wire n_57;
wire n_54;
wire n_37;
wire n_21;
wire n_43;
wire n_35;
wire n_33;
wire n_38;
wire n_50;
wire n_29;
wire n_55;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_12;
wire n_24;
wire n_34;
wire n_44;
wire n_28;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_51;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_48;
wire n_30;
wire n_56;
wire n_16;
wire n_15;
wire n_13;

INVx4_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_2),
.A2(n_11),
.B1(n_12),
.B2(n_19),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_2),
.A2(n_19),
.B1(n_42),
.B2(n_44),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_4),
.A2(n_11),
.B1(n_12),
.B2(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_5),
.B(n_14),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_5),
.A2(n_11),
.B1(n_12),
.B2(n_23),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_5),
.B(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_5),
.A2(n_23),
.B1(n_42),
.B2(n_44),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_5),
.B(n_11),
.C(n_32),
.Y(n_51)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

XNOR2xp5_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_35),
.Y(n_7)
);

AOI21xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_24),
.B(n_34),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_16),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_13),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_15),
.Y(n_21)
);

AO22x1_ASAP7_75t_L g31 ( 
.A1(n_11),
.A2(n_12),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_20),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_22),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_21),
.B(n_28),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_49),
.Y(n_48)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_32),
.A2(n_33),
.B1(n_42),
.B2(n_44),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_57),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_54),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_54),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_38)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_45),
.Y(n_39)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_51),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_48),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_50),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);


endmodule