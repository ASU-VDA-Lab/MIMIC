module fake_jpeg_3928_n_175 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_175);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_34),
.B1(n_27),
.B2(n_25),
.Y(n_41)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_24),
.B(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_28),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_38),
.Y(n_48)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_17),
.B1(n_28),
.B2(n_27),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_39),
.A2(n_47),
.B1(n_52),
.B2(n_33),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_31),
.A2(n_29),
.B1(n_24),
.B2(n_26),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_16),
.B1(n_14),
.B2(n_19),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_29),
.B1(n_26),
.B2(n_21),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_49),
.B(n_23),
.C(n_38),
.Y(n_54)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_34),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_31),
.A2(n_21),
.B1(n_22),
.B2(n_18),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_23),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_20),
.Y(n_51)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_15),
.B1(n_14),
.B2(n_19),
.Y(n_52)
);

AOI21xp33_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_36),
.B(n_35),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_53),
.A2(n_54),
.B(n_66),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_57),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_30),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_40),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_34),
.B1(n_32),
.B2(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_61),
.Y(n_88)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_63),
.Y(n_91)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_64),
.B(n_72),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_51),
.B(n_1),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_65),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_45),
.A2(n_38),
.B1(n_32),
.B2(n_49),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_15),
.B1(n_33),
.B2(n_18),
.Y(n_67)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_49),
.A2(n_15),
.B1(n_16),
.B2(n_14),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_71),
.B(n_74),
.Y(n_76)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_69),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_87),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_41),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_81),
.A2(n_94),
.B(n_3),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_47),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_30),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_78),
.C(n_79),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_60),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_86),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_40),
.Y(n_87)
);

NOR2x1_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_50),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_SL g98 ( 
.A1(n_92),
.A2(n_55),
.B(n_42),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_60),
.B(n_52),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_93),
.B(n_95),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_30),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_63),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_96),
.B(n_100),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_98),
.A2(n_101),
.B1(n_108),
.B2(n_83),
.Y(n_128)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_30),
.B(n_42),
.C(n_14),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_99),
.A2(n_90),
.B(n_83),
.Y(n_127)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_30),
.B1(n_42),
.B2(n_9),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_1),
.Y(n_102)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_76),
.C(n_90),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_77),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_110),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_107),
.A2(n_94),
.B1(n_95),
.B2(n_81),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_8),
.B1(n_12),
.B2(n_6),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_109),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_3),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_3),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_111),
.A2(n_114),
.B(n_89),
.Y(n_122)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_113),
.Y(n_126)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_122),
.B(n_114),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_78),
.Y(n_119)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

XOR2x2_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_81),
.Y(n_120)
);

XOR2x1_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_111),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_129),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_104),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_125),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_109),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_111),
.B(n_88),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_127),
.A2(n_128),
.B1(n_99),
.B2(n_107),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_108),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_101),
.B1(n_82),
.B2(n_106),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_131),
.A2(n_127),
.B1(n_118),
.B2(n_10),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_133),
.B(n_139),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_140),
.C(n_117),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_107),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_136),
.B(n_142),
.Y(n_147)
);

INVxp33_ASAP7_75t_SL g138 ( 
.A(n_121),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_138),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_125),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_130),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_126),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_6),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_133),
.A2(n_119),
.B(n_124),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_144),
.A2(n_151),
.B(n_137),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_152),
.C(n_140),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_115),
.Y(n_151)
);

MAJx2_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_120),
.C(n_122),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_7),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_155),
.Y(n_166)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_156),
.Y(n_162)
);

AO21x1_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_138),
.B(n_132),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_158),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_147),
.B(n_134),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_159),
.A2(n_150),
.B1(n_148),
.B2(n_4),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_11),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_145),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_R g169 ( 
.A1(n_161),
.A2(n_165),
.B1(n_133),
.B2(n_153),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_162),
.Y(n_168)
);

NOR2xp67_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_13),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_164),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_168),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_166),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_166),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_172),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_170),
.Y(n_173)
);

XNOR2x2_ASAP7_75t_SL g175 ( 
.A(n_174),
.B(n_173),
.Y(n_175)
);


endmodule