module fake_jpeg_18226_n_45 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_45);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_45;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx6_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx2_ASAP7_75t_SL g10 ( 
.A(n_3),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_2),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx24_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_5),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_16),
.B(n_17),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_15),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_1),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_15),
.B(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_1),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_1),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_12),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_SL g23 ( 
.A1(n_7),
.A2(n_6),
.B(n_12),
.C(n_14),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_23),
.A2(n_7),
.B1(n_8),
.B2(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_12),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_8),
.Y(n_25)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_21),
.Y(n_34)
);

OAI322xp33_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_37),
.A3(n_27),
.B1(n_23),
.B2(n_29),
.C1(n_26),
.C2(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_26),
.B1(n_33),
.B2(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_40),
.Y(n_41)
);

AOI322xp5_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_23),
.A3(n_25),
.B1(n_29),
.B2(n_31),
.C1(n_36),
.C2(n_39),
.Y(n_42)
);

MAJx2_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_23),
.C(n_31),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_44),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);


endmodule