module fake_jpeg_6573_n_314 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_314);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_48),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_41),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_15),
.B(n_7),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_34),
.Y(n_57)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_40),
.B(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_33),
.Y(n_72)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_22),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_50),
.B(n_68),
.Y(n_125)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_52),
.B(n_56),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_57),
.B(n_62),
.Y(n_103)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_58),
.B(n_64),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_31),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_60),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_31),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_18),
.C(n_28),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_61),
.B(n_32),
.C(n_20),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_22),
.Y(n_62)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_67),
.B(n_69),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_39),
.B(n_18),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_41),
.A2(n_29),
.B1(n_16),
.B2(n_34),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_71),
.A2(n_95),
.B1(n_99),
.B2(n_20),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_72),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_39),
.A2(n_29),
.B1(n_28),
.B2(n_25),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_73),
.A2(n_97),
.B1(n_19),
.B2(n_30),
.Y(n_119)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_17),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_75),
.B(n_77),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_25),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_27),
.Y(n_78)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

BUFx2_ASAP7_75t_SL g124 ( 
.A(n_79),
.Y(n_124)
);

CKINVDCx12_ASAP7_75t_R g80 ( 
.A(n_36),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_27),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_83),
.B(n_86),
.Y(n_112)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_42),
.B(n_24),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_87),
.B(n_88),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_42),
.B(n_16),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_24),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_90),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_42),
.B(n_12),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_42),
.B(n_12),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_94),
.Y(n_114)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_47),
.B(n_20),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_47),
.A2(n_33),
.B1(n_26),
.B2(n_23),
.Y(n_95)
);

OR2x4_ASAP7_75t_L g96 ( 
.A(n_38),
.B(n_30),
.Y(n_96)
);

OR2x2_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_98),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_L g97 ( 
.A1(n_44),
.A2(n_33),
.B1(n_26),
.B2(n_32),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_41),
.A2(n_26),
.B1(n_19),
.B2(n_30),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_62),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_96),
.A2(n_14),
.B1(n_19),
.B2(n_30),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_71),
.B1(n_95),
.B2(n_99),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_119),
.A2(n_85),
.B1(n_63),
.B2(n_20),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_55),
.B(n_30),
.C(n_19),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_66),
.C(n_49),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_53),
.B1(n_64),
.B2(n_81),
.Y(n_155)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_132),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_130),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_131),
.B(n_113),
.C(n_126),
.Y(n_172)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_52),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_143),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_62),
.B(n_75),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_134),
.A2(n_128),
.B1(n_105),
.B2(n_79),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_135),
.Y(n_183)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_136),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

INVx3_ASAP7_75t_SL g191 ( 
.A(n_137),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_100),
.B(n_57),
.Y(n_138)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_138),
.Y(n_175)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

INVx13_ASAP7_75t_L g199 ( 
.A(n_139),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_140),
.A2(n_155),
.B1(n_160),
.B2(n_105),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_141),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_110),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_142),
.B(n_148),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_57),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_58),
.Y(n_144)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_144),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_100),
.B(n_54),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_146),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_100),
.B(n_75),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_104),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_147),
.Y(n_198)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_149),
.Y(n_201)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_154),
.Y(n_179)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_111),
.B(n_70),
.Y(n_152)
);

BUFx24_ASAP7_75t_SL g185 ( 
.A(n_152),
.Y(n_185)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_97),
.B1(n_92),
.B2(n_82),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_153),
.A2(n_159),
.B1(n_161),
.B2(n_164),
.Y(n_167)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_112),
.A2(n_84),
.B(n_73),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_156),
.A2(n_103),
.B(n_117),
.Y(n_170)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_101),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_120),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_110),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_163),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_119),
.A2(n_53),
.B1(n_61),
.B2(n_63),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_103),
.A2(n_85),
.B1(n_3),
.B2(n_4),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_112),
.A2(n_79),
.B(n_76),
.C(n_65),
.Y(n_162)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_162),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_125),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_126),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_170),
.A2(n_192),
.B(n_193),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_172),
.B(n_178),
.C(n_116),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_146),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_137),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_153),
.A2(n_141),
.B1(n_156),
.B2(n_143),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_174),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_153),
.A2(n_117),
.B1(n_125),
.B2(n_104),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_177),
.Y(n_208)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_109),
.C(n_120),
.Y(n_178)
);

NOR3xp33_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_193),
.C(n_175),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_184),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_110),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_194),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_0),
.Y(n_227)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_195),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_153),
.A2(n_51),
.B(n_76),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_148),
.A2(n_51),
.B(n_65),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_0),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_159),
.A2(n_128),
.B1(n_106),
.B2(n_6),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_176),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_166),
.A2(n_150),
.B1(n_152),
.B2(n_136),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_203),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_165),
.B(n_129),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_204),
.B(n_205),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_164),
.Y(n_205)
);

BUFx24_ASAP7_75t_SL g207 ( 
.A(n_177),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_207),
.B(n_212),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_213),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_170),
.A2(n_132),
.B(n_139),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_210),
.A2(n_214),
.B(n_223),
.Y(n_232)
);

BUFx24_ASAP7_75t_SL g212 ( 
.A(n_173),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_166),
.A2(n_195),
.B(n_190),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_168),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_215),
.B(n_218),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_192),
.A2(n_149),
.B1(n_106),
.B2(n_135),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_216),
.A2(n_196),
.B1(n_186),
.B2(n_178),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_217),
.A2(n_214),
.B1(n_219),
.B2(n_211),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_179),
.B(n_116),
.Y(n_218)
);

MAJx2_ASAP7_75t_L g220 ( 
.A(n_169),
.B(n_116),
.C(n_151),
.Y(n_220)
);

OAI322xp33_ASAP7_75t_L g242 ( 
.A1(n_220),
.A2(n_171),
.A3(n_194),
.B1(n_200),
.B2(n_191),
.C1(n_185),
.C2(n_187),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_221),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_147),
.Y(n_222)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_222),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_174),
.A2(n_172),
.B(n_167),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_181),
.B(n_8),
.Y(n_225)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_225),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_106),
.Y(n_226)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_171),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_180),
.A2(n_0),
.B(n_5),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_228),
.A2(n_191),
.B(n_198),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_218),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_237),
.Y(n_256)
);

NOR3xp33_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_242),
.C(n_219),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_224),
.A2(n_167),
.B1(n_189),
.B2(n_180),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_235),
.A2(n_238),
.B1(n_216),
.B2(n_215),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_220),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_224),
.A2(n_200),
.B1(n_184),
.B2(n_179),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_250),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_245),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_203),
.B(n_197),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_208),
.A2(n_191),
.B1(n_201),
.B2(n_188),
.Y(n_246)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_247),
.A2(n_204),
.B(n_206),
.Y(n_251)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_202),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_251),
.A2(n_265),
.B(n_266),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_213),
.C(n_223),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_253),
.C(n_258),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_209),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_187),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_255),
.B(n_229),
.Y(n_273)
);

NOR3xp33_ASAP7_75t_SL g281 ( 
.A(n_257),
.B(n_10),
.C(n_13),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_206),
.C(n_210),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_246),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_264),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_227),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_263),
.C(n_267),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_202),
.C(n_205),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_240),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_247),
.A2(n_237),
.B(n_250),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_228),
.C(n_188),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_262),
.A2(n_248),
.B1(n_243),
.B2(n_245),
.Y(n_269)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_269),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_233),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_281),
.Y(n_282)
);

XNOR2x1_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_241),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_5),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_267),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_254),
.A2(n_243),
.B1(n_244),
.B2(n_241),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_275),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_266),
.A2(n_239),
.B1(n_249),
.B2(n_236),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_276),
.B(n_198),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_249),
.C(n_230),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_278),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_236),
.C(n_183),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_183),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_279),
.A2(n_260),
.B(n_263),
.Y(n_287)
);

INVxp67_ASAP7_75t_SL g283 ( 
.A(n_279),
.Y(n_283)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_283),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_284),
.B(n_288),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_271),
.A2(n_251),
.B1(n_261),
.B2(n_265),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_285),
.A2(n_274),
.B1(n_268),
.B2(n_6),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_287),
.A2(n_280),
.B(n_278),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_291),
.Y(n_299)
);

OA21x2_ASAP7_75t_L g292 ( 
.A1(n_272),
.A2(n_6),
.B(n_7),
.Y(n_292)
);

AO21x1_ASAP7_75t_L g298 ( 
.A1(n_292),
.A2(n_7),
.B(n_8),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_297),
.B1(n_301),
.B2(n_299),
.Y(n_304)
);

AOI21x1_ASAP7_75t_L g294 ( 
.A1(n_283),
.A2(n_270),
.B(n_281),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_296),
.Y(n_306)
);

AOI322xp5_ASAP7_75t_L g295 ( 
.A1(n_290),
.A2(n_277),
.A3(n_274),
.B1(n_268),
.B2(n_10),
.C1(n_11),
.C2(n_13),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_282),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_299),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_285),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_289),
.C(n_286),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_304),
.C(n_292),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_292),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_308),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_298),
.Y(n_309)
);

OAI21x1_ASAP7_75t_L g311 ( 
.A1(n_309),
.A2(n_310),
.B(n_303),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_10),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_311),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_312),
.Y(n_314)
);


endmodule